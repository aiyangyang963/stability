
module issp_Ch1_dat_abs (
	source,
	source_ena,
	probe,
	source_clk);	

	output	[15:0]	source;
	input		source_ena;
	input	[0:0]	probe;
	input		source_clk;
endmodule
