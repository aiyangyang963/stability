-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kBFK1LoH6M77sVErtgJSfdnvtLItFsldt0xqXdZ7mTDQK4MA2Sntnsm3YYiu4cSGbuCRY/NCGufH
1dvjkay+UEnnrBD+F9oQNsyObT8vAzhiGSugpVHpJNd0nxtNo5SgWGXnUiAaZ1JdGDV4X1gz5dxs
u4BshIpXYRRi2+Do643wkY3nY1Yz4pvv1ueGHSwMm0d2wrDlouNHcv4Eu+M/w/2CzmB0FFF0ga5y
egtIVupf8tUlf9Fbrz0QL1i9yEDfRzHKF2dEzPKFlQKNpO85BvYmElEOhJ6/5L6iVl+jmZ8HHFmd
YXlyFq4kPIn+9g7up+Vk4/TLiLbjJg9f40mMKQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
zifMk3QQG5xNzec465EQaGuRZYb3bXgwpP8QEbjvd0aD2qdi/2pHgkfq9ngT2Ps72ZI2ZQT5I8V+
K5MAiLALZSqHyX5izTjOYjqoAoFiTc7WkpAbQ7Zj18dhI0nomVR+O3PrGC6oZTnqzz5pRsdIIanB
S0xHki+trYFQJikJDkv/Zam19iLGGJ3VA0tb6iLwkISvbf53oALU7u07RtDP75P8+UuWS1B2lZv3
O/WJyPKP3SMxJVG9GoD3MXR00Q8IAofGOU2U2W8wSsuJaovhaCJK2MUhb0pBUnammtwcP9W2nN0r
plFFfR9wCOhKpx7m8wT9iywzx+W0gSyIak8kTsRqFm2wLj4AaJOKOr6JWKRp7cyRm4gu50PIc9CY
uMXHNHaBXoudIomWK+cv9ZrnZgWltrKthO0UGZ97JreytNib5NWa+z471uCX9ea6QIAsztxoDBNy
VfnAMfBtawyC4mv1sGagP/VbXzTHXelCTIfQOrlomWaJcVnRsvFX9yEb5v04SMTDiUwFJR3SbYIn
6fuFc+YqkEZx/GuDhQYW4DCiBTb8C9Zg3dNmLAtsiUm5w2x55Uj6T5IlzGVDHggCP0bEj25jgQNO
K9XZMqv/2Hj0tVNb8rz+2wZmLmmyRxb4il+Ev7KlRet2Bbzfh4PSzU8IYBmt9HX9SUvqeHaRxVfD
bQRCgnmSY6OiNzwoNDTy2EbTYkZNUJDC4mbgjElMGHppDsjwNuGN5wDwhwwR0iXed8SHY0ay4D4U
ldF3l1xOXsMpCWqF/zJYtjLa0xLhFqnDKQxumJgydLiJiTlgsvpxs3DV9D1pvadjq37LDgNIh6zW
k+HrdaXvwWtddvD4GlT6jBuKxTNnsW5Qmbe/pyfqzq/I83h2FdX9j/DYWbip9R3ifmiqSKzyoFCp
tCKo8mx1/BBRlH+M6J8UaiytFcxWhjTofEtvsOm2ZO6+3Mp5TzVrMWoiEiUHxG+Th+F46Y+JFtaP
UzaSTy4aTHN2jRAWvFEah/KrRmfGqAwGf4l4RsPFLIqZ33SBJXyfXQmhMaj/aSexCTs6o+aCQpNC
s+lktbR3JGgrccv/XIMawM/F8JhEP63zyZkt06NlzqcjU8sfIM16ylRZGq5iCG1L/EeT4vmyUFyk
xWmFKTUbl+eZJ/sPJ/rpPTOndX9gTLwqLZkfWZP/btgbRohkMTz72Lz6gke23ORBwkYteLkiy2md
IGUbSoc43Myy64xSTswg4O7c5UhrZGrBwnGj9IhmvBmjlkfh4h8B5aq28FutP6PXCUUX54zo+ISj
GsLF/0CJcntN0KGK9WoDJaj+uTaMiiSHDYbInwWAnH1SUWV6e97lt8rLT/GVsr35xCzinPBO6rVk
wGhyDOo7XmHWm+OkPCW0Zb2tVDAY1s1q5O+qttVGROviekTfXjOnfDkduvL9jxq2SfVhYZrE8kGg
EdYVwhxUlgoC0EsSDxPp9aZrUkC6dt664VqpvVmcMo0JS2ljU5fQzB1tbhh3FPTmx8V78c0NZCv4
MiSLlGMknQnU9P4ow+Jnu9iumI/kZVW/XgoybRZWd+yujzeQ4gmVxeag18Gx5is2pSrV/P31bGaN
822cIfBs6U4NovwTPtTeb7toYEO06L89L8O1RR3EKLqEvPKhZc6QesHPfTR5tcD1wvYDOZjptMpk
2sCeuQ9Ltht19fJwARKFgG+pOktHIkErNMjOCJ2KuBWHAe5N9/e2p7XAzfyZxKljddUim4N+KirT
AspXOf8cpYRW/woa/YUXRRSDCTFP/OMZ1PCAEuF1isfv3h+Bb17QrnbdhwJgvYPdAy2N7B1+q3RU
x8YZgoUxbazUazcXlhzBA01K5SnLJD6UAFYa6vfpwgGqyFWEgnL2LvGA4bqwo6mu7QlQokILGbIJ
ktRvqW8XlHuJKKlsnsWvU9WdbazDn3ZQbh7BX/qK5HVDHJ5G/+my880QQvgzti5PrjQ2X/MPjZmV
+xMEqqeveiRwciDjaiwA+tmjBPYQNOafV9VGVqnembPIGfZ2HVA6BX9YL4d2Wg0SUy75WDhvXqc4
dzcrpPxeVJgBJWFn28286mwqhJkrMB1KloyNKkdV/BY1IlNzhRVuFKkQul0woIBmvzbxrFsnGAhK
woArVUtZGuMji0XJnN2d8Jx3LMfxy0Mg7/wV/UPSUyAtpixRaTzAn6Cou0zwLmjbnZS4d0CxtU2D
iAMVv3SDra2Ed42ovHgS1HGmHdlvYwQEgyV/DqCvmv6tjtOwID2iVCfiwga+ZHgnxiPsoL2TLHjx
s3vowYSWxl9QzrI3qifsX3GbDJOjNphtZX1SVeedyTFEp93knGn9OGMCH7vLymORRiwfpfJ+5h/X
hBZyQX0D317DCgGJO9OmxjCOOh0keIWJv43JEyPOJnO8NfY98jrUzS3GcQ5zbQprJZTRaT60xWcE
OzkNKgaACo11lmAX6fcad8drVu1D7kzcwhUImkMTzhbZJ2d3rwxvzhJWRiyG31KA7OoHye1228f0
s9CKZYAGaVonrhpyRYiFcHjoL2J9rFdZmKVhmAPk93Ug+oxsrttqmGioO6MJRQgh7S+VsN7+Us7B
q5t8ske4F1/GVkXwG89Ia8qa2gCCZTwGXeXMYyZ9uOfY9wbL4pilBaoo1bXH4Trr8cgXeveSfOJB
Y+GEQpDcyQFIi3X4uXpyIeJ/iKJ+S3lFt1E9pfP4AYOkCvhG3/8oZSm6eMQOwxgOBZBpUvf31nvf
IV0AfljMjWWDdI3ppYz+nUsM+eah4tQnbex0eNfLtx+YbaGY3KzU6aM4+I5/yAiv5kS5QXvLpLc4
nEFx+xGWFwdihpFlEsq3wprQBWseKL+Srg9wjtCEwtiGJyAGG7dJJf7i2fH51t0URjIB3EWccty8
yVantrS/cBWdxw0YBUTcfeS8cKPNSSkDuKzEe6c1KivTyei+iZ7wQdcvZ2egEIRti0DWavUP21Wv
h8R8onee743xELNp+m8qt3yMnSIh2rTtXLPVZTSI9oq5wHPc/rL12X+MJEry3IGHwUgbXp/WvQFt
py3nZAH6HtwryMas5kA0fsn1mENs9X1pv0mDcBnXX4zCUgO3V3Nb+geDJeNFelYmMFSYtK5pupHa
HeHVvilUIqGhJuxWkYhn1wrIDGcFCB/kbVK/+ThaCrrRdXxGYCcG9DmO11cq/LHyI27evCJwlhQt
Ytr6XvvxZatDyZWd6n1SCjrjdpcaHIzXw8YiktO6Kwd1myerWyC4GClmhX4hBSrvxaCRlIzQmebX
lohvESGYCxnRzJUVe3uC2mI01sQ4A+wGUlSSp4WdU4ZAWG+EFGxHWrigCdgIoCepuI/eTLJOzAtB
GcHUp5teJUNoSewJszNNwiAeKi5YdN1teskCZYVD+aM8zJO8ta8b7UI4NJ1V6gM48LEbNaWViKQc
Q8zQuaRJybocVmpg7NpBZ+aIkKzFM6ALDPpnzqtbg44tMDRGXuqnsmxmMKKFR3vFMUx2DWt2fqBo
qIx3bD+Ym2s7vM5VODayknCOg1GT/1w9g4ni4GXQ51stNM2TJktUTFzcXt6IA+ddMW4Yl3kFgP/F
2lxBpzFvof9HmaPZMfkTOsMeF86rvGxZzLjGkiSHkOSF9emL3FTE/x5sz3vBpJtiXfwFcWUqBioQ
Bo4D6HBD3v1Zf+F5jGah0InhkDmo541e2UH7pHtaYdoVA7z/7ttTUN5tJVXjnPMdLDlvRZ3k5EwM
zyxeYgGBSNJoFiqRi1P7+lOO9zS8Z8nnENkqMoUFm7GrlBp/JhDO3PEOx2EfhojHnztOysL6C9c5
yL/QMCIv8Skdhrdjrb8gS966dGz11XCnoe+08pyOpxATB7d3qTV6SV9ciXjZy5B+K6GLOtDZmyEu
7qds6fNUy5WLZmd9RGW2hShoeM8jWEJarEFlG0BvQ27pSlGYL/p4BdOSVHduLeRp5djFZHjIdSBw
PoBevYTTOygnDjb1vxL2CURKVdY/qHQOD5JMag336MTRPyw5F4ZRHqmMDoEI8JgNDr0h97zs9Vf+
zoyxlsNMOpsWQ/PZzPBhffxtXGOgwk/lewZv1wa6MHfS08kOrxievxNQ/WYHXQfIKnE/pwnzskmr
QjT+rUqibffaje/RvWMByQudXl/NbvB1kADUNUb5JIuVNnT32gH1o1FcyOnAsCV3pBJ3ak1CWKIN
Bl7qwOpidaKIETS7nQILXTDgkrWzCVj4NTKbsvdmTAh2bLPJgoASsSInx3oaSBqeCMpKKvg3acdC
OClso9u02NygZn364J9IDg07ppJLrhL884i2AJsLv33kVpIeTrwFiBWk8D0k8MkqiriGvVCLSgdm
XBmWKUYtX7+7XYPvwCh/6QBaHqUPr/btFDP0sX2vDY5OpkAAQZXQwYH4t1apyUCLHMZtrzckUfTP
Q6ufpVZkWiE3SYd3tOmr5JkiRRUDf4q4UH2aOPAj7CxxPWc6ehLSyz3bMkRpkKEJ5Js+K6Y19KwC
JnQIo/GIB60pTjdggM7aQ3SbFU7ykJ2f2Bn/fvV4k9MGTMh/kPEh7Fytb6obNoJ2K4zv/NP0Tjyf
JpzKXaGSWe2H2/ulbLHeRmQ8PWlHJlSe7qN9/F8Y30OWv4MEhvOs5k7LxlbSe3/70uJZGzD46xej
dJ30TCZputVujfDn9DevIugLPh2TG4mu/SMCddRXNokllyuDYVYWm8wN6ZX1Z3cjClAKTa39U7w2
nleUMcdfy9vWVlpjB36iw7MGzWD/zqewwU0eCbTgZ7l36R4TGQ3OJkBU/ts8/U/5D8TrtJ0/nFCo
3CUYBKuv5VZqu0AAYkESJ8ushj3h75Z9FXmxiVYIsIXnMzikLX0b4TXhoKbehCQOgSL5Xw4vdyjF
zeubD8F7rJFGqHi/wBNpjVOa3hughMPMo03eugHXoXZmH1guCWyGGlUZLGI43wZVwOuVjgRIN1SE
L0hexzVFpluQX7MMqNRSOl3VybXrNrbi/aZKwQsAzPUBolvY4RX9VY6y8FAnZYTvQtbsa8CMx95I
qdMxR1jMoSIfgl6l3HzpmCEtHek+tlxhlsVctpmLdcUPq9/DZwNInSsCjtaBAuOaliAh0cy8R7vf
VFWZzRzk+nFWqwoXsvcEFkq9v7Tz+YHFXPWwN9EGAGh0neUrLoeKQJI0NcO5ehhmhXIW2bERWUnJ
90jOeQEk5PRx9k9qty99YildlN8R+bIIjYvkwwQ888FubEoS2xGItkafpWFgGonhGLsIlafXciBC
rKu6iZYlw2toITayHu5ZTim/q7RFFOro16/Syw9BbS2kj/F5xyGH0zXkVBT/rfy4+2XmE/ctdDJ1
FybGki2YthrgYu2XHLstBD20m8hTsvJJMlh6yT26oSJafe7+UgUQE4tnyhaz2H/PrCvRJbxUXWMn
UHxNcYtpBFSTgv5xxFKHP4ud7IZQyHVAdhwK7qPJHpUKQHrimm5wVXhU30rJR99unwrEqDMd4B5n
i18GgxBeQ1gfKAooth/QBz4cbbfIOeYiGm26EhpqS/UZ5CERtyR8MwUK8ukpRDJcgPNAa42frBzU
ORhmqE6wl6E0/dJbDoRbktSHDdcNsvaydhMTzJ9I1f+wbt2uaVmFBoXYOF1wuSuHNEU4Kpl0jIyT
PYJoE+0J6DaotlMtkYsmv+JMWpA202kFCXItXn4dyAmsNCnHItGrLF5FhGQK9uTE8SbAyPV0tsb3
QiR6p2s7PY4JNU/AqY3L4Y2SozIhFVtHxG6fJ4qsUM9hXhGik+pMlv0F7O5YtmoRWY3F1HA7P06y
GPDhzG4cRKICvYwSokbozN87LgrPd1n4wgZ8BOS1bn7J74HL2QOanDPnAKKSzLAxpUwDSCvm1chp
FQZ2dyGecKfSezHxYNu7J+Wks3NpSgCw997c1hdZCUw0FevZwISDoj8BbuzpbH7A67TgLDt/5x9E
uWo4gYW6N+TgIn8a4pTVf0CA3e74EY/yTeE63Rc3UHLJlN5MziXx4zDuB/EB7Ojam2iziPFvRmXb
Em4pl+Ds/Q24AIfpRXM5+57dHmMTGy5NGff4GzTWxnpm9H52xQVjc6BuONLKzkHOM2kFNEsblKef
qAbpk3Ct61e5iWtLfn/YwidQg8YdRamPbf1F8GPznjHehWLUqqB/F7xsZag4C8VOL64bDM2nlJh2
K7zxjB+gNCv7PNlcmEZiJRwPjcu80PI/yeb8C8zMvs4/4VNNXxK/FDduCrk/aV/JXUdj1qy9Ik7S
YNT8DarC9vTLfrVWnKmvbHCb2kIo3Jou8p+nq44p7s8/j68gzsHgadJ1xUbIV3xQpnEV3f62N6iS
s7/pZFYZZlViO20G9kvVt5srAZYz38M72Guf0SZTgVPWfGo0S6ir0Z/tx0ja9sWGL0FNI7Ka0i8z
iiZtdZdQIOgMRHnHDi4DIKyZsApZcKT9uC6WP7tqQM+M3yZEqCCjZam0kPyDUk9v50Gj64Xz9OE6
svhNDcHHzfKejai3RU45E89B7IXqEKevcLkksTBlooZaU/wPzh1JMIlqikxDe0n6Xe+TOIaf3/Sd
yrZJsa8LIeorLIjjkbf/J+uOPlZpYyDJFaQOPII1pjiZRLIaf8zfE4p5P8p7dD01dOl3FCaZ6ZoN
PUYuknrxtyLBrm+ezvN08t21QGo9drHmnzwKFtHa6j6K4jMscLkqNiQEhfgZIZnRE7yNMLIgJ+kf
ZgGPkSZLlj2OCCuAxWkVQPoHhUAhqlq4z14V1tAk1pnbh6XCcKY3Uy8DzLbKVqV4L1ASe27uQF/S
BKRZKj4EQqnCfx0Za/7+qtxkcK2qdUmLx0wAacupmOT5m8oaYRkW8Sg+kz3b60AiJswHisa1xS3S
WDX8wZGPGNLB9MVvXUFuxhEyak1mtc6kUxnT3WuAPrO/cKctjzw+4bOAL4x2nplAvCexTMw3xrZH
Vu+QjUGiVPY7Qmby6wD/xwuadNlM43siya3+mCgCqCHVjoESlZpK/g+zU0CRdD0vaQnfEBDtq4S5
ijp56SX7SeEs+M+NuFptfl3VfMD3Jk0ammotjRi6l0xHjWJMsEv47lVot1LUKsk5QSuhBPiIct+h
d2XS0Cn9QvVvL6N4Pw25Pg5WSHGyIw/m8tgw9vOL727sG8cg44jilw9Ev9BexK3RJYHgq+GZ0Ulf
xMBI5QOK4xDejcJHpOKasH7N+Uv+b7tcLihRW2hra0+WCbFvZFwYodNCeR4tNev6JMpfRI1WqGPN
wGWZsCZYparA5BYb6LV1wRcrAug+Ky4NSFaofalxPReFFYSv6MNPv0zCWJnBoPfI3g19qQQiLnU2
NW9bqIwPo16/z3Usda2ChSxcavZSOpTROvHOmuUixh7APNyKpnD9h+uORA3TlnLLPzkmyOnzF7Ju
G+jDy/Q8zrN8K84n4Uswy9NibJSK/MMNZQevzCxLhKiZWunI1CDo7DpaGpDQqBbtggdW1KQGmGq9
JVBgmRBCd5w4i09KcXu1jo8xMPK/uXYzmRJVfxKeIYiqp+iPhU2+LcM6xg6+u+5bRXoUFhyzFelL
VAKOww2V8EKhSykwfedPprhnd6UnE9ODBxW8NpvhcNC6gGa8NRBnz6bLmPE/JsvPhTuqJ6DEsYeO
+FfcTIfhJ75Ra7+qB84XLtCzIehK2bPOCuSeGonUdcYQ5N/C2TlK75AUs4UtSyz3YeTuoSs9VT0g
/JZFqw4g8zUZLqoecGv7qGhV86R/s65JJT5lvKc2IQBZZroUlyuUxphjSqB1inZ5oM77WxDCY/LI
ubtnfXtecWyeJuLMSjnqGSayS98fIcF5oKnewnDc+Uvb3wnw9qjz4jamD5JxqkGAYi6UzrFMGa+n
pzrs6Nupz2XU5RSFtIoCBHLijNXXDHsKN899XRZ+e7Z8M/GlgiAfxtDj6Ph/Zygf71KKAjDh5+B4
cxbBsy+WxtWRuFifLiMo9MS93dQBnQhndz7b0GKlH9BD2mcKu25JEhoBnJniiruh/uMs68X8ftcS
ftOIvJlyZNYoMA0dANXM44Qb7X/0zq4yrsfwmSOuvhwMLbsf8pNMtYthFtCqR0xY4gfUWFZEapiS
l0UzHsVynNbtZfNrQr4HIaXjxtYRQgyF/v8oA+i+rspE1/BH+JppZGj8/HxHw9EfbeElyKOpH+hY
7IW37VYaJve3mXA1zgizg2qMUKZTD3VXm3B3bWC8Z96FeMoMi0n1p2YYbsNS5blk4X20dpXgyotO
6DhBczd4HFCUSCw+x4Tf+9O5HPAnnGIR/SPECdNHtdYmxdQTooMj4tAZb6DPthZOIVzbnsBowdoW
E2qWRWmDtOVQGm3S05seoJfp7KxCFvAgdqF3ojbLh03V/Ubdn5Cvb6jK2yLYA3lnvpy7ziNe5/cc
8w/xlTg1GDmX36kGhzfqBoiOe+eD5F3P5M5ii0dG/G71JD+KhbGD7hqdRp5sykkrT/JklpJXtzyg
LNR0567M1JvRqz6mWW5vgFoWXmfCXt910PsPlmB9FM3EDfpzHmclq/Nj46SvXLogTJN2p2nPMZFA
/A9hM/sMPkZ/5BVxm5k7uFiCymBHlx0vGbb0sJqluFmoR+P7h4abaGrrk2j7Aq8GwbSXdD2mHiG0
Ci/M075dD1ND7N5duUA+hr++ALV98LEobLBgrZIcZWZ/CS61xQBlPUln4JN3jZnqY7XPwAIWCwfO
FeYZ2XjcK9x4gHkdfhlracP4YyBmMiipbClz20nVUMLrC2CxIFLgcZRtLWjjEYa093W/LJ9ukwNz
i8eymETUI0iZGeJ9fpJctLxhyy2h3ghPs0SYsCuu2ZO7px2bshanUB2Ps3U2SiJgNkKvpnCs2v5J
mJ/l+6KpXyCP7lNsUJLtXaidZiCFU+mbb1pVCUA3uPpYejzb8TH8f6kpoQeUR96k3uN8SdnIVZgn
wOwV57eGc+vX4YmTnGoyyIjRWyeAFcoKCWSVQ5LZKuPb2UC6OkvqgyZ5227Yo9oJM7gmWNeLGK/l
oFOxDT55gZadz1HkQjEE136yK0zn1vHoAmt/6FtWdNwAgc0ouowWpjd9Yx+1+l8MyRhV1YQVXzfD
h40IE90g8H8sWmZPpzcGvSWr5HEj1CkptNA/diTlpanwPAYV7gh4n4u5Eg1VIQaOChkeZpO4JE3h
xDQLWGzipmAfbxrSakNbHewyTN6uJtRAIWtOCNo9UZlqmBrUpUY7b/6eYHaxa777TFVFK/SW4IYy
VPUcw6+Zj2UUdqpa5puPHHHvKt4cG3jvrRVIa9mmlE0zTiaqFHs0apVeogksh72IyrgXcZNs6Caa
ZmbpDfbJkyp+WXySmavYoWJUUmpWwII6AE4rRyfmoC/hHGDKdZYBPjgZDHooYrs1EXPbOFhCbASB
fz/zDVhHyXEE++yWdJIAC+ukyIl0fKx8i6Lx3QFH66TlqAHI98adYpSCw1zQcvP9M/gWEpgivaJj
4Pg3OM9UrN/RYXEamOZzVwAXeiNux9gXXJgH0Fm1Q2jhmOxqhwWYQqxhvawtg0hahopYnmwda1lM
JPQcF8esTRuJFCn8CSvhCvPukP9wTsU8SNbseejm/n45yPbEjrsc/bSeGtUQKGif1yWHB6Ll9l9L
+VF4sAKNLYHOrhne1yce61EbhRc0s6C6oD65/0XpF/ez6L5M33e3IERlyv8/9XQsUGUznXDN7iOk
oFm00RH/JmSO4+UfGDUBvjUjJK778I2uJiztT1NRzxGOGpD90aI163bEghA/RxABzlzPlK/9cYGn
wW7uaLNlBD06tWpHBwvzvMTzslb4/wQtP/L+EM+/QGqahl3n9PKkb9k1mPqFxgGItug51NMsZw0Q
eJocBAD0vaHWL5BCwvhfKkz2/Dx/EjFxFQ679mwSrn+PXtj1DIFU1M1s+9gU+2h1VGjRWKWQ6zYn
dg3Dkj2fuj/xCuOYCUyDLCkY0xfJWdDPvkPIZg0MTWcnAzZonVsQiCE80PrlHmf4ms88XGo51DXz
gYkUhO3LKdkXmHUVzve8g6+dsOd0DrfRlfmk4ZUlBUYtoyCzOHmgN9Y9uXOWIdv4c7jRn43gJvCZ
Zd9UlUNP3DLHYN8o8J1n6fSWEi+UydP1sr0c4NISuKKMHNPZsEGQjsKq5WHVkkL+99a9DRWHxByT
maV4D8PJh37IK1o22daXQtyt8Cw/T49gY0wEmTgPDm6TlOmVfDiAbEEgR2Sh4BbVAmbKareQPO96
nd8R4hz6I6mtIL6qHM0aYW0WEf4vcLzo65PNBIDP8fRk1czYM1OhQG1kUXMi9vZIt9g/WWMPWXJr
je0jEOvhgKWN+sx0UbBVnEV+xj/A3MxX+q8cN34TvOX+RrHRnNMthWVRA32Bjn/kFbpiM9nPeixw
0w0Bk37dBPxbmjA/5jQaWdvqhV3sfAefwkSWdPtTp/BZSVxdhGzcms4G2E3GKzJz00K55C3s9w49
wqFyXu+p8Rze2c9c7zKtFpXD4wZk6aZM5JQGupnFl8xv2uK9oHr9JkMWLu+xkp+BCrt3yePUR4Nj
NlQ6vzWCYc4PwGO+lxTDWQ0kIFpXc8OAXsszNZ1c6lhMIaa/hEbi7nyh/c3TqLtoxn2ANa+ZcUlx
XcNjfZCJrEdhb6/KW28mM+22Z1w9QrFPDt5pOdzjANfdEoY/NJ64Tlft2COJGc8usHQBaeDeNlds
0+vwLKYV3mskBwxX0hHs2OmJ6Y6NgMH7yeqXVOwq14NU0p+HtqxD3O2eWSP9dNT/S+4/ZDgbfelY
8BeGLXO/TXGPwu8vmsnhXYC80uu0uvK7J9lC+OnZ0/z/9HeWpTyZLmdrT9UOCSQ8vhe4Och05G8s
pkCsXg/0uw7DhSleyPepDCndP6QA7KpJBkYnvPhPHlmp9PtM7yDEZHtghcEn+l4Ex3xpJjWQjUl/
I4FfDMZdWfPj3AiQhMSwoAt1vnjNK2EXLBhLxcPff3jrFB+tYJB3V2dA2A9DDNgZjWNkfKZzVMyA
t91lRQb6acATmyA6B2pR0xEHMBSB9UbIkSXeH9vTSDaPMrU1ftkGlR7DJj4MMDkG28zDXKHuub8X
iwC7N9xDefbroWl+hjOekWTEL2xDtZzb3x6yl8b4lIPIPmshSMC0mIs9yij39dcX6J9Knliz+6ym
5dX7N0qEJNiDnndG57uJNIkkisNTySHM/3D8PX5aZZO4N3CHrkswJu+MROIq3VEJafZHj5E8VreQ
6mLY9s6cCI09knmDyNLakX/Q5BdkDNvmrkd5b+NDeWlCJdsP/y2XdTKMn2MJzz/FNuRZ4uZNcefT
N9XZVKk8/U5MyBFZPo9kDDD1cMtF9PiU3KVF5hKDA2LWOJYtSJXZJoOFDdXXQ0MGCJTCAC02+5cc
048CyAc+C3y/HHT8nt4Byr3NMRUREJz81iGk6+1ULNOYsTmVshp9gzMFZUaLut+AyjDg6L6Pv4cw
wFF0cr7cP9pPY/DiDkgLj30E2WbrfbX5n3bRW/EveHpknwZgSJ1wMoY1lnRJzcwfqI88aEgiAne6
KfnwupCAYFGIxZsugz8oeOXduL1R3VKgPfynOuUPXM2Xi8zN8RSQC/RfNWET0c6JOhiKXBhpwJ1W
MBOFLMyAsmRaIBGBKTEikGlDA8SF84JqUJ2hNCZ8X0rp58kc3IilgBvFyUj44nzIrPSDvj4wD+UE
wDsp2/N+4q0T8PLsZbVmoPIMu6fK9FWBY4P6LZrUDNZq1Rzp5fyhhG1/Afu50aDi0tiqs93jdsq2
vePp3ViCHAyAW1+5kMOtuogVH9zklPZClJJBVUn7AddtyAkIqQiB4pmymg9KpOZjwYe3VMUrk/R2
NsCMWmPvVBk+j2zIUg/Q03liGplVKbKPDu9iBGSOK9SAsjWsgZnLsiZ0NYiBRMhot35PiI2gbHfG
e2Gv2OO/XJ4Wnl/z5Ie5CTqZ9GkctYscPhnn6/ExdkCjeL7alEdahMqj9AZhn4q05k//Cd+EWEaW
NTjAmkTTwcLcZV7fh+rSHR3+VGIWLM9lHDDDzrqmocY9odULSnMEhZWvmjfB87lRJb/U4HdwWgld
XfBTKUc7t2y7SQz6KmEww0quW+rNtrqQ0SC2YuZX3JyjURQ5W9H4AJf1arO09NCI4fNQyNjCJrcN
OQBYyIwX/oL15dKPlxb9njExhNXny8go45wrvDW156tkrrcwzDKN8D87A6gGvxy+piYVLfd4Pl47
QS1cu/CbSxM3dtApM7Ipv+f/Nsnbs8syuoIGJpGVGqlDYr1pDBms7KESrTSoKnm5wdAYwN56u3F6
uE88BA4Bfjk+wt16Aj4isn52vKiTjMCCXQpVstLkpklhE4KIMZB/WVyqgdPYHNhKJM1wAAR2PHf7
GsTPJVi6onJKRkkglkpuJqUyBDSRS0QejN/2VkIrVwilBKZhKdsVJHP21xqbZ1k5hrDcmluqI8SU
MJLoZp1/X8sakRA1WeBjalq3z18JWdq1doesOCbjGOEhsK7aKSCYDO2KeK6Q1HW5tcY+Tpw+0lt6
vcIoopn637ZrshC/rh7/u84k9aAKLn0mdSyINUArW/p7idpfyuSVNDYuLvCeVh63q0maYHNnppFG
2JgsgmBJ3pkgLVuVhwvHEmBJFd6WK0MkgD+/2hXjcXxSD0i7QDywUzFPVQ2npuP+mq3Nr5S+yRlf
GDga9C2yRh1F3g5/8WiTcZ7GDJetOy1DnefJEr8KIGnR0EWKp5MZI575+IBAYxPRv8doaVe5WNrJ
CtRIfzYEo9Fh29uxjptxaRrwlWR0Ufht3MRczujgwLq+fUm635nuJz2ijHdNBrjtjtihEa/rzf56
6sjkPQNqEq6ZedsyrPsB/36eBf1xjSmpinTmeA4SRWKDKXS+qPZSV+G14dg5B8z5XzDlkgAMgNKf
s5UVaz/4QXnhkUCyt+TofEWK2Xyz4/x5ZrG8YNz9ac6eYMIyCxIJt5mqLlxHdy2PQPIJyBFkJK1s
8+oRiwymZTcDf47T6eF6lSfLGxrYxXdO0fa4/F6ATag9v0e8tPyW1PVIJW6HZflZS8HzX5khpzmG
0ZjWs8ztVoKLZmGQ30fcPbtNCpp6hC+tnqClvh6IHl1SYHTVvAaXKd/VCCHzJ5q5ZzPVAtm779S+
hI+g54kkaTHuKevYBiDoGCp1TIy6bbmcpyAdvcxsGJ2Ak0cpJ92u/7R6CmvoWPoII6FNZaA0HxFI
jIVuN0lO/4X2XN6N/HOy88XSo8oAE7gEyQvDVYFO11G3ZEcMd0FMH1vXCUVZBRe1u7FhNIS8WxQS
qFL1Qf88uj4NkanRrFFqWOFGV90eorTdmUlIu2aextbHpd2Uiom6ds1cgfCg0F/8tW2o6ZvKo7iW
ZmSduFLTLmX8t+JJ5qN9cXuBMuLJoYWbVe6x9NJYzlgJhyIRs1tr9QSkfHy3rj5+Vq+UB1LvBzzW
ac2gUhBswIVJCsra8ToRSYUdzOfsB+ea6KmtyxPNBpqt3X3xTn9zZDP4wWs338OFamqz/44bZRTy
qIhDFzwbePnMYjxTM6Vmv/xU/al7wMw+s4yTwUrd9yD3XZor6FGBvp99NDWUKIf07SK+vrj88K7J
GYGnHUc1jdypotr2oW5Gpjy78WmdbMfUVJdTDUDlyTKPksP3OR6EYqYquP5f+XPoPTOQ37RQWIiR
TY7T5Pc+YZkVv1RVqxOvsOOyyXJARog6w0EFxBonjOrTE1JfAqWaCsQPz5MbjaEE71hnKAV/Vn5O
pdTQif8rTsc01dNqLZU8cYDAql1YP3iBKkU6IZbRS0vggYCpAv6PKZfEIZ+wj7D24nrN+QmKrXWP
jxOmljEnvd8lxEBjbXf1PRKDrutejUzRxu3idqhL83FD4DAx0ghN1x4TDFMJLDIwXJ2zos4PQKKb
fordf1w8rjc4baGoFdKaBFqr862P8Q10PmbbGoFULoJSo4dwebCxLIeVwM4l6IBbNJOaIM5JkEiT
sPRAKCcetEBIiAukE03S3vOOWbR458hHWznhoN5GLwmsZ1waH0eqLUsbJ+RVmeY3ZBvzl3jGDshN
oTKnZMpee7t4HdTXC6m1oL0HGNne6HklDjgm/fvY/h0szs6KtOIqxInGRZRg8baABEnQVnE5Nmf4
JushdPIOB1EYUfmHMRxc6inSuZjpvO9SJsUYNCS29QjX9BJANQEb+wcx90FUJ1Py+laWl/T538ae
zC+9eMYs+7CYPPwE8Lo+LjN9tUBZw1FHIm/n5olgzhNLqKhSA8U+JEhcJ7uYDkjfmc1XPkicj4am
yewUuoe8XByIfkuQPZcaF7/4Fp871IgfSqY5VIu7zCLQZs4vnRfSiu9Sh160mL7gbVocqP55v155
0miA3u79xwR79E+EuQGLi4qubXXGHdV+b1iu6Qsvuk7f7u+7CG5+ijik7WbWOBt0vID19LY6GKuD
dPTX4gVbFXQ/oIKvszWrFMmkwfElyWyAAyI/2qSbPqQMTbrAjLiby7gMByuKllzdv1OSevdLBGdd
gL+YdIvCeiTe60fkfjHpS1PkMJ70FR2sdHEsHqpB2unapJL+9oQd4lV6GEjbo7LXOCL8AV0faN61
67e5rGMQVnDVr9v35p4zVVPZJqzGDXZV2O+xveiwPtRXaEER6vEzCMqcdUZxJGSSOm5S64s7NENi
bpBky5Zr9izGFewddfwiAJNaji0Ug0vyoUITKM6GP467iC10c7RLyBsgMRkDMbDaPHI182pXp4TT
ufbERUwd98+IoqNmIx5mZn6IcHiHlWLKmPMs6+BC1+/Qtrp6hEk1IJFMCscdvEep3UeAH2aqTSJj
lnBB4fEDRrnh2qqKcR2C6OS2I0uBwrUn45G/s33Hk5DM8erM1qQRGKZD4k4Pev8oz3dw7/MyTF8u
05EAoQ7Ti7UjBK8rukva1KA9MHoprFX21H2Er4Ip3Uvba0dcRhcxOS0UYzXKltCYx6nLi9cCwaMd
oExzETouNWO7a9TN1MUVOeMJfhMGC15s79VmtG2eol6x/G4c/J0opkWCeadfkHDRH1u/VMgmJ1/2
ygEO1ore8PyR17+HogFqYduUBuj7ZL4VT45+uxClZ6zM87ci3/b+lPt1qsfjlxtgpioCkTYcNZB0
Ed1Ynb5qOkPUI1gK3bEgckCiO0sIYEiK0qQfgu1TMU7iXte6sFOqAu391vUiHQIVMlKJ6jmIeSQu
dbg6KveBDY0u/eawiLFZVYvucuNR/Fs9b5GczWLLbQs2nWx82Ni9Ngty9CVlJhQNvPpWD1ssWvkD
jtIdv1ldxEdPu+2tKdgNrXgkRDNbOfRY+jxQVRqunfo9uHo3GqeoCYcagYx9aXIzgq/eL8Ey+yD9
XmvkzBNiccOSuH0UTzN+fCiBZmWbxwHG1Ud+sAY0eN5/NcPG9rYAxuP4xQPPdStlOZeIzm/WL4bM
V1IDECewKbmZT3nIQF5B+NEtiPgubRDQ6LWqQaVctkHCzA6EN6vP6vtEu8GMHAO1smFr8rmQvUdJ
o73OPl2ud1i/HHl9cmpEMTtC4d+CyGCsg4cFslpCAwLgkcVwdkoZkKshKL4A6VSJt+gSeuKE976h
pzwb1VsA317RSdiZcLd02dKLT7rlaeNaANsve2Tqlra5fOLUu9mpB2XmKmU3U9YytfOhPsDc35BN
h3EON7tsoHK/TxmPtr5vevFLtELvK1+SjVVT67XhvYwjeb4Z+oEFCx/rSRohB0KFAvcLeDdHVlSG
N5sexTpogbywY3zT57/vZ1rUdWikI313416f9ST7TW0VqlBjLYWbjijmV0wdUlErB/hkz3R2Eftr
1hWkUJbEuDkFOkws/LX0Zq0lOs/R3Jb85PDPH/GKkNsgjHdsuUWMQpVjK9++f7mdpAuLOOxrbJgg
iBtfvPOShq6WGZdXskmzroy0dAfd2mPvVtKNdjotM/DiUMP0pZ6AUUmFU1Mf4O5K/55L9cRjH+RF
XzLU6eI/hQ+D3YYPbzlpUJsac4mx8FPHST057iwdpkmSCcNMTsXriIB3upOxK94U27SfCaTbf6P4
/uFrXB9zDkF2bMJxqKW193oiCIK4HXNhJwhXTz+f40RJNB+bIz0Y3ZXRYn/mx6zZI8V/NOX6sH60
E6e99APnwTmrGM16WeTBNuNlm3s4fJVCskqHsKzbR/SMYwkbBKi8bjzmKDOcljh9ymUYEgb2PWXv
kU04oaKdXOE9HW/LS7DB/J3TwPL8KNxHb0a6/h0gMCKSRtZ+CVPB2ZHIAxJPu4gKflRpXAhY5+V9
JEh8akefu6QWG7PB/dIDE+OBbWxUV521XhpOsMb4hmtB5OMWxPxBA7wAA2w5ePyLVG5Rtk6+pGIM
znNdzLBF00ekgHTCAyTfFYkX2a0KQHR6Y4GkDiuGctjXSGyGXDmhphD5bt8UdTla5ltL2DI8o8k3
USXIQvZG+eKB4TM96FQ8CwMcyJ6yCIj6GJTHWEH50k+Jokx95A1flg7lQy3OlaSZe13jS+YpavdF
iaUutRlXc7fY2KcNJEnFmt6/10IQmVfNmuGhS/0FTao1n8pzf2KChahZmVvuEb25ae5psvv5otSY
9+wVfMjsa4V96Ic8YCC88a8cyg1OlJLgDmEtbxloskbVuEx39F600mg+Y39igmFHz+T/nFB0wyHG
l0QojOf7fu2DmOBrIeyryD74Dy02YuroEb56h1pEhEsMMKeB7im5RIBcaIcuXg9K/7J2guvER8gK
vo4HWWitb/MgpdonRblZNxOHuYb4QGle3Stz7bVLFj/a+Uzskms5K20VYB7Dfr2aLj/ckdyJljQW
kbe8ZVUlbAVNZVMi+WVR/l95PYRiJqZWxyha8/ik9uNURUWHeAfzsowppyMALD4DgVeoFCiRpcps
OGYsaqlrfkS2C4FL8BkJ+ijvWjGVkS6B76inbYukchn1ird1nSO4Fi+jUICZJ0fMGAdYT96Vzwiw
NdN36ZnhRBjrzcp8378tS1s1/eNAzzcgof+way3R67v8CwEnfn28/aZgAfmtReoYkL+uCxQeInv/
Q/QdDzUjQxHwL+ZZObSvficgr48nHU0TeGUFeIdRFZJ3yqxNvo8xBMA8hyH+trn+NhlsBL9DJzrW
FDyo6ZPEUbANk++LMA77O86wGLrRyVgPPfOp9hWIk89heBhsJkdokEU50omS2rPU/HrAPiVeyzLK
R+cHpvAWFePqG7FUAd2+Ee+LdPCY8xyE3KKYgOJbh9PsERCkyIZXIxqi0C33s1X9AdvjG3Y9mVkk
DZTocr7SHsCB3akRKAzFJQNfCBo08Z+NONjaS0r5QpJeLPeCfDb52xpn5HJBtYBAL/xqJo+s7xI2
wuxX0PVG0x82YnZnMeVIagqV+s/zY0VHr3yQBRenFriIruPhcpSZTG1jXFy72WMTvsgtdh9ERaRc
iBHMPyxnJCjPwkH42g9QNdmSjYXs1fcK79XPW7SmrZhMF5HL193M2g+zU96CYYRRdQPwxWVoHbjI
wFJ5zHNrwMLK7ayNrTY1W0GjiWMJMrQf2ufrNrzEKr0fjG/GnMW0Q0vMeCUaek/ZbKkV1OwbI9zh
WIF2fKNghsEo4aAyImXvhzxqF8u1Jm/WFHiEcuqFFmxo2x2dbvEGlm+A2KDODXHU1dKPS0DF6h2J
2eyJLqoQzi5eKdEIbEG2Op92sES6pPwSfR5eF83rLyyM8c59GfS5U3aLM+yLkEF/yfzov7EH31Si
RaStONQhGFJJTarcPK3fUD7OFQBJyuNQA4Fup0GISi4ROX/Mb2DObyJWoM9gKtHhtzYhEZVoYpfP
kc/YwptfDzhyGEV/htxpgQg6T4pAsPmiAQbNsjV34smlJp8LMCS4FI/28lRgq61Up4XPiJpJRZ/p
vo1VNc6TXPvNoHVLT0sq+lXimq4LJ5pyssApeA3NSDp5a6KxvtdBn91uKqjlo6LPBv6ZL+oVzP1G
g1akQwcFO1/mAY1wa0OP5kYY0PgzumCnUfAiqHamwEUpKWpBemJ3w0i8QIF2ZWo8kKGQdADeJKXU
4RBinev/xVqdDI71+ek9ta+BadWvkOLa6vYPafPaLCHtlxj5GRMLI9cIBH6jVdypSnVwE5hRChHr
GY2bDfJDGRsv2OuKgK2upWF2kjObgSDDfwA4nTB35ZH8z3etQY5gvzCaLbAoF/TKw9Awq06Kwekn
XpcXonJ4J/0zF1LEkj5++TkVtwllSyuOrs8Jo9UYfpEEFTxEWYJQz6l2KEGyANF35vGU3qEK5EA7
wS4b1i4uyw9ckYCwjNHW4ApI8eDAA85a8/GsA8IJIZB0ms3fPPrC2vl/0FeyS7Cww0wtLmmxTq5Y
2iEiSti1AfOWpvmpRaqpvxbOMIUQoDvroU7pShZXLtnfkmx9Kl4Xn6CouA5YDurQaVLeAzFNtUfv
iQidnocQuDJzf4qZcPmr1Z70NnMmQU2PPnWJjn91XEKaSSeS/1xRZ1HstPOWXmiKdqBLHm6VwgEs
9wL0HqyMzvhWczNotKtrmbFj4xGCXLokjYkHoZSJgWn8khtbfl4pm3PsnKyIGrK0T+I/b3c7/Etd
MC1uaiq7aVwqJQSoWYVP6E+A4FHCAeZnGyp0t+x/8Mh8YXFSBaThdYyAY51oS/v6F3X2iAWR3v+3
vmAl00eynVJUzBr4IT2m6lzPKkmIa0xWnF0fw7am/9mTVdldw8+j+yoOp8wqCeeNCLdiSgaFl3Y/
EBQheG5ER3hmQHl/UdAvjllbKWZvsSr4brlgPvTWLckyE8sUaScVf/6r80g0eTtTMHwHOv288pY7
q9yBwY/pA8p28LPvIbrRt2GmqeBKsVVzhtDpccnXx7i26kcSdpU52yBvRpbQEBL8aw5/eYyLiaBt
s4okq8GgVIRM+7uq6YBh0FWliIGPxnacq4Dsz7C63jZBcA7IWfU3Ec0DIp/JC4eF8qrzUaXk1nrs
9XF4kFkswnKwTvUQ6ZsnKQt+1yxgHl5D6Jzx7/JdEp+Ee7w50qmjWwgLH23qVc8WlSYqDR3Yl92O
hdwkCvYfSn3kUj1AlHOeV7U2PjjpmusaALS1IRO24M6P8aIV5Lpw/4LF3adSkT7sWxVpJ4r+siZ9
UI28T/QxCu6t9WXP+6w0sGAfsbyx3dnS2jzcEUC2wAntxX21LIqMp5aoyeAVKZMUCVK/K+1L+UOB
mQXGOMOLqWqdgtOa62ukkBjjOBtvPweeLsDWM3Xza8pfD8xng3+wgFEEcEoVZ1t6yb/G0rtmbs+y
wlTesyprMwEYPfM+bAQoAC28f4Gy0NxCnG4GIfQ2bUl8yj9vwr8PmKx/jzjahlNkJx7QZ1XmQrRQ
pm+Thh2ZpkX2lU+Od7z1++bnGVKUurcb61pi6z13BguDMV7NgIl0PsM028SGSWgCMP07ckR9QGWD
AKRRGvgYFqdmESUwCpeT8bZZoLoO8/rHWPMdFeqr59fjLZoGy/3CL+SJwILXvfgWmdOwEVnkycWb
TQRDhpKUUx5pUFVoivj2yCUpYdJkszh62Gl5Eqhcn1pUnO4toST4A4CDmmBBdeunF4+D0HjoBor9
ZSYsqaeTjvO0TEhKy+ckjoZ/+WuPDEMNONcWQ4voM4Fi9sbAcBsjL39W9IceKZZ1tFZ9Nur3kZzV
7BKAbmnKmoODHE6Egvhh8KyinlU5cklPq3NW/gcQGOueXbv6KkbmifoMo2ZCcQQq3ULGjDAXKOgv
O2Bjd5o5nVq/aU1rmZ9elHqwJTSH7GAi7EuP3Gs3uaz+bIOM/b7V/zeY5bvWJipFrQcw84GMozSb
EYjIGmnNGR6lhjm8sHDFRuy2BJwYJzZJhhJ2z3Y9XEznBj4N6/c4IVc+lL2x+y5LJBd/Jnwl9165
lWZ/mG1ny3KqSbx/b47sRgVoN56J7jFK7qY0mFZBypBNczz+Ud1N3HpvbuNHxG69rS4xAZ1HLk9W
pIUMA4kGuuhDVWtWOaQE1pQVUHbtey+5qnWM8WIXHcn6sYHAYjabhSymVaX8edqzusdjYwJxiseK
UJB7fAVNZVAs3me56cn8gUFYlfTkU1sweL2+L8hXOR2Y0hu6WM3Hg0WDuKz6pYV1E5kf1DBXXTyo
8RDZ7vewHHtNl/QK4MPnzCy5PVF9qgRK6wy6CalnUWTj3u/XeAOnXmNweo7qYLM28rmRSdl6gorH
Y14yOVuKXco+HJvg/wKXPHRnzlnTHJDnpAMCHNsNW/kcFH2ss/wRuk7pRuR6sYa3JwVoWT1qaWeP
Wyw+ysOsodSR54VdnX8kN7lJG/LcZLqVeIciVinIxAWDwYRoe1FsVINFZf3h1zzYd7M7MF9V8/uD
H8mDawXk+HDeJCSEs/1pKmlAE88YOHxxLASGR463mKpC8Y+dogvnCpAC0/4xXL0W3zh/W2VhJur/
CsdTgNOVTwNEANaG02oHduRDRCqqQU9gXoP3LHUZCgYrWxD5r7ix59n9VCCHR72X55qhv+WTkEl1
HeK65aI8wNrJ8VjZQyDEVeeK4oRwi6ehQo+seobe8PLCYe3QYfFpL+12cxlOZiSAiAKhCOQMT5Y0
qAfdmDFimtwr6qHnSegLNFtspbHsUROH+Vdjl9WLLUl4gcmTOX7Ni/Y1/uQbtjts/86rB6foCZSb
22asCo+YoIxjyvHIcoTQBz9q+WCWJbbCGxPkZmy+loFPepUfkubezfIIcifVx6u7P0ez1/gwY3ur
YXpT7CzVmV5joeFX9ewnuO1djrChVZq7cPx8xYBPCVkcmAb3IDTRoMqscVnF3lyhRSMEStAyJPiy
hGAdtGvIvkXTQ5WXWpbfzamh+gR07+G9yNxq44p5NYxwxY6a+gMi+UOyijDMFMhZ7ACQ1euRXDFk
IndGWJx8YrfAnsiINwYLKmC+GP+d8Vetfhp0YXX8XAmQmHTggUg09ER2js1CNEMMjJ44IOGTG0O3
8Th2/UG3gzBBg3T3QUv6SrsozAJ8YLmmTCievTD8/kWe5n/efWJ1z+L7Wm1FqABHz6xjd3da9eTP
Hf7XiRjNHV00ZoZ9eBnDVk3oH7MoAUEhk2gtvKykXouaUCEyJQRwDqIi2hnH7UfTIxEY7UzCY0rK
pH/2S2ltGqUNO/MHKkxVXi79xEeT3MbZ/qesuCwRyF6qTQGN1pGD99V4XxBWa0MsmTp5fNEm5mcs
BdsVKzDovpAY2iMpOVzzMHcgFtyyPv0wiYWxsFHr5ZZ4Ha/SmFnvCUDT79FTiGSTNkils6Cuy82M
HFx2nhaPUifyNM9FIfh0/iSomWRXl9mImdhpniZhj4kDaPClfZp3rB9diBo/q/iOQ54ylou1Uz6/
fGrCmVMjQdbNUJdWa8yNrjgEvvypBrAu9wXaEx/k4uy1G8HdDbhagXX8DR/eEoBDNjLcoi8UR3PR
oSR3byE4pr7KDsfMpallqh0r2t87HvsfVekmZDD42WWGJXx0NPJpy+GptxQjGGaO9CKWs4f1Go9X
/YcntWCvz1Xugmp5GThxjRuf+dOVJDGJNER2BkgDVdr5owNRxeK0DXwLgGvjIM6ATiJgbCbElidH
UxGfQ9TUA7k1RjxNR6Zbsc0Zpt29pg/RgaqugB9iW7DStwdR40Hvp63ntzQM5jWZMuYM1n3CqCYR
0U5kTPy42LdAv+5O3y3ZHSNE7UX0wsxmjPCiN5Kt57Gbc91SQlC2Tw8MJD2vLTFMox2utbn0R9Rm
QAunsQ2VSrPH/0sbxNKNViMfKG7qj0GYw+Zlo3P2pnvj73DdiO9LF0adF66MNkcQZm9qUYXjZXU9
P1w9c/cQ2O9KpEpZedG+h8+nXrlVeAbYF5tAG3dx+XbKmjFfjva7/oTBubBP396BHGiZA7F6Xs7S
D6KbmTF3tmIkUZ/BhGPuOlBnlmInm0krUaEmfPhrV2FKbrEWq02O1R3x/D54Phb4n136MqL8D3N2
kkqJSweaMgLSjg8huJtC1QXonu7ft9MyYpHXYCjwt2AuQb05nxmar0S4YV5W7ydo7yJ1lXrNzZMR
iQ8HMuIEPSv5SQxEHqTS0EdKR3NN6wwzYEWMpMIrMpdIcdy42a5BVuH0mguXSIa22eCtPrJBDgmZ
8GaCM9BpHyCyN0nCGOdGNop8tT6SXWSPWpQOo9V68XTDMw0884CpSWAejo8tOjaBdKT1ZaHSlPvp
BW6KEiEdiNTpdbiS0baB5AZfld6+4LzTtz84lexjaWKHOnWnXqlOSRKa6XMwVyGrE8qPo95clpFC
DhlfO5hRMSwWJy/fqhLUCJCZEsaet9aqsRqXVSLZIsUfb5CL2jOZt/7QR7mm1ROPbeyI/siK5a+S
WNBMN7l7wkhr+6k+w6vrlALQherMsLXdCQsRjYEDHu+h5bbSSQoq4q+U56jMcmaIJ6YszZaOQzlZ
sfgJC3f/6Eh3M1znnC3y25vUySxxWRHEHHz1QlNpEL1Qvm/bM7lTkfLTM4+mUWhKwzAG3qFFyVNp
hI32IlG0x+nUIykxI+qclKeNuCKI3SKag/2XwtCPLJLLhU/XX7OcyNxfLkl7J2PeJSiKzf1Jtdnk
aYzVhn8eb1li1DD2WBb6nJmivCWGbJnoXYFcY39YLThnT01bIBlJGwfQ2HcUqR3zeJNFK0OOdOSF
4QJWU7c7lfs0wpUhrnSBRXRNUj9z8BFAU0/c2bKYWezGgOCb/8wcXkk0ozzhfPQ+e1sDgeTCrCwX
5f4bLwc01+xsM68mxus7V0RSjQbvm5lQyAEX5JPUaTXUCWSTf0LpxwNJxVDtA/Rfu7CmOAi16Lw1
aBbBfgkPUuvRMKboBUt6YqIECIUU/iTrDaXZheWBcwFGtTSayJ4mJHOK+dSwr9HNyn52SI1VI3Ym
gqCrusWM0G+b5Sak5lH2v3pjSiCw8QAEjKmWMaOE5w18pShqusiFzutGp9R/ln9AzvlMe/k3xdUp
LFGJOMYiYCxC4sEYdbFdiGiRjDUj4vfAxD+1rJjJ9M3s9VLicE6LPvMbxiy4LNfBIRjnmJhPfR5P
s4AxANHVS57uzfgBfd1XdGfOHufpEINz0XOEIr65D8SpJtpnQBcpMOxStidTGE2LjBgspadLw8Md
jDnwhB9HnW9/rAySS8RZDPSlpTgxVOluA/MWTgCggos/t3wlC8Kw7E+90lW1CqSY+PYfzHqTo6vs
O/pmiA7tDk2YbPvLESTpV5XcPY0Qfx11SJwSsQnXb62bcci2A2/GbH3TctapYVWLnW41XTScsOVh
0LbN1TqXYgFZ413pdJOahrB8xUbGERcosr8nxMzm9S5BSWa/fwNxzA86v3V52a3sGbDA0MFJD2XC
/RRYM99R3/sGEy9pEW7atttUs3QqMasBNMv8EduHghseFAgNGbbwPv5o9dNdUDdnSDT4B800/bMX
vtEKwlLdt7y5LrkjaysWkypnrYkpVXy4vDSJvpAAWtO8SyXnRc3kG0IvEsBQv5MKswGeWf0C1a3S
dtYpVemrhzyLhziT/Z7o5BpN9DMNRwEj7P0ZLE6UQt8Qi/KfuLaUoRzGZzUVbVeKZTPULMVdNQ7M
wIkQTYiOIAl3HT5xZtC9NMCdHcB/3ewJEB/7GZR5zeOr6MlYSXGJoD9l8VOxbwSFWUTja9qsCeX4
7zDcAkAOVc9qNfA0sHJdI22CjP10Nc08WtWNjtdp9eTU9eOwekBZZMPX62DV8YpRj/7wa6pnDhbt
XRcwl1c5U83rpJBjscJTMUlj80ujVimzLKoP1aqfXdSOS32wrGLWK3/yAIXRzaXg9tGT7lUrFbuC
ueWGfWYYR91old7CoqrTQ/50u/E5MdTv3Z941VieekqHBYaC+BBBI1xEvF7FaHOQ90PqZJYS0syz
6s0Ltu1vjSTigSyVsQBR6QphAzfcIJ1JPki4UmVORIQF4wZOBIJ+ZC95mrjewZCdDsVRm084ycig
EeVbUb9HENIKlbuDF9Zr9VuvQaK4JH360xuxPTysp4doCZHHBQJsy9YHpi0fsqMD0mHaI2oUIvxD
56Pa5yS+6FzGZ/cZ5pu+uLTZFZrrj/ciVKC/pOokjXmCs6xwkAPbQhwQqMl9qWPELaUE+n7+jHZ5
7cTRa90oz0FL+XNBHfxpZNMpOBnMduy9z5goRnzlAfiQIN3IjmNWqSVuU+HaiycUApp74Ya69pyE
uPqmS2l7f3wuGKu5gGAC/Yb5ReSg/TTWWYWu003ZaiSD8dBSG8SCP2svETGt67ZCohG8EixR7Svv
Y+6sN0+9w9+w3aXiVFJG6kBWPOOEx5ym1jzddwqAnLFts7DHzUPVICIRAlBuRza5eN52PWSB7quJ
wKLTL1r/ilGOjw4+B5YB3G97RRcXv7Z/1IVlnd5orLdhsYZ8hVbS5iYUCa7cgYfmE0do9HaTiqNW
ZXu6NvlbcIdnCAN6T5Iis4DA2tXs+zgzHFuc332/pWiH7RRINAMOAgUJ2U5gUp/FQg2x4NYzZNEm
RVBGVFHRVlSxITtFnGop8ZGsw/xMNk7deD/KTk/ACFVatrBeMqffqGgx1HMXZUF8jFrzEnkUIuYY
ngIr/w5Jo4VxLgTs0S6bwVeQBoFM+nLLLmojA/h+dAtu3S2i6ADJZjg8pkUqBn53ZuToVCDlu01d
SBNqZ+w6p/Vb3c+PuOdbyAy6l3vdlvBWZmGi9bOonGJDbhujbuRU51UeAJquWPIF9/m7PrE9P91S
jAJ1nLh2eouq+C9UZvoF+idmBkE/EsWrlgK20HB6esFGTOVS5fOZkYetBbBJd8wuE/p9tyHzbCvc
cI8bWonXeRa6MIvdFogmo2BWBO/ncgfM/sMy3K2AqBslpyZRhHYu92kYxy2rsHFZGvrSLHYCNZ75
X4iaYVLJdt3bXvqM0jKIo04B33V1uvb+3rc9EhNPo1NHrYhKPJmKyi9fbGJTUIMbLbV3W/nyzLyd
aRVHUFQGG/nPv0kpjH5CCXgNt+HWTPx3qPthpYpxBo+iFXI0NfJkcTJK2UFGO3TY7Rp4M2etxHNw
pisOTO4abRDx7Iq+Svr5om+U0+p1guQpjIe9X6W2QgxVC6wCQwIhuXmX5SJ6BnS/obDiJ6tHu7gO
P8vpFy5ybS+gQThWtHPw7WC+RU671E3cgJ62GnvmtBTcpIOt0zIkC/CT3Y0WJGR7LPXNgBXlXrFW
9LfgGIuTypjZUzfAH4c8z1KnKQ/Oq6ufGjtxGsfDdZ53XTc2uaveqHzbdZeq3+Sxx8kHoLLH2kWl
vm/nJov0OZ4cch9iOiDwICuuLkuwzx6+DiPnh1gPe2f0hX+B7XQ2SRcUoUNu2nRwpENRK4fiJ5VH
Ub2gXImWIS/55CqMmpHfjaaUu85ErB15GXOFjIKdHaUHKZm7Irb6hS3R8duULh3q+QSlPC60/beN
KGCbNweZYZZmzjvk7XDvIzeGYS59Myhm1mVpotSj+cOxIZH+429n466lQFlOl5j96/hWi36RD+Ro
1aqlgQwu9P4PcwMMy55Jwrl27mXTCVHlgOESmDRntw2t14Uy7RovDKZoCVJ1WRMWqMnGFFt5Cwgy
16LurAyUjJHefG/sif/bP9bgswOCVPk0Rjivj35YmwAx7pnW3uQ9JFw4K0sRwvN/olw+olE0BKcY
0S0qNO9Yhpxzc9M318hOitHoEF9x7oXoGC4wYeX39sqzi2j3yNQhPUiXrE1oVwYoWXQaVBq2t2/h
R/ljLFjGLt62Rrll1XsTPJyzeeLIKXZcgk3f20I1k/dMEs7R3gU4hhrE+kNWaIItF9+d7pB9lHjy
mYF5hiuNukULx7OolOdCwuM3V7PXVFEN6CJQFnWxASJYIYYsT/BkqHhkrGXTim3s3UODGoVpZzQj
SFhYoBPr5i0Wj/zqMINb5v6dvco/MT2jPyaQYvwR5lAvYXVIdJWDqbBdei42tYCrOLAZaxvkb+Rd
37eBG18bwzjm1F2DX4spbzOgDmxQvvNoTmH8d4+xGw+NxyOXGyBx0DEzDk0Qlg25xAawgEIuCozW
MQzSaZhSJCrA1Q9KokIKyP2z2akhdlMlPybTleHY4hbR42F9TzO0CSbgUziBo+sov95xnEnxsjp+
mciklsHX7+FjOOHl4oga0KdRFEclLruy39C24ohRb/jwIUw24nwYKXat7I+vWOcY/LCuNXp6396H
7TdPcZgf7yRVximkLlpvRcjgPMV3Snl1b+z/3R65nQ6N7uP9pIcYCwsEm3HtIWtdt6Znm4HRCRQG
wochRtvbVE7jHd/ervynYS33Y9exKVnENd8ylHaMIW2HKlEYvLmHCnWqDAsqhurvr4nbYsxu8NSd
TGHXiHDOGekFP04BRU7EU78SN1JUQqlDR5QtOMFwUmoAE8T4KIuGxGvjUccsD/z0ySmEJCL71wyT
QmfbfwLtpOxXJMh4qTBiL8/G+F5ApkqSrTNsVfv8B4arRjDrUNvOGVuz1WgS56nMJISIq+DfKF3s
fVSJbeefNv2Sv5GBjEzWAQxKDVLR1ZRjOyZhAb/+pNoCVh8Hh57CvScXQiTaC5ZfCFN7QlEUlZNr
ToTkArLu2GJ85u+Hx6rfwcm4t4ltf4ky5f4k7guyRaQRxhZNiIkiV5zMiq2kujajaEjBCabXpJce
U87/Mh2sTzpEQn0FTr53YuVkJDziZ50yf+OYOL33E/jOU0H4TYJlXFPic+q37yZWWnuYY2y5UNZ8
Cdggmodqd3AOij1+Q7xCvBZU80j5RkkZ7UbfLruzWdSjLLEiwLvx7lc5flmCCrAQn7wiNOgMRJf8
1b+ttJTBTD42o1FCnXs8vjEPXDEQBM/GKxk/rtnEHzEJWZINEbYIqk4ujiAEsqm6CJ0ZMnIjlbSt
WPREv87+W7b6mm9FTX4fcCkBA6XsAVxzSb5ecAgavOnJ9/FaQky4w5k8Ip155INvO57zH5PuFyMc
gG0Ms6UO3+qnp51zGolXr1IMhqbUfsTC6PSkMOjJX4S/IjQqAM4UrEGt9Pxzph0HNYAe8JHdZMwk
YG8EYhvmQHMcdteODsJvLb8GkaaMrvp/YxF7AzKfRuzESc+2NcBW6v8gR0hYK4AJoz3o00salPI8
3BYrvy9GnCRQo5rWlwsWUGMBWa6/WK8p3z6krT+a11P5NSWXbL15GF4pn3/EDabCZM/TCEuCjrln
Xw6NXNmOuRu/gz9sQxxxBhjUHxE118aosFTPx0QtqlAyuqmUuHqpYWBK1mZdUhEQYKbBRpR2OIIR
dGHm4xzR8iXw8+nnpXKXWCAfv3ZqI+uZW/zOFPSY7P+tskD2iQEZRplDJzxoKzQX7zT8XIXKtjPz
sQUuveNnUEQsDvDT6hGQk7VL2X5XNfogMj0fr2BiqskmgHmiZtOf6T04kIrXHeSMYWWLcI591EKU
yi3aWMY3eKHifxN+YlAQ9itcjFgy2oULBsSkUsRFKc3Rh1Bpz3P/EVe/wfsG5BUd9fpBptvyptOm
7pKMsN7IDSB9Go8JBxSRxPCA/Oq+tU0Way0KZkaWAKLbUEtlFT9PMT5EYRtUwg9KbOvJ2rt7k8W6
KafmXWRn8I6vqTGEJNoIhJECgzwAFFuqQVJN3THfeYRv5gNJl4AEFSvW8zewg8jVMrOJUFnKQQXr
EBzJwVPiWfd2JUxqUgWh0Jq3Kt7dq9xIc/479ke/8qByWfPdP0B3ZH8dlcGIlQCOPQVx9eqmnzMQ
n++Aol4b8YTqM3qcR8UPdChaP1PC+lEJbxN+UcpggIIVP/zojfM+0m1NqxnqxMT+SAqAkVEJzfin
KKWOTpBs6yGAgKUa0B6QWDKfCJKpwoPWz/RhK3MRhf3t1VyYrmEfrCXq7EW0dTxPCrPwZ3jnGIWc
d40m8UNQkAIRVMl2+O9rnXEpfPGjKHqCXelk0+ysrVTpqy+sdvG/1Sc2MPyXnp1vIbglQSpZ3yPG
Jkobycsx0kEEZTPkMk86/q/OySCMkT4HhbvLCctshBm8J5tTNCNULdpzk8SxFweITZPaNiToZpMf
DBSrLfS9bUgb2bCfOtAmNarR94CNfkMfKfnz16cB5tR0a0ZS1F+Mg9dlb8gsidGNuKQrIl5hVu3i
HCnryIENiZF80fYGR92pkctdsG6zum3TJsspENRYm8JMSTiyvtY3ebcgV2P0ymyuNZdB9M9NGNAG
/5QBF/xDRDmCStcyZED+S9TIP9aYFv93pJ8dE1v0+02RqhfeGxVjebXg61U8WMGH/cvARSzk2cWA
pUXtEB33/SdE7+h8KLYsD/5SrX7ewRq/11wGfq38xCdkNIHDDmPWhwfnVxyY5gAcVS6qCO6cl4B7
bcwirOqqw3dujk4hsE6+bx71U00I9xdB7RQdADz5LwIrnUkPbu7sKjHo+lx1Q4TgEJXeOpIKQWNG
bv/J+WwtVIKM0DH02O/+46lc3uOxNTePIkl/AVrcuGXkntacEN4THapMnLMbAuqj4yg200FEt0SE
cqWIgqCaS6vw/jHj+eb+5FjLRRJLQ4c/GAa4mKSkUGWm31nCAsIksrTFuPfaKWBS/+AUjDibm7hj
4JNKMLT7fMS0sjKSxTk0a/SjV9+kjdvO6v+/Dep6h3FHDkRLTI0MF4jraQU05XbH53+AoYtSver0
7n8zYhl/yHzwXmvuT7USfxWok6X0vZLSilUx1Ghvf5WBbyinb4WB07wYn8AzLteFRCcEmRwQ4vVO
lEFKD2kBUHYEie+f6hngRt997t5sz6Ga4TBquwTL8JyX7J/kKlJSXrvsxUCTuQ4q/JXSU+wsOR/3
U5mpWtUSrxorIt3kQVI6LUn3u8QTAZBrALgRsBnJ9Lwj8TOX1uD6yF/xKB3nhH8FLzN50XwCKhqn
neYlQRnNufWhHlF7YNEpLBWvGsSybCnoIG9uGHUfTs2Df+vCITtAREr1ZXgsbMxSW2EXo4Qfd87o
mxOdcn1j9duwHJ61W94Uq0rVk84p7c/VKEU/iqhFo+cdhdptJ2SmUIj1ciyBREIkE6DzpCS69Wx5
78ROf3z2xIffpyvbSpcKnO73nL7EzDNjf6L5dtNFFaq8bv4pNdUaWhFkCknwPTSif08JlT9WPofF
uV/azW0ANjXOZmsxpKEXa3uT1p480ARZ1mTDaDHfZLAsET/Io9lg+B0mlEzfN1OKu9Blzq/PS/kX
ZWju8Ms3WJL5enwCcZCjdPGA4259qJg22EDmSlzPF1qi0gvSPuLs9un8SJ5FiBIoZibgapeX+fpi
PfsGFjM26TDnNM/ZivxyK8kT5AnXIn7KUGOwxihGI0lR515ZeqyviNz8MuylmuMVWrHES4rKZhzn
BV0AFwUS6H6PnK6QiuJ44feqOMw9sSbcTNzou7LezvgZxrX4WdnBPVFcOhMYHMzqdIsYgb2aJF6S
GLMbtDd2OLub5LfjYB8J9zynitV7PBLSyqE1EkFTIMM/Reozoh1sYguDpEwAEve2svJYEq2Wwifg
iA4MLchYu/IBkTO7gkzQtNZXlf68v2/Ey0KtGMVnyfeCpDj2bp4YqT2hzrDBJ2WWdjyMB0XKbzQP
yZzQEPd/e9t8iXcJuB3VygzSd4IpWiXCSXAwh367QkF7UZMQjwaaybjybtG0LtPM/YYt1bzDMedg
3Ulw9eVdrRtoZcIUfsEqDyJxzsbAVqfPrGLSH0SZTQIizue3I2eRXx8/rJ13xc87pAxTjnaPCufm
n0IeXCuNHnPUlQMgbcBpcG26VDyAAEx/pBjFc9UXFJ6rRdhpHbiicHK4VdjNhsBIWs1LZV3/hMtQ
x2ZeqCfKNVrGbUPV00gjZsKvEpbu7LUcjjTGx0J7ATzFFbURIYFB7fWuw4XeSIKvXDJdpLdp8FAi
dTlfawkng3nbnQ6Zm/t+HvehqfICNvgvsF20EXCwjRBy1b/ynt/pz6Bt+3JTffrWvEvts5Io+x2r
D34lvH/5DXUx6JTl8A5R+tNxii8u3W68ZkqMSbI3JpOw1j2XGleacTpFQsCqSyV2RkimR6U5EFkp
vpTeNQJzpv1/KPKeeof9uv9rsUHaoJ5h6E4DoJeuHlrlqEXNcSvGnBdL8Xv+WNq8uCy6CRo7n7em
D4M4piPvu719BkAoclpEmFVm7czbX9nbWOku9SCYDTglxcWKz3AFxQc3OKr9Lbepsk+0yVXOvdvg
0dtlJVYsU0mmACbBcDwgvecDSZW84aCoSR2UoDygF5+R1r6DYe/VE29B6nVrkRIu32ZcPAv5uTdR
OxF1RGtU4rtdllKbMdEfz+K2sO5+jbS3Wj+/1UXXBFTZ+v6kGM0ncojA09oKBXSRanIRxczaHwtM
KW9zl9KXgUIdlZC/XB/rytHM2sHEkYarhdjblx6UW8DUlMdcs6+eK2RUru9DWMRfLiXTESHWlX+J
J/qIGDqexz9mCrZ8Yt+Z7Gxgp7BKB0NWxlj0S/4n63ltX/wubmnBxpfovlRnxYovuB1/KrYi0WC6
jw570lFlQES7JygdWkyqXhiFXF6Y2DAytMiSFiZ/tn1svczdnLIjXbhIdCJV5okGszh6U1Oc877B
yur/CBepv5x32ZJbIGjJ6ZYiCyj1CQUW5h1yo3RD+ttkRn0DcVmW9o16WaZ9lF9edNLqKvIvJqKh
mqElv8CVs5Dr6lX/5y1HPFXIN53wlu6Oir24n4IPOSQQMORZyBwtmp+W7ERaG06tJYYw9BhxznLO
GtF6kTqYGxJonbHjKw3b+0d4ovEgBZK0aClwwzOTfPXBYIeSu4+lrn6nTcPVcX2gsEATfn/xaTCM
diFlTeFzXoGZHXygWa2SudL/HyijX5ARCwaj4N9qkt7NNJ421eGoOga/HtjT9LyQ8SkVxn6zK1Wj
9bOID436K5d6nP4em2UcoD3tV3s00rFUXILAVqQJ2V7tjYmA1qYx3LdxdFGFquKE7psG0B9J3D4S
LGVq8hBgSoADdPfKS1kzYSrIj4bUbg5W/8qSrO2eTjbtb4YDoxdlbXu1xflqtws4Kb+tEclGyuO0
H7HBGZJAAgPbHNv4A/Uc5H4klNKO/OKFX928MkcN6JHEUZAeaEQaIrZpSE1ZkzN6tZCQAXVdS/6y
8dzR1dBuUSApYCDZ7rLFTtLGTD6DKShc6psHHrjl6zeLfI/rh1/PeWBksibxz1L4x8MaY6Qjpalp
Qhhm1EpHjXiAYQkxaROyAVhNDRib9sT4S2QXjYD4WLhvTYGZ442B74bs0VoDG2mdrY/H1SDsfRMj
AY6YL8Ojf1aI2Mo6bUhNCOgYyZSrG8PHo177lTRzOfuQSssJ6ZHQ5uR1S/CBaJv0bPuo63b+ayxL
EOnkBbI5a89Jyl0ksFWbjKjqkzqytQkhXjAXEZchJ7Aqet8H+h+LUUJzRWiXWLH7AzHpxdFLLxPx
DFtmkJq7lunfjyZ5wq3m/j9gKkTjiVjUzZo40ig0JAF6zSl8E6zwwIF8idTCY2VefCT4RI+mEhgl
4rsh0QFduknxihGNx9aQFskxO4u8h1ZzK0SxRiybDQuy66uINk/QEhhmZ9i+/ecPfjQv+APxw5ms
2gXvyvVpcE5/eSLQo8WWcB14WPLeewOoJrz6H7cLeLQuuQM+KYcnIqtji4/R071IIm/HZQIIBbMf
hgGQH5ruVuDsqz1zUnm/fli29XBNvbsVIFFRQ+fGgpa06zE7/JF5rk8/AfQp7SkX45ffG0gPlIbM
LDSVGSDXpkiRVqIW3wd4DBDgM/lpIzwbOPPe5yY3bmsybWk8hNdFLWqhAvm1N0/nptmLUQz/N3LQ
5c+iaSUZwIJfZb0iwuvfbd3UuAQrcSTu0jGEclSafPM3yjtngukfxjqm2ZtaZa02M4Eo0+4ugi/n
o+qB44RHuDVwEI+zdffL/T137uvDHdNJgK4YNLCwLhD6gRS+epTJgEZcdtuES5nAHiHdanpvUImD
we+xemK9eHayiznV15DmLAdigsMJdMypMACfNOw/9P1vc2d4h9FS6YNgZks51sI/Hs7CFWoiQ0JD
cQQzEK9Ws/irFSKRzU87prN/vwMrH4g9qWy6VpMPLqzLU9fQE1cI1lPx6sRRyJkdkOJQDpcCFPKi
fgHKopZ2v/cgrB0SsWjUzpoBK3MzOIkZio2yOD5PCdTQSk5ROROB9N8QGuWp95kwDluZHUx02IB5
UdhkVjpFg9ImokZxFiB31BKTzzQOxwwZCRF8OT7xYC1lozcBDvcuNl4puX8O8YKTU+4iOXOtbgVq
wHLKIWjRdE0c9YYqzoY6+iItVZpzEo9kTVTo+znSBBrSeExnyKFziHphURBCwQ9eGgSE0ACjcs8Z
nsgq7Zb7bgAEscF/csPEsU0Spm1LIDBWlMEQKpWk5Y5aE6mZzuwJiuaATSOAvYi6EUgMO7ChoPxk
W8XlwiQPNK70k/yXKyRgCevX4jw4YbrUDIkSBHKQ5TQvUZnBaZDsC/zCOGOwik/0t4zDOxvgQ+lH
LKIHa36bAYbjcLa113y2wqEUQNw0iF+reHfKHYq+Ok5qdEGt29O5PFIuKLTNs5dKhM5EyCMOFYve
nE7xwNBqj0zCp3/H9jTiqShTpplaXsO10B/Ezw8E9agxftkyft0WUaB10rC4vj0i/84TH2Mbe+wk
Olds05Ohvpx5ZXHvAh3OxhUsdIdAJeP3drvKqwsioV+1LIKlk2OQsd+9mCxYf9KIl2ux4mZqzlMF
I0vPg/SiXhoGfGozJW//X2tMsWcp4f3VLGPC+cFsYE0MFwKDBe/YzY4u1o4wbyifMdk53sXzQZi+
QrWnKMwKtgqZWUnDud0JDm0Zfkm4/RMzkXp31qdIk4MgIPHzS29sH73jMiXCcrdB9z14atShvvpl
zjtb4mTLrFf30CE6rUPZFyctIbl5Zt7lVmIBWRGPg6mFZuyZsqtsVO5tsNV73+n+s8PBED1VF6wa
ROhQiCx5La/hGLqH7eUZoBrVjNh5tJqA+AvbeJkbHxEnY5pRD7Q5cv9BiQM4UVIYPbhyDxc3OcWx
QzxfN/7RJ4ZTUK7OjOk/JJ/JveSXSmCU7RaOBxEiRoqLaccfkxe+48J/w8gYjYdaQzRq3Je8Bc7C
Q9bniGBLgr726G3sxWEXRGZFVdy4baJ5qgVLpjjTUE860OHju4w3XPHBtgC16ajcDYFeqlbI4EQ7
xn3H223KPf+IcvWj4GkyMKx1LfbPWGFcc3XU4sQG8aaEoGkZ82NHVgYGEUZDaaFV0c7ZsgW26Bam
lTGFqx1/yu0LRnnVy5RrFlpEM2KCBCDPLik/TfRwobEkC0OeWdswfGUeA/2N8Z8s406mnlPlstDa
CqYnl4UiPQGYgtUWhkGRlX0WfTd1Hcc1HdcWr7Q6PyFnlI0MWR+6dwnNX5HP6kCnTkHD308CN3A0
nVKUuIyR3Xqi+XIU+fZjgoA/H3DjX9BDUrgcqEc9SQWgLoxpnOdWDTVYGT3qwS82T4oh1wzl19ZP
oHocq8yTZ3XLhtPp+olQAsyoGMd7+I6zINRNRgKldghOBfVyZ4Ga/CGv96fhGTnXtTrBkzsUis6n
uHx2zG1u1pqxiB4wVeHpC3f7Pti6qGISOKPCJEwDXXPeI0c7imzzdzLcji6x+mRrXtpR8+Kd0cA3
JuaifIvOGVPfD0iLkCNYg2Fzi5GNdnVdtyOSxAA24KReCuS2xFu7hQhuFj61ub49kyNIXAiutB5g
MjoFGQXXrNTROvzY89nlOxZ0MU1XZ6/rXe+Sg1QOAUWywkZxbEBPj8HFL60oHmSbww1kg9Llqk2f
dF1BrKAD/rHCfXCVULeKTTa7JUVCvqFTYhy8CPiniKEkfsMACfIrbzg0bE6K8pNSNnJj5JN5XjwF
pBVLoV5q4RrH+8euuelaiyXY5hXJvGnHYNqNKwgY0ys/+khkchA8FgcvWcym5SjWtjHrWmDwN3qJ
XUirV733N4SmE33FR/Zb4Zc3EYWrrvpqzBHFhHq95i8P/gZTTCqZRMAtP4CyxGY7iDq3rkE6lTFZ
nDboANJOtb+4Xg1bowdCMYP5xuPq0gOxoHTmIoLfPW6PsxZy/KTdpXqX5Je+MoMvuSMP92v3/nSL
zlgLIAc775K7oB5O7OuftGsoeBfoSZQMDylC8ejjH1fL6IfLXM5qdHPlsBv7SlyIS1Zd35CRpZwh
bvDBy+pr5RsKeznNLM7Qn9aU8koAmruJDl4hSGj6MGoUUftQ+UD1hOgdb0kLTr281eSEOAUNUBwt
iHHNXmtXF/0qLO+GJppJBzzObr8iJBkFN76HL0yN/hS3s2QBUcVVvtrubhQGtvcZ+1DH9W5vHX0M
RTnKBBRHT6AdhqWq+whtDZ6e+srbC7T4luZKGKCf5cqBCkB0Zo0J+EpD/X7qgU4q1k37hl6WVCt4
oCBS8451sdei3LidpRy+o8oohtnhFsnhznySLk/myBTfgqGX67JZxgerhvBoS5V/vUnmcLyRGprn
hMWfa+YdSIrQIyt0uyD6w47zbVU3thLGZtm9hskuZ2G6+JMiztlnefzSZFGtUsqFwt5CskyDAf53
HHwngGcCK0vIrMZlSGAtQqPB45GKyesTihC716fbjXO9ru8KQu8ODZ/7o/cYxSZJU6wa3WtO7NiH
u+ueVZiLzf1FW0YtmY+TzqbQrVOeLeGLvWHFBF2urnEl2QJ53ohRmSvfLsHKoRWar6mMv4ugYMuU
mfwBdCVuV3Qo0DDWm7R1RMwIdQzXY9qOsUu7ZIg+omdTBHW1FvLZSpy6S8PttPwtfD1ucu8p2VvP
K4AjHJ2Dwge1yP2OdVtn8r3c9ZnOzyr+Ek/CgBr8OP2ug1zEzmqtX11jIHzYicOywI7OjFf6SbVT
ID1FlP9drDmbSIaKf9UVW75s/D61a89pbO/TN9un/KiVaUrqWHpSf3X1St/2heXXkXpFQsisnbcY
mXP9xX57INTjRvtU/GM0hbZDf9p7Nz0+GdBdGf7cFCPXUTt0XulmLMFsbSSbnnN87af3uGhgrj6I
sp2wq3NEFZKM/T0UU+w1ERFtny1bOt7hCsSp3+fEZ/HJSA/5G96qdu63Ql+LBZm5ihwAwjJSfmmc
+fdBeqkFkCsyq30uS/L0RSEseMCQAzglbn6f3N3EnaxtRK3YXlBfN2yQRZ6EVs2SfLhRxZmqpGe5
3hWqz/hEcc4aOe9bjjZZaYLhmZdNifRQ8q8TrLE3YJOD3WTEln3/JcILyXOVKRGQ6Za2108oW36D
n54USLFtUTUpQzPXE+7oEMbr2J/wsM0qEVCTOsN7XUpzzTL2oRSJK9wIJUnL7PrNmpqtG9Xw6quT
vDWJqwDeTRQ+cvtoAU++QIO+otlUi/G01E3Mnf7agpbrWvD+eNgn9lrVnHLbdt81UpkPMa3ClcKi
URR4ZN6YNSnxcNF/5xYQTgjrrCd3Il9wcLe0HvbypVaTVb5hORU6XApWC3VoTr/BKNAPhAGysrzz
suNaZCXCjOuvAAIv+b/UrfvwxnpAo8GYuR2uS7urqps/TGisB6lm+Gz1qdNf7i0FD60cHE2/1SCc
J/xUIo/6Gq929kMnGFrYMALJafx/c5PDJMNgu5erP9b1EsYWwmeNkxwBd0fJrZBrm/Ej3q3DGhvA
pD6H5XQ+E7sEhc1vghyQmnk330qNDWxaRHG2wjP0mS1tO3/s5MtXzI+X1xgZzwi40k7h9prHOnI0
fXi4nHXEfdUybnzeC01Fpdrd0cIgLnjcp4KGuqOlcEAW7UNOMQ7x9pUTkyHPOlrGwxzOdYNUMDUG
AEWARe3T74IC5fVkrE87R2yhw49/jSlUVdmc0L6H3LZvcIqpmxAxUI8nfm941KFz/FOcdNvO+oJw
EFZhrXW7Ev8lcLZHzOekeW78fa2w8EXWAsc9YDpcRhM1YyhHc2JBvI8oGdyM8bv5o4gtFTDdhhYu
IN5BLbFnpE/SgW5NwNAaW9S0fW6wbhMd92UjPMcerleklcOL/j+2NyuoySe1GWMeYca3u1XIwN30
DBtBp/Boskip2GZbfHCAVrWyQ6NHFiGi8JtRLEJZrEW4npO55P3TC2bI2CLZV64RraujSOQ3MdZ1
hNA2jhRUZLEdyM4BA2RfTeCK4f43tEIqDYkUQ3jzfvLBwGT9sB2cksy3/L5I+8Rinv7tgDuDhUd6
fB4ZM3LIVFy8DPDNTK12SxPLFKWkM3mmoNtASpxtn4rFWJi8LM6C/jLfFOlLsY9IVBnloh0mpVSU
w59BZsQcwVtL3zbZdXfllUN5bdxwJfQGnc4DNx0ndyb0JPm+L4SzwTng+xnG4fkDcwUq1jgDqBnp
KL+Tf/CCZiOX+SsTjvri1K9GhDtV7xu9FpqVAXFUi/mVhx7edUTDB5Tus6SepbirvBEKJ1S2lpnC
G4T1xG5KcgMEufhNqaug3NrDeaNqKmyp9ZKU0G1DaxbtO96drzRWYDeNknpUWNbCpv/PMjlkkFIy
7ZXPT/YSM4avM+U8YT/u5KHywnJlO9MjFlAvW5ekE4CVDFy/v+dM6uNJk7bxTdE1XeFwxs+4W58B
9MRRc/PxQ6e/YQnd4zMN57RnF0HEsU3GMX+QNoNIKZ4eZ1mB1v3B3+xK1gAdUpFnaoUGK5Gr5CRc
jEQyNliY+qob9Q0iLVqOCs7/IZfa+2+DZv4itWYANRArxaoTYhGMTfZM39mUiSs6m/YueYBCuwGz
f/QHqHagX5NekYgRYSllw36a/urwHLceU0CL08M/wXd/M5EEskHLVYxzcrEA1JkoiXfZHZk0UsEg
yjr7XAJnIREwzaHJR+GQbhLzv51bbwaBH70YANQwwpbG1KavQcZzyXdACkFTiug3Jh8+Jf0t9/ne
JAXioeSV6IqeyBsGjbvzx5Yhof7QjSRfCGELQsn3Vl4DomsE/DHgR8HZtggdJrSPIDR6i+Ta16mg
IEM4xjE8NyJhzerYDlq4o6VxMS3KK604jPdJZssVBavYaWLI8ab4Qeyg5p3errvFmGcxyz1DYYt2
nURLdc0OyIxz3b71YDjIFQ/vT3d1Q819JaUpJ8Px4Le24Xid6/3yWaQ/2oiU8pTHiJT6oSM751Ur
aILouxynbqlNt8mebGPQ+p7wH+KBU2KsDHxhlnJ0xd1cU7JWhCV3kbRFEqHCTNvxO1pfFKMczGbN
wMrgE5AIiIWGDQH3keqn9vHL0nnGLmXnwxZ2UUdUtEg5/9gXRDBs4WZLqPLplMDuiBQ6gXnyrBjN
9KllhPTEChFZacyjIweqLQ57tKLMNvLGEFWY0ZKSTIPaTiRuvqzEXsRJhvQ1hNGJhXZNmmeewBkL
jUtJz+JlnJEwmyn40zAqm+H+CwXMVwJ27y88TQFOVtjcH7wk3dn9qWO8iyzfA4cvjAdt+7q4cvTD
oSngWmKCB58xBaFVK4mEQ9EsX4IwbVb3OakNQwnjDSZ8IWllZb0NzsQcmaux5/b0wE/fOSYP7CwZ
fgoPy6zbEN7rgcRe+aHWtLrPqiTELnjDWq11ltanNfCAM0TijSDouymktuDuULikzE3AucT4oc4C
6be/5gqFGk9Srnrctfl40Pko2TvLZnkhRuRBHQaDW30h9omu7wdxLV5uay+AzcnZFkgs7hy1Su8H
6ewL6HgGVl4ZLVpONVq52lwwo1UasbqdQo5CFBrcb7jC34Oc/Mq7R6bKojmk7wIv639lqjujXRkq
fYLwR9qV7C6kUFcZuLEyaCkhhsNO2jhLFKNpd4pHWFZOXqs6iUW6y9/ZNzfk01McqJ9fDwyAW0P6
ArFqIS0NbRcB2n5vsuew19bjyK/fv5urSLQ9jfmtWc2Ng2h3FRJxeT5qIgNbIdlGe6s+SZRnUYfz
hWbcE6XYaWXKvyOMijgQI6BdQISYp+TfT+tZjTv8U388HdP/v+gE0Yt2zmQ//z27IYGk4OoubuDS
TTyTb+VfteOhmO71FOZBTt+v2XXgOHiRoZdPtvSSARIUclWeYBbk8JQoNrdOvQ/prhhZoSh+M2VX
6udQ+/DXwnaorPIWC2NGlxRnJhb5Y8BOOFnAiYAFMw/g+8q7RpqIeTL7jqcM2cn7k//Wf0EeaqWM
02y6orrShunYrvvxNlVDTGFF5ODWYt8rMZMjMrudZWbjoVLSQWrw3XNMNj2BeoWskImjXNwGX1VW
CVfEce/qzs/asy0ehMnx4Oy7xMf8cLHVs8xRMTFed9bMj52t+mUpfZqRpN1lBvNNxl6W+nsKTl+v
YeKDF8QLu+qgKs68c/fR8DKJhs2GfC693lzesElthfuUtSHYo6mh+kIcPlcEsCR/zVv4AwwyEmgS
cQl590APp42my0SVothG0K1tKS5sSTJMApdIMMybh6tyZ0+No0bUdq0lP2SOD83lCrFpQaW/5W4S
p3AFixhGUpHMX5EwsHT5chLmMgyOo/JzIghH7Pw64ryh+8/p+KRzOADtEKlOVlMXTVPnD/Y5484t
QwKme+2mpkR/uGXb1/D8nypRiimmhMtJ9gb/tyDFm9TIpHkUM+aj9uqRisFX6J3F1CjXyn/bQQL+
+nqrPMwemLeWX388+dRZU0Jind2NRGXthuqgUbTqDK5Rd/R7wGLy7Os2IZSHuyD2ty4j9VQ2pO5Z
CTT5mDqhpUCi1WpnB6G9ejCgqeT5uD5mu/6yfkaWKY3iZWEgy2Veujba6JLgTpEwH65eV6w7Cz13
3Zmc98czcHglunbJha2v/J4nGDt+xn9ycl6CRPcax6RwYLp0VSmkVUA3MLDaIcRi1mW48CbrdD9l
ANilr8I3xwTU+5jsBP3H570LjKZC0v2FypIEa7pkZ9Upb9aZVQhD7lh1nkDgKHgaGjoG1LmJ/+Et
R7lgbPeIrFU8oX8CENvBR1rgR5NLc+Lav+fe3nI6Sf0t1K6v1M/OQy0J61i4fYP2lE/xfDzDTLva
YDWqkJCh2n71rFrfo4Yx29qU2tYkkHFVeNeV/6HOjVITL7eSvcrnscBrzEajtMdnVSf0xDHL72vG
maPyxnZLLA6cRJb6QNSMRpJ5X96FG3R32IrqXvnb8Yv9TikcerVzgh20nj4AWkJIGYXhoenVqHn3
pBmMMFq7NAIO0ZnnRA0Cqc5kUCZnG8qKF9uWSmBJPTBSnDiToJQxmcksi1VAlX49xzgKc/T+kHUo
EaksnbzLC3p5d71e4tlYsEB42G2/IfiHIdsCigIORGrSHczDP76fYZ+0AYHoFud9OzW7GEqJTpzL
R9KakaSGpLBQ0zqul3CslmdgbowxQNG56MC8sR8AEVRC0z1sUAAkkzlRCpAsloqc9n9Q+VQlCWHx
vDx6trQXoRFSqYCJ4070vNthF9GXxKWZnhIIKwrk5JOW5oq+AlfC4wA+X1NseDvc79MewmsxqNoY
rutrCxWtNH4um+RnBgMO4Gx+Ya4AkpyT3wf4xnrXC2fp6LwMmMMmnJHry2L0dWHg5IpWI+n0PIlf
kalqKIyMyYP1zduF5qEMZ+414QhJjQjhsNDZXkizhgtWPRm4QbQP2FO8tgm+Rq7haP8+GGnagLqO
UFDSUZEVoM5ckYhfddlXk4aDoURZrL5JE9mOSTaQx/5S3ZfFdDs+RUwEaS0qJH+sS+t54j1uhAXU
d6o6CNOT5ppBVPJBfVa5CEXQ5kyfClC6oQ3WP0Z3XQ/LXygyciYELo5p5qlLaKBcqF9s9OGcScVr
R1jg7BvG5zQ0RBkHbadaolM31DnSmY+Mb2ZpmNu8Q7paK9DX8uGTtV1okmkarsGso0qv3ZybB+8T
fPwy/YKuoZbpwhgykc7NInXhXifIqsSrrlTPMNTygCBesltbIF+xo32UYTwev2mVhVOkgTjvt4S3
qGuRd4ckCqKt7KfuSA1PeecNOF50wPzW2Mom+vHlyhUo54O9LHRkXUnBYnbc716qv1jYCJtPbnKX
Ufqv8oFIh9LWSoFWb5lkUn1W4MfRQq+ksMcCKHE1N4cD5KXfXIZyPEL/KHgXWczaD1xur5SGWVsE
pIx7cScCRON/mNW33iwoN+XDxNyb2VmGtzBbiteJH8CywAnNdrBjQnM9rZDi03GSGQoZcG/og1K8
YV8D8Sw+esNF7F0EoKu6222YRzdd3LWi39KREerjgVdCkQ6DcX8iR6qUG+AaIhh8aRqDqkL7FeH4
83oSAkZGROqSVl2MgIXH9Pn6si77zpS9uzDGT6i4Qf9ojET3QOMpiFPATX3sexQcUyAdlsFmR6ST
ot/BqJpYkaMMSdAlgm0Yamp+iu74T9HnMzQxDp5s/HL/H3QFEFz3Yk9ZeYSyb1dC0k0O4s4q8h1m
vlEeNrfkbPbHh+xAmZSwffzjNyDL4pqa0dB3HzAo2+fcWHqK7vRU2R6BQO7Ot5UNkRWfie/sT6ic
LAD2yB32kKegLG0lo7WkarnY9A2QxB8uKePTk/K6aJsmLk6bU28bVmWIdbAiwQZcYdjb4juc3M+F
chlyo1CkDXgneGEiaRO8zfkwQeza8aWfDVSRhzp2hrCRY4GqXmHuDeOICNqvAn3VMUE7N1v1mQOm
80oUQPgilHusqHQpI6gAc2sck13D1m0o1SAGycGOFYNzTI/AGMXdcMNNZpeUMUGDPAkQdSRvI58/
pRLrr64646rmA6JxCt7k9Tjlhx7yez99+o55JGyYQH78klk3fR/9cGeSfanH5pI/uKbjZ/BC7WkO
O3ObCROda4VmEJB9uINAHbpy3r0uJTFJIzvWW7fuAzKCzGoCHrVn8IlxIa2tUq0gkvd+j9kFFIS/
6bzNJG3qa5uiK+sgmRYq6X4g/MlKq3MCTj0NM2xa28/YX9uTRWZa0eGYB3raltGrq/BdLiTK2Kzu
P/a+31V7XZI41uOWXtX1UpQLHEhGxr8RxdI36feK0JFnX8eYHmtGNBYSo/uPNKg+NzbwqK/UTYBx
pxRA7xv9dggaLJbS9WrTIe4IpbhtrswdVi4syKxxLF/Se7X4BbREwzJNn3QfkWV9AHfEAMJF8qQI
Lf/N0rIh0cFKOebmFBAb0hmbded2wsv+Ef6q4QjUtWV7zY31wQPLZZ95hnj/bf+DOgC7I7DIrnIN
bZT3Q9LjfxpVLbxhOdhTYW7hcCFosrG7t0c2JP+RJX4h35/mf7q08x5B1JQhEkgtnegIqYySvjE4
BpH+sYGSCig2i1mYqWpuxfTfNf8I4dz15Bt/A7ixhxb/U9nLsX9TemV+SmUe+MjIJwpe1tW7wa4o
97NxbS2pgeZeFmYarZUPXOrIcS/xBY4WKZxmiRN+VjRW0vLZSzhtRlTdcmKeh8DGqJ5XbKSlKIGH
dw1sjnXh8FthDzVSVWpixE8rEbRiBLRNyGIuhfP/BogWkSWk1E9wqQePj+V24MG8xf4V4NJLpb2x
9TPpHqHC0A+NqHzOg5WqNyQ07wv6gzotpuKj94LAH7lc16rD/OJ4iTKjCL8Xa75MUizc5vF5XQcz
mGozFnJQVP1/vfgdaraZoGLVBcIeMWK9F3Bnn9MPHdcT61jFUnxo+NeniigG5SkKIJxyszR+heUa
9nwyBN9pJPfUEkSFzZeIIqaIHGHR+XFmXG7zQkjZWponeMxJsovML5Ts0E/JzhC4psfESo4wBWzo
ar+BUBE0xtS9o6/dUemxiHHpWCsMsqWp/xHMt72pagOVGYuWVRgdGStVAU3HoL0aV/j4WPbufkHz
wteZcQwPSJv6pwHe2G6vftxu6l7PzFASTxz7nAQ6DUmqYRiV5eUskWyANFRpnTSpP/toeYcUWFtl
tcbHPRRvE3sBEizaKAJp7xyf6f1YmoFJS8IpAc+o5XUcv0WUnJ3KgOKakqVNfCCQVAjyBJ29tO3g
PFSDjuWWFFxgvImkJvaozS2y4yiAyz4d2NO10vaBcbZqb2KGHFmHNgO2C5UTTSVTzyANIoaOQNwO
zZg2S+VPTw7zw3JYGOceEfnobrxLqNYalomxFAV2LbHzybrUOB557LPZ9qShkMAxXVdIKxY4muIu
M6moYN2NnOJq3iYPcW2AlPXFKsKPCnIpY+ARnLJuMrOYxzKaqyT6hRwAFaQe8N3Ig43jUoK/aCls
N6kEnwYLQ4hczq4MDU9I5+u+12zPUzG9OKKRshpgIbD0GVVYfUqhJ71LX+gWPxNKcgwKRRrUwEUF
vi3d/X+H5TH5aSBqPfd9R+chSJ4SCtaVOUQrGZw87RJYqTSnm5k9+9C9Aw/qOMhLyFMKHv1RrXvF
CYl5M8J8tMhCK2B+kj4gqwok4g+fLcvrMxoW8ztUe22g0dzkKGR1EDHeDvwG/CARoMaT6vCK8OZW
7CApcv27eKPbeyu5qx6bsR+fNzbCnRFmlYrTsWqre7x5G6bjiARCFfIZnGELz1B8qnXQfQZdpX9k
MVqZPvmI9EnpzZrVQ6aRSuMiSX1gsvnzONez5Tro2QRz8GAWqaO8U2kbJJPhSXSf20kppFZfcwtw
nhC1LIvOZxQ6XhckRhwvS/HDUawJrGIjn3dYwwOUcenutTgGtGpUAuNUyGj7tDhO/0BIS/fnEZrO
k02Pcnou+BccwEpp6kEKMDN4m0iifDQVxewU27k2rU9fGN9URRGSDCOtgjfjWFxKJCP+X6XIM/LQ
dhup1zJ9b2vg/JUGpPpkvulQbe8q3daojerwNsKki+Jn29ZZYWyrUTV7qG13CtnJrdJdswk5onQS
JDhXHTUcKH8oFMq5bO/OiSn5Wwkbv1BlOD+d3EMkGwc3V13uoa2MK8zEKRx1vth9vm9WM+W8f+cq
15jHQImWPzcHgTQPnlnDcPTKf6LRyUKcq1saD0Mt5ZZ73Fgd0qmJGPUtBTCS8QclSV6yFVJsuzy2
XJ5cgAIh02Aurj8VtGi3vvrX3HMoLzOjpuWMuvOc7a1smuCGMQYQEoCNrhy/MipTdM52BRLC6hf8
NSizsYz/YAXu0djF6k+HaieNK2weNVzKW6NH5zxTm3wwF6wSW0bq+QXAykJlYA5bNYV3V1Ai9phh
ppGtgWagj8WTx8GyA9bCEv096jKDrbpJLUSU5LGw0UIcbZzJvhmbxQ7uuu55KG4Cl8Fb01JeW1lC
YaWdqu5kwqfcFXe7mWRUvd4GvrvmivMUb2RqkAiyXSRUteLZxbgNyhuS0tFE1RrnZdGbSb1MXGmL
LjXsmDSYhbshKfuu1mOTo4LqC2sjvfo3wR6tXahvFH6yn7Nlm6XL/68wvmeUNM1XYPeCOD2OUrob
jLYNtM/78g7n7lf11edzEGWVIIrGOjvBc7DYguu/bClvmxMbnKB3MMygitZq4QjoAXv4IXzIyn05
fonn5TOlF0O0PokpvZA/dA9PbqOsdKW6Efd7BguNypmYqFlSJqCOhlfptPw9gQ60O/yPkjSNp69t
EeKErqTpYEc1lFQGBIK/olHaNjgSzSxunixwF+SnYHINgwP/a66Rh9ocUoXAVUzgJePc83VsL+lX
CE6+rAH5IAwZsb1EqIPhzY03o/FRAJOZFoaV/VjS3RAWKXH9VR2k54jCj0GfGPBk/xl8woleCXj9
DdmyPQsgypATwHXyqh2arZw5Zu4aUQsHbww6QzivndfuCNBoptz13MgarQsRve4zUnPTA0pPByzk
cDuWQHY+GhmuMMf3bwPWWlNWH7e2gY0LTui3+qphKv1/nse7QIs+UDpLRdOKHHaDGhxiOSL7lto2
+k3SHvo6GHzhqjQE6eUo+kGDojF5dn4ixf4qd3zqUDSE3i9kt9DLCfjLfmm4NFjINSz3xpEJK/nC
9z2s07Zk6TAUNnqe7Q4jAhczSRwpl1xqbJhuuFlbQ3169/3rbL4msubgCz0MoA3yE5s4MvU6SJQt
yyR3LgoDeWo9dgBaTMQ4HTTb+bC85tE0u5/VhWoQrNRJRtrjNrqgxDgSBOHkdLogs1nb6pqMpzIa
iRZnjTk08/BHHbqdGxR+aHEiss+V2qIPBd3IlOMoQr02+svvJ/jJB24n8zWv1Y18M7klwQDmFDYJ
Ya0+3GwUEXhbeXfpajEPeFEqQdjtcYb/CgjsRuEccErqkq+r3QDUq3tJkpTSRmZ7XoFX4KW0iNoj
HTD4VQvG3Sa+ngJCkLpt5WW9DdEg6QzHbJPPfkb4bUPoIZbyr7+Jkd0Hd1yKXGN2qvE1DfMOVHgB
xVKvJyLH5/Ja9G5wbEvjwD4zwvMwjmtQXKlYGugjBCTH+qekox2x7a/SD25Bz3QuGeQfG4MQa/Aw
+b38hAuLHFX4D0xAY8KPbqP925jH9HcCiYtHQYzyrNLUdvx+m+vREcJ9BArjfdLo6UjzSL7DPrD+
bkofvLEppgtwbE4IT5czk4TcU7C+T4qWdbmUpPoppQ8uO+w+B07smTWMsHG9Tl5asDqxgd2XKnJC
elXtkf4iw8n7NS4fu6P/JuhcLda4UYm3mAIGCJpYFQ+hQaoZ2+8O3o9D8iGSirHYG2Uf0hsZNXIF
gzieDZJxF4UBBXLgFPJdLpous0ZfOe5GL9l+0U7/ywaHkg5RhvgbF2B/dAOoNgqGn1CrDryjULvb
6Uxu9Qfjuwlxmf93xBa84fduUQ6VAia2qgSoV7Wwq5oqXC+qysVGTEMv/Z3BKtadIdMT3qxrJ5/Q
FIRp5YbZDRZTRLaQVCn5YTv4fJVb+Q9Sxopz9BAEKhmcTtWK0qfQtKIhFUGu5eFfxOGAxg5bAMVu
YHGVScVD1DxaKhXwqEW+NRUqYgYNKRKu8erj29tRlO8xiUHYfnbo4SJxMhOMYdHFGuQC6fDGd8lj
5NqPioSPd2IRHJemDnH/fmN7uAMTC+7/WCaqBw4Z9iN2ZqjavD2pI2BL6I9vhXHqGRVcHQ+QHd/Z
hrylRnYfMU5hdfmdb5VdVZqa9bw08lb+5+GO72BX8nvVvkIGxLbSl2uaFDSrsrCEHUxadcp0W03Y
PsQHHJOe2AC23U8VdYaL3FQo2SVVTEXJ38Ru1fShiRO48vv4gIUdjVQVgijZFKkI0x83N6NeaBLl
QfFa1UKxz3xnVjdUD5HTLDzAhL/ShRfxNFV0Uxy69zehl1QHflDDmyzhtvGPRMgyV7AjMql6d6Pu
JeltRXXOF31eMuN/hRAsbWtjlAeE3M8lNARiRIcQnbal5AGq+UZlXpyvFv23Y0pvSFoe4IngFNmi
K2rY7Ptfsd5ovA25VaTcmVFFPba0XhxA/h/MW9bjAK1r/gCOlt9Uarz0ucefld8c52tvCkFNAWog
H5OjZ/uxCzcZEpldWDUtZW9BAOKvBedKL7ICEnYUS9VnjaX9yqEZn8vdsdqmMesfdJexT1BGh/m1
xnz33QQ6c2XG4s3/JbK30jQghf/kwilrqJSgLXHykYCccPWgSSYujFNl3gCIgzBWToD8UavVUHuH
ZL+y+s8o8+t1FNObm/SJ0OvB8QNM6GoFnPd49T3xVYpffAXrBrPni2xkrxhnT5uH2SVqJb5Q+2hD
srJirXVnOUQH8USzwAVbBT68CZmqgu+jlwKTVSVAZfhw6tTaweAoXegmk73/QF3OJdomfI/+3P8j
bt93oqLFezQSyznOVG5dI/TZ05wwWSygIYeOiwJSSJjNphLvFF8t+tc4AcZrY3XmUdl/eWv4PC7I
eYAcLzOCORPF+W8RJwz38NeefBaGNO+5weSCE7q3mb8RriLgFg1R4NSwKZ48Oo/TT0zB0t7A0Kz/
bfo5Fq7+7lIw/tkGU2Vmm/n92wngsrF+nzKlCcMSoLoCaM9bhLHBG8XVjGaGG0udb8JB9aKFtYet
F0cZ06sDVS2bexlxeHRvusxzkNNwzQXayAWI5liznL2SFu4RpiA98Qqy9QqBIGyGFDhSRu+lqW6H
GvF+7JvjyKinG4+cK+kNnnBJEtUqg8LfZ0CbCnhgaWA392vkDGZbezkAdtFeqBseIjsVk7iUlesc
r1FzjwkfO6XtaL3NA5LDBWBJfvtVKhHP3qwRJ4iAH0K9iuYhgSxm3eX09wbCcuIl7qJZEAqtuOFe
Ef1MhnJNjBWUDCxEMWKzalXyiOI8tuIhiwyRz6z5HAiRxi6W4o/DGQAENhgvfCx/EaXDP+kJaXu5
+opn9m0mU7RTahaZlQLMYrTNlmaAbdE/D7Rh6DU7U8Ng2OWNDvVgjTWYW8dNyDx2ib6hNUHr29EU
GGpjVtmgx8ZJ96dCOKJ6W76PHBcbQJPA7GJ1lHnKX6xha/hsj+ierh7W9Nueir2LwEsIoRd3b0bM
nuXCv6vRiExGaDRTR8DTTMbs9QuZ5lJK/R+gp+6lw6SUuGX/lH8g+nbsPZTbAXj5USnfudWr8p8w
TJVE5Dw4V+h8I4eHwkLkh1aYPEBlTOqTX8szgQn8/Orff1txZUb5xsy7BYfiTkhmqV0kUzma/BrP
34Bebni0WaAT5SlL8DBH1eIo6s77Mm5hPZzIqTEEJXEaKSUTBmWXewtYv1kKhaW4yZxWLzf5LSky
4VhTpxA1HBiPbzrUmGQLsc8NAOKgDs1tR1jok6D0P8Ch2KK3RNCYWbGnvfJjokFMVZBPYhgv6Cqh
SAOGtaRdN7zoox9EVTc50P3gCSW5ND8jpiVJaJ1le0sqm2yu3ScaMmMl0gH+CZDLfX+QC2kMCnyq
M/QtHOXQ1zv6D00he56xkw9XBJ5ra1y7zDV1D0sTvneRXTVvlEKBS73B6cVv26bY/WlXCmHLlTta
xHInBX6ykMrRF956JP7W2p+jgiVIY8nCE/4yerGFL1vrF+adnKfCAazH/fLHADMAs8pWgbX3MvIv
FIt/mwFBeVliRuf1b5Zvpr0KqT687t+NVbJNYPLGy1ij5gXpYSYieM8vnZ+wtwOcNrMmroMZg6iL
ZiSKA1HaX/hj2RHDy02xcg0qi9WL2wbYVTQmF9QnkLZsUt6Or80zLKJ4dsXLgn3XezdlDOsRGP/v
9giNYXtv9pqbKUTmyK+P92KlelTBxpulXR/8j93aEj0NuhdD0u5VnEigC54TRhfxT8HSkjr9pM6J
Psyw+B0zVTFCx2sH6nT1x5uESOd34Dty4l8RuS8uzYsZcONZG/v8/tIzGAAHTQDUIwZw/x7mFE8I
9UBGqG6Tuau/dXFm6PYpOFCwuVmz7gEDj1nV7I/elE68xmi/rbTIYsVg5/YIPY6RPaA2j/BknDn7
DXMhjfkAQqq6wKsbj+i51LttX8lY4r1xZMQvc8Cn0X0ERgbAZqBNlHTsdBXMk2RRsH43xdi0D5hr
hPaFykOJJ0MHfhZYl+O7zGQMmkI2u2hD2J/Pn3EkxA3bq+K3bY2QPYtFUZ49IKi1FNHhBlhfXsVb
3XfdLFohADheBdzArcoQfB3cMH3k9Vd9UkAWvWjw8xArb4WvpoM09UewGCMECZ9nAS/o+GFd3z1v
vh9YbbnnFBuZNvyuUk2PL6zY652i4Ec4uqtcC5pTy5fKQyKHCGGCn1tdp/+s3L826B5Y8H81Ejbz
GMh0+q6aTMt8+YHI+B1g0/xuq8Ori6rwwcdVoCSDgjI5X/X7Nku/Rw8dpoHUOCEqdhm80f1JusLA
Szpv/sOgyqQ9wDSPP0cf7nFSriTxgD2/Az2XDIB3edHptb182Ljowb2/uNxGh4Uy0looUowg2KD/
dLtJAHsqGEONQgGEPWwuwFg0hewYpAMSJFFMgBFzw7irb5RUULNPbJ8CxkM6BalZk7qjkesSyhSD
vJ97pzFRd6G714SCsC4WOCHAMYfqQKPwt6OjoSw4hjintVdB3Fj3lMUzMbBUuszIB+RwgUrheV0I
QskgwMii/r2is7yZ3pWfT3sRY0S7bxrLVRhTNcvhBUJorhpPy4fp+tjPflvo2ko4pihNg7Wny7Ns
hRe351J4UzGW1QwEoeE4q9d21W//KDBvim4/LilXJXaynKLq6MA11dYNLLXB/xmRtzSlbEuBgR9v
QQa42HOgixmQF4FRiCwchdxP1mjolrlwT69elSifztzeiJTEN1FTyIL69DYrmLmq6X8RNVEWu60z
5K7DejBV4xWKm8yioT3w62I/e9W7XyR+CzyN5Wsc6rgnTYfUGZjz5LBED4qMF/6h1SD77lU3b5MG
S0JkT16HHMuVUtn1C54XE3WaEWoCxCgCiXSlbelm5JsWyi/oc/G0kdhCTy5egtlSnN6kIy5OE58Q
fHoPKIie6r62rzp6Gu3jDCJKuT3b/IgJwgTvzy5nF7k1qpLn6R5P/skxyv/E/bDtxsBPjnLeJHqh
4YZGyZpgfwI+VhQoJyGNn9JxkthyQMLHOYwO4jg+Y6CY4JTmBVISiuoPBaNOv4xc92PjxYa0w7QZ
CBjhgxfbWcQH3PjktzosPYia6AzkER5OAtP7Rl2d2wH7n+MvH6oIZjxIjh8LcGrWICWFbIvh3grc
jxoW/PqgSb+MmhoZTqsGnw9btZMjO3org8+R9JfoY9/jLROx8FoIxuk98ooj/TY4Ojh6EHMT7iAX
plWGydmECWUe/AelfojC+3EH67WJQu4AKKeyGDAMcIlPEy6GXUCLUrbA7LNtR27QXmBH5qtGRTii
A7O7ENSoUJpOxcBEnjll3RdSsl7Lovxol2I1xi4xgt/Z2Yw8EuD93utQ5WLBWNAns+QYICMbMqRt
HSmjdS8mjptqpBQr/zu4c1TmAVJmbvjYMiunihyLcpkx55nsfU+fxokgHsBkSVpJUS22ydCjiEY4
tdlasnnrSPyqh8b0JQ2naUcmDY73+XIrA4UN8JYqI5dfiWMNTw5bbZ3wvpWLRpreiKt+oPrVr54x
6pY2QGZ7k/LIDUbY73xNvIQHsEfHaGLUMV6G5DFaQVeaPyajpINrgEn//MHLPghb5g5b5bTOXbzG
Lg8HAdjzUNkUrHlZJfXnS+6FOd8vLFAzJkyIdYr/dCO6lcpHT7Z1BZCj0JXhFl9Cub44mX0waOab
JowNf8csMF52U5/gOVtLRKElyAfywrjbXZMNVLXQTljh2sVIP91fvaodxONlFPJimKywr9SJ42Tt
nLiuL9/g7XTefbXHK/cThdF7v7AS+Vq/SCgxba78CpJKKVLW5H5a4WI6NPrjtOI09MCqbbustHq2
/uatwNTjXoFVOcuIieBp9dz1DocIK7O+VBaIsycicZZAbqWCTKRBIg2w+DXVPDjC3RtPwx2aZtKG
/JEinpB4jXnvJCufgMXmg8sW3HpstxFlIIEA0GsqD7he8PZBX3qPltCghuBq5zgX3sLippebEys9
AQBMTZrFBok2YqIZEso159XEDZsLOV1CKU3YcqbBaxjPovDVdZHgHh9uni6ubrU0TKwm0oB0MJJJ
3RXbI/5+56PHULic6M0mSFc9GTOt5JCS3fg3rtRFOfrNBCZti/scDU9I3Az5+PPg9MtWuCRidZhp
TjpEZtvKJzIv/eOXgGSGbf3Pw9YnGPiBlgPJh7f9p5jtRU5ZOinLeJ7G4f6UO+j3WI7VQWZE0HAp
DlG27A5OCx9BBrFwDZOVlZv6NJPxR1XsOszk8DLuY95jYLWQFVWPF+pzIa0t3EzBDOT8puaTqyDl
TAPk0U+AXM/zWJryBAPH6Iu5DeTrBUEbNrbV8gdNdlxit9llt2tPzTRXaurJ7nLrY8CcDk8Sk948
DgVt35rVZ2fUYvFGUr+NL+4lZqSWfJT8bJFXYbtbj/5xBArNcCh3ga1QEk9hixi9Y5w+JotzC/65
oUyEs+WKcEUvJRsk/3ZyUMJcmKEwcSDqdKLBtL+UsUqMNwp7yws0hZwv1SduSZBl6vl/cHXNk3uX
NM2OKqb9mltbFxkN21ukcp5xi745HlvgRp5oiDXa+J4lQrDpbAaeIoEzhWyK4r91qRZhlUeqFEN0
/ip8SdnC4Okk0dB2BGa+lD1kIjuhvETUo7drXWt4fPGlmevtFSBl6Tkq0ZDt82SgOHv2rowy2Mth
4+0o7gkwSBTci/kSvIGXFnOVyIjPeRD0zNj29zuZOdPDnOpE1svCyiacSTraDTnK+meUztPqRbVM
ltBV0GDikg3317xUUUNCUtyhTywmRhm8O/cIRCURb1oDWKb6tIq7PUeE7n5yILgFHLetEgvqNwIN
76no0Jm6mfAkKf2JFluf/K2Y/SHRmY1gncxkfhRUvc4Bnthk8ZcDtY+r8co1lYROGHOASArD/w0E
b0Ue7Q6GuoiLKcRXj+YJDifn1ybT18gyhODqGhc3YT0w5RZ6GFV5M5FA9vKudYHKo0qNR+40aL3M
PWEhvz4+rO0niyVa2s7MhMmyjqfQP+8VBWexU3wsPJaCztByM87SlQlcx4Q2GygD+oMkOVWwKFBp
+j1eWbawhzQ/UBmk5xZ8nfaatg8dXeftgEOBJRaaBI2ZI2Y3lp91OpyHPrPpaBuKoI/mYryzLVuI
0UmrKQ/2EvmHMzPc0q3HMNvztyf/VLGs1GHqdbLuZUaxe5NF9JmyMJpd71k4/0hyVbE4usb1dTSb
gY5XtXVb0Nf5Fv3Ki+qlmGVlebSk/KbTt84/Ol/uYdhzQZAQ9sJLYRDlElScNcWvewRoI2rFUEou
M8OaPDR/sLUS8AeizEInSC0G2waf
`protect end_protected
