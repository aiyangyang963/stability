// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 16.1.2 Build 203 01/18/2017 SJ Standard Edition"

// DATE "10/27/2017 09:33:56"

// 
// Device: Altera 5CEBA4F17I7 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Qsys_system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	pio_key_export,
	pio_led0_export,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
input 	pio_key_export;
output 	pio_led0_export;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \onchip_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_rom|the_altsyncram|auto_generated|q_a[17] ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[4]~q ;
wire \jtag_uart_0|Add1~1_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[20]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[12]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[28]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \jtag_uart_0|Add1~5_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[16]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[8]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[24]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[2]~q ;
wire \jtag_uart_0|Add1~9_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[18]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[10]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[26]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[5]~q ;
wire \jtag_uart_0|Add1~13_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[21]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[13]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[29]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[7]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[23]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[15]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[31]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[11]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[27]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[9]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[25]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[6]~q ;
wire \jtag_uart_0|Add1~17_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[22]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[14]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[30]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[3]~q ;
wire \jtag_uart_0|Add1~21_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[19]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \jtag_uart_0|Add1~25_sumout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[17]~q ;
wire \mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ;
wire \pio_led|data_out~q ;
wire \jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|tdo~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ;
wire \nios2_qsys_0|d_address_offset_field[2]~q ;
wire \nios2_qsys_0|d_writedata[0]~q ;
wire \nios2_qsys_0|d_address_offset_field[0]~q ;
wire \jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|rst1~q ;
wire \nios2_qsys_0|d_write~q ;
wire \jtag_uart_0|always2~0_combout ;
wire \nios2_qsys_0|d_address_line_field[0]~q ;
wire \nios2_qsys_0|d_address_tag_field[1]~q ;
wire \nios2_qsys_0|d_address_tag_field[0]~q ;
wire \nios2_qsys_0|d_address_line_field[5]~q ;
wire \nios2_qsys_0|d_address_line_field[4]~q ;
wire \nios2_qsys_0|d_address_line_field[3]~q ;
wire \nios2_qsys_0|d_address_line_field[2]~q ;
wire \mm_interconnect_0|router|Equal3~0_combout ;
wire \nios2_qsys_0|d_address_line_field[1]~q ;
wire \nios2_qsys_0|d_address_tag_field[5]~q ;
wire \nios2_qsys_0|d_address_tag_field[4]~q ;
wire \nios2_qsys_0|d_address_tag_field[3]~q ;
wire \nios2_qsys_0|d_address_tag_field[2]~q ;
wire \mm_interconnect_0|router|Equal3~1_combout ;
wire \mm_interconnect_0|pio_led_s1_agent|m0_write~0_combout ;
wire \nios2_qsys_0|d_address_offset_field[1]~q ;
wire \mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \nios2_qsys_0|d_read~q ;
wire \mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_begintransfer~0_combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ;
wire \jtag_uart_0|av_waitrequest~0_combout ;
wire \mm_interconnect_0|router|Equal4~0_combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~1_combout ;
wire \mm_interconnect_0|pio_key_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart_0|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_rom_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_demux|WideOr0~combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ;
wire \nios2_qsys_0|i_read~q ;
wire \nios2_qsys_0|ic_fill_tag[4]~q ;
wire \nios2_qsys_0|ic_fill_tag[3]~q ;
wire \nios2_qsys_0|ic_fill_tag[2]~q ;
wire \nios2_qsys_0|ic_fill_tag[1]~q ;
wire \nios2_qsys_0|ic_fill_tag[0]~q ;
wire \nios2_qsys_0|ic_fill_line[6]~q ;
wire \mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux|src3_valid~1_combout ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_limiter|last_channel[0]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|WideOr1~combout ;
wire \mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|src2_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux|src6_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ;
wire \nios2_qsys_0|hbreak_enabled~q ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|save_dest_id~0_combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ;
wire \nios2_qsys_0|ic_fill_line[5]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \rst_controller|r_early_rst~q ;
wire \nios2_qsys_0|ic_fill_line[4]~q ;
wire \nios2_qsys_0|ic_fill_line[3]~q ;
wire \nios2_qsys_0|ic_fill_line[1]~q ;
wire \nios2_qsys_0|ic_fill_line[2]~q ;
wire \nios2_qsys_0|ic_fill_line[0]~q ;
wire \nios2_qsys_0|d_writedata[7]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \nios2_qsys_0|d_byteenable[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \jtag_uart_0|ien_AE~q ;
wire \jtag_uart_0|av_readdata[9]~combout ;
wire \jtag_uart_0|ien_AF~q ;
wire \jtag_uart_0|av_readdata[8]~0_combout ;
wire \pio_key|irq_mask~q ;
wire \pio_key|edge_capture~q ;
wire \nios2_qsys_0|d_writedata[3]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[16]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[18]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[19]~combout ;
wire \jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \nios2_qsys_0|d_writedata[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \jtag_uart_0|read_0~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[17]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~combout ;
wire \nios2_qsys_0|d_writedata[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[32]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[32]~combout ;
wire \nios2_qsys_0|d_writedata[20]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~1_combout ;
wire \nios2_qsys_0|d_byteenable[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[34]~combout ;
wire \nios2_qsys_0|d_writedata[12]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~2_combout ;
wire \nios2_qsys_0|d_byteenable[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[33]~combout ;
wire \nios2_qsys_0|d_writedata[28]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~3_combout ;
wire \nios2_qsys_0|d_byteenable[3]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~4_combout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[0]~q ;
wire \pio_key|readdata[0]~q ;
wire \pio_led|readdata[0]~combout ;
wire \nios2_qsys_0|d_writedata[16]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~5_combout ;
wire \nios2_qsys_0|d_writedata[8]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~6_combout ;
wire \nios2_qsys_0|d_writedata[24]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~7_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~combout ;
wire \nios2_qsys_0|d_writedata[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~8_combout ;
wire \nios2_qsys_0|d_writedata[18]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~9_combout ;
wire \nios2_qsys_0|d_writedata[10]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~10_combout ;
wire \jtag_uart_0|ac~q ;
wire \nios2_qsys_0|d_writedata[26]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~11_combout ;
wire \nios2_qsys_0|d_writedata[5]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~12_combout ;
wire \nios2_qsys_0|d_writedata[21]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~13_combout ;
wire \nios2_qsys_0|d_writedata[13]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~14_combout ;
wire \nios2_qsys_0|d_writedata[29]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~15_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~16_combout ;
wire \nios2_qsys_0|d_writedata[23]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~17_combout ;
wire \nios2_qsys_0|d_writedata[15]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~18_combout ;
wire \jtag_uart_0|rvalid~q ;
wire \nios2_qsys_0|d_writedata[31]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~19_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~combout ;
wire \nios2_qsys_0|d_writedata[11]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~20_combout ;
wire \nios2_qsys_0|d_writedata[27]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~21_combout ;
wire \nios2_qsys_0|d_writedata[9]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~22_combout ;
wire \nios2_qsys_0|d_writedata[25]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~23_combout ;
wire \nios2_qsys_0|d_writedata[6]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~24_combout ;
wire \nios2_qsys_0|d_writedata[22]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~25_combout ;
wire \nios2_qsys_0|d_writedata[14]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~26_combout ;
wire \jtag_uart_0|woverflow~q ;
wire \nios2_qsys_0|d_writedata[30]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~27_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~28_combout ;
wire \nios2_qsys_0|d_writedata[19]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~29_combout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~30_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~combout ;
wire \nios2_qsys_0|d_writedata[17]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \pio_key_export~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


Qsys_system_Qsys_system_jtag_uart_0 jtag_uart_0(
	.q_b_4(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.Add1(\jtag_uart_0|Add1~1_sumout ),
	.q_b_0(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.Add11(\jtag_uart_0|Add1~5_sumout ),
	.q_b_2(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.Add12(\jtag_uart_0|Add1~9_sumout ),
	.q_b_5(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.Add13(\jtag_uart_0|Add1~13_sumout ),
	.q_b_7(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.Add14(\jtag_uart_0|Add1~17_sumout ),
	.q_b_3(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.Add15(\jtag_uart_0|Add1~21_sumout ),
	.q_b_1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.Add16(\jtag_uart_0|Add1~25_sumout ),
	.tdo(\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|tdo~q ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.rst1(\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_write(\nios2_qsys_0|d_write~q ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.d_address_line_field_0(\nios2_qsys_0|d_address_line_field[0]~q ),
	.Equal3(\mm_interconnect_0|router|Equal3~0_combout ),
	.Equal31(\mm_interconnect_0|router|Equal3~1_combout ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.suppress_change_dest_id(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~0_combout ),
	.av_waitrequest2(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.cp_valid(\mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~0_combout ),
	.last_channel_0(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|last_channel[0]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.b_full(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~q ),
	.b_non_empty(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.ien_AE1(\jtag_uart_0|ien_AE~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.ien_AF1(\jtag_uart_0|ien_AF~q ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~q ),
	.b_full1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~q ),
	.read_01(\jtag_uart_0|read_0~q ),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~q ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~q ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~q ),
	.ac1(\jtag_uart_0|ac~q ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~q ),
	.rvalid1(\jtag_uart_0|rvalid~q ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~q ),
	.woverflow1(\jtag_uart_0|woverflow~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

Qsys_system_Qsys_system_nios2_qsys_0 nios2_qsys_0(
	.readdata_4(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[4]~q ),
	.readdata_20(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[20]~q ),
	.readdata_12(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[12]~q ),
	.readdata_28(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[28]~q ),
	.readdata_16(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[16]~q ),
	.readdata_8(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[8]~q ),
	.readdata_24(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[24]~q ),
	.readdata_2(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[2]~q ),
	.readdata_18(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[18]~q ),
	.readdata_10(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[10]~q ),
	.readdata_26(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[26]~q ),
	.readdata_5(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[5]~q ),
	.readdata_21(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[21]~q ),
	.readdata_13(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[13]~q ),
	.readdata_29(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[29]~q ),
	.readdata_7(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[7]~q ),
	.readdata_23(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[23]~q ),
	.readdata_15(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[15]~q ),
	.readdata_31(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[31]~q ),
	.readdata_11(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[11]~q ),
	.readdata_27(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[27]~q ),
	.readdata_9(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[9]~q ),
	.readdata_25(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[25]~q ),
	.readdata_6(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[6]~q ),
	.readdata_22(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[22]~q ),
	.readdata_14(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[14]~q ),
	.readdata_30(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[30]~q ),
	.readdata_3(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[3]~q ),
	.readdata_19(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[19]~q ),
	.readdata_17(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[17]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.sr_0(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ),
	.ir_out_0(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ),
	.ir_out_1(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.rst1(\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_write1(\nios2_qsys_0|d_write~q ),
	.d_address_line_field_0(\nios2_qsys_0|d_address_line_field[0]~q ),
	.d_address_tag_field_1(\nios2_qsys_0|d_address_tag_field[1]~q ),
	.d_address_tag_field_0(\nios2_qsys_0|d_address_tag_field[0]~q ),
	.d_address_line_field_5(\nios2_qsys_0|d_address_line_field[5]~q ),
	.d_address_line_field_4(\nios2_qsys_0|d_address_line_field[4]~q ),
	.d_address_line_field_3(\nios2_qsys_0|d_address_line_field[3]~q ),
	.d_address_line_field_2(\nios2_qsys_0|d_address_line_field[2]~q ),
	.d_address_line_field_1(\nios2_qsys_0|d_address_line_field[1]~q ),
	.d_address_tag_field_5(\nios2_qsys_0|d_address_tag_field[5]~q ),
	.d_address_tag_field_4(\nios2_qsys_0|d_address_tag_field[4]~q ),
	.d_address_tag_field_3(\nios2_qsys_0|d_address_tag_field[3]~q ),
	.d_address_tag_field_2(\nios2_qsys_0|d_address_tag_field[2]~q ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_read1(\nios2_qsys_0|d_read~q ),
	.av_begintransfer(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_begintransfer~0_combout ),
	.suppress_change_dest_id(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.jtag_debug_module_waitrequest(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr01(\mm_interconnect_0|cmd_demux|WideOr0~combout ),
	.av_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ),
	.d_readdatavalid(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.has_pending_responses(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ),
	.i_read1(\nios2_qsys_0|i_read~q ),
	.ic_fill_tag_4(\nios2_qsys_0|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\nios2_qsys_0|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\nios2_qsys_0|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\nios2_qsys_0|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\nios2_qsys_0|ic_fill_tag[0]~q ),
	.ic_fill_line_6(\nios2_qsys_0|ic_fill_line[6]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.rf_source_valid(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.hbreak_enabled1(\nios2_qsys_0|hbreak_enabled~q ),
	.save_dest_id(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|save_dest_id~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.suppress_change_dest_id1(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.ic_fill_line_5(\nios2_qsys_0|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.ic_fill_line_4(\nios2_qsys_0|ic_fill_line[4]~q ),
	.ic_fill_line_3(\nios2_qsys_0|ic_fill_line[3]~q ),
	.ic_fill_line_1(\nios2_qsys_0|ic_fill_line[1]~q ),
	.ic_fill_line_2(\nios2_qsys_0|ic_fill_line[2]~q ),
	.ic_fill_line_0(\nios2_qsys_0|ic_fill_line[0]~q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\nios2_qsys_0|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\nios2_qsys_0|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\nios2_qsys_0|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.d_byteenable_0(\nios2_qsys_0|d_byteenable[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.irq_mask(\pio_key|irq_mask~q ),
	.edge_capture(\pio_key|edge_capture~q ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~q ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.d_readdata({\mm_interconnect_0|rsp_mux|src_data[31]~combout ,\mm_interconnect_0|rsp_mux|src_data[30]~combout ,\mm_interconnect_0|rsp_mux|src_data[29]~combout ,\mm_interconnect_0|rsp_mux|src_data[28]~combout ,\mm_interconnect_0|rsp_mux|src_data[27]~combout ,
\mm_interconnect_0|rsp_mux|src_data[26]~combout ,\mm_interconnect_0|rsp_mux|src_data[25]~combout ,\mm_interconnect_0|rsp_mux|src_data[24]~combout ,\mm_interconnect_0|rsp_mux|src_data[23]~combout ,\mm_interconnect_0|rsp_mux|src_data[22]~combout ,
\mm_interconnect_0|rsp_mux|src_data[21]~combout ,\mm_interconnect_0|rsp_mux|src_data[20]~combout ,\mm_interconnect_0|rsp_mux|src_data[19]~combout ,\mm_interconnect_0|rsp_mux|src_data[18]~combout ,\mm_interconnect_0|rsp_mux|src_data[17]~combout ,
\mm_interconnect_0|rsp_mux|src_data[16]~combout ,\mm_interconnect_0|rsp_mux|src_data[15]~combout ,\mm_interconnect_0|rsp_mux|src_data[14]~combout ,\mm_interconnect_0|rsp_mux|src_data[13]~combout ,\mm_interconnect_0|rsp_mux|src_data[12]~combout ,
\mm_interconnect_0|rsp_mux|src_data[11]~combout ,\mm_interconnect_0|rsp_mux|src_data[10]~combout ,\mm_interconnect_0|rsp_mux|src_data[9]~combout ,\mm_interconnect_0|rsp_mux|src_data[8]~combout ,\mm_interconnect_0|rsp_mux|src_data[7]~combout ,
\mm_interconnect_0|rsp_mux|src_data[6]~combout ,\mm_interconnect_0|rsp_mux|src_data[5]~combout ,\mm_interconnect_0|rsp_mux|src_data[4]~combout ,\mm_interconnect_0|rsp_mux|src_data[3]~combout ,\mm_interconnect_0|rsp_mux|src_data[2]~combout ,
\mm_interconnect_0|rsp_mux|src_data[1]~combout ,\mm_interconnect_0|rsp_mux|src_data[0]~combout }),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~q ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.i_readdata({\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[0]~combout }),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~q ),
	.d_writedata_20(\nios2_qsys_0|d_writedata[20]~q ),
	.d_byteenable_2(\nios2_qsys_0|d_byteenable[2]~q ),
	.d_writedata_12(\nios2_qsys_0|d_writedata[12]~q ),
	.d_byteenable_1(\nios2_qsys_0|d_byteenable[1]~q ),
	.d_writedata_28(\nios2_qsys_0|d_writedata[28]~q ),
	.d_byteenable_3(\nios2_qsys_0|d_byteenable[3]~q ),
	.readdata_0(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[0]~q ),
	.d_writedata_16(\nios2_qsys_0|d_writedata[16]~q ),
	.d_writedata_8(\nios2_qsys_0|d_writedata[8]~q ),
	.d_writedata_24(\nios2_qsys_0|d_writedata[24]~q ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~q ),
	.d_writedata_18(\nios2_qsys_0|d_writedata[18]~q ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~q ),
	.d_writedata_26(\nios2_qsys_0|d_writedata[26]~q ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~q ),
	.d_writedata_21(\nios2_qsys_0|d_writedata[21]~q ),
	.d_writedata_13(\nios2_qsys_0|d_writedata[13]~q ),
	.d_writedata_29(\nios2_qsys_0|d_writedata[29]~q ),
	.d_writedata_23(\nios2_qsys_0|d_writedata[23]~q ),
	.d_writedata_15(\nios2_qsys_0|d_writedata[15]~q ),
	.d_writedata_31(\nios2_qsys_0|d_writedata[31]~q ),
	.d_writedata_11(\nios2_qsys_0|d_writedata[11]~q ),
	.d_writedata_27(\nios2_qsys_0|d_writedata[27]~q ),
	.d_writedata_9(\nios2_qsys_0|d_writedata[9]~q ),
	.d_writedata_25(\nios2_qsys_0|d_writedata[25]~q ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~q ),
	.d_writedata_22(\nios2_qsys_0|d_writedata[22]~q ),
	.d_writedata_14(\nios2_qsys_0|d_writedata[14]~q ),
	.d_writedata_30(\nios2_qsys_0|d_writedata[30]~q ),
	.d_writedata_19(\nios2_qsys_0|d_writedata[19]~q ),
	.jtag_debug_module_resetrequest(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.readdata_1(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[1]~q ),
	.d_writedata_17(\nios2_qsys_0|d_writedata[17]~q ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

Qsys_system_Qsys_system_mm_interconnect_0 mm_interconnect_0(
	.q_a_4(\onchip_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_41(\onchip_rom|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_201(\onchip_rom|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_12(\onchip_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_121(\onchip_rom|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\onchip_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_281(\onchip_rom|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_0(\onchip_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_01(\onchip_rom|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_161(\onchip_rom|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\onchip_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_81(\onchip_rom|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\onchip_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_241(\onchip_rom|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_2(\onchip_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_21(\onchip_rom|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_18(\onchip_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_181(\onchip_rom|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_10(\onchip_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_101(\onchip_rom|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\onchip_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_261(\onchip_rom|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_5(\onchip_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_51(\onchip_rom|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_211(\onchip_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_212(\onchip_rom|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\onchip_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_131(\onchip_rom|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\onchip_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_291(\onchip_rom|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_7(\onchip_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_71(\onchip_rom|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_231(\onchip_rom|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_151(\onchip_rom|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_311(\onchip_rom|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\onchip_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_111(\onchip_rom|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\onchip_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_271(\onchip_rom|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_9(\onchip_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_91(\onchip_rom|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_25(\onchip_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_251(\onchip_rom|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_6(\onchip_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_61(\onchip_rom|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\onchip_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_221(\onchip_rom|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\onchip_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_141(\onchip_rom|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\onchip_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_301(\onchip_rom|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_3(\onchip_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_32(\onchip_rom|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_191(\onchip_rom|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_1(\onchip_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_rom|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_171(\onchip_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_172(\onchip_rom|the_altsyncram|auto_generated|q_a[17] ),
	.q_b_4(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.readdata_4(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[4]~q ),
	.Add1(\jtag_uart_0|Add1~1_sumout ),
	.readdata_20(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[20]~q ),
	.readdata_12(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[12]~q ),
	.readdata_28(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[28]~q ),
	.q_b_0(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.Add11(\jtag_uart_0|Add1~5_sumout ),
	.readdata_16(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[16]~q ),
	.readdata_8(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[8]~q ),
	.readdata_24(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[24]~q ),
	.q_b_2(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.readdata_2(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[2]~q ),
	.Add12(\jtag_uart_0|Add1~9_sumout ),
	.readdata_18(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[18]~q ),
	.readdata_10(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[10]~q ),
	.readdata_26(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[26]~q ),
	.q_b_5(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.readdata_5(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[5]~q ),
	.Add13(\jtag_uart_0|Add1~13_sumout ),
	.readdata_21(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[21]~q ),
	.readdata_13(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[13]~q ),
	.readdata_29(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[29]~q ),
	.q_b_7(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.readdata_7(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[7]~q ),
	.readdata_23(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[23]~q ),
	.readdata_15(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[15]~q ),
	.readdata_31(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[31]~q ),
	.readdata_11(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[11]~q ),
	.readdata_27(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[27]~q ),
	.readdata_9(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[9]~q ),
	.readdata_25(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[25]~q ),
	.q_b_6(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.readdata_6(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[6]~q ),
	.Add14(\jtag_uart_0|Add1~17_sumout ),
	.readdata_22(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[22]~q ),
	.readdata_14(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[14]~q ),
	.readdata_30(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[30]~q ),
	.q_b_3(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.readdata_3(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[3]~q ),
	.Add15(\jtag_uart_0|Add1~21_sumout ),
	.readdata_19(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[19]~q ),
	.q_b_1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.Add16(\jtag_uart_0|Add1~25_sumout ),
	.readdata_17(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[17]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.rst1(\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_write(\nios2_qsys_0|d_write~q ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.d_address_line_field_0(\nios2_qsys_0|d_address_line_field[0]~q ),
	.d_address_tag_field_1(\nios2_qsys_0|d_address_tag_field[1]~q ),
	.d_address_tag_field_0(\nios2_qsys_0|d_address_tag_field[0]~q ),
	.d_address_line_field_5(\nios2_qsys_0|d_address_line_field[5]~q ),
	.d_address_line_field_4(\nios2_qsys_0|d_address_line_field[4]~q ),
	.d_address_line_field_3(\nios2_qsys_0|d_address_line_field[3]~q ),
	.d_address_line_field_2(\nios2_qsys_0|d_address_line_field[2]~q ),
	.Equal3(\mm_interconnect_0|router|Equal3~0_combout ),
	.d_address_line_field_1(\nios2_qsys_0|d_address_line_field[1]~q ),
	.d_address_tag_field_5(\nios2_qsys_0|d_address_tag_field[5]~q ),
	.d_address_tag_field_4(\nios2_qsys_0|d_address_tag_field[4]~q ),
	.d_address_tag_field_3(\nios2_qsys_0|d_address_tag_field[3]~q ),
	.d_address_tag_field_2(\nios2_qsys_0|d_address_tag_field[2]~q ),
	.Equal31(\mm_interconnect_0|router|Equal3~1_combout ),
	.m0_write(\mm_interconnect_0|pio_led_s1_agent|m0_write~0_combout ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_read(\nios2_qsys_0|d_read~q ),
	.av_begintransfer(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_begintransfer~0_combout ),
	.suppress_change_dest_id(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ),
	.av_waitrequest(\jtag_uart_0|av_waitrequest~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~0_combout ),
	.suppress_change_dest_id1(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~1_combout ),
	.mem_used_1(\mm_interconnect_0|pio_key_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[0]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.mem_used_11(\mm_interconnect_0|onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_12(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ),
	.mem_used_13(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_02(\mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ),
	.mem_used_14(\mm_interconnect_0|onchip_rom_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr01(\mm_interconnect_0|cmd_demux|WideOr0~combout ),
	.av_waitrequest2(\mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ),
	.cp_valid(\mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.has_pending_responses(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ),
	.i_read(\nios2_qsys_0|i_read~q ),
	.ic_fill_tag_4(\nios2_qsys_0|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\nios2_qsys_0|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\nios2_qsys_0|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\nios2_qsys_0|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\nios2_qsys_0|ic_fill_tag[0]~q ),
	.ic_fill_line_6(\nios2_qsys_0|ic_fill_line[6]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.src3_valid(\mm_interconnect_0|cmd_demux|src3_valid~1_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.last_channel_0(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|last_channel[0]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.WideOr11(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.rf_source_valid(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.src2_valid(\mm_interconnect_0|cmd_demux_001|src2_valid~0_combout ),
	.src6_valid(\mm_interconnect_0|cmd_demux|src6_valid~0_combout ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.hbreak_enabled(\nios2_qsys_0|hbreak_enabled~q ),
	.save_dest_id(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|save_dest_id~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.suppress_change_dest_id2(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.ic_fill_line_5(\nios2_qsys_0|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.b_full(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.ic_fill_line_4(\nios2_qsys_0|ic_fill_line[4]~q ),
	.ic_fill_line_3(\nios2_qsys_0|ic_fill_line[3]~q ),
	.ic_fill_line_1(\nios2_qsys_0|ic_fill_line[1]~q ),
	.ic_fill_line_2(\nios2_qsys_0|ic_fill_line[2]~q ),
	.ic_fill_line_0(\nios2_qsys_0|ic_fill_line[0]~q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~q ),
	.b_non_empty(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\nios2_qsys_0|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\nios2_qsys_0|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\nios2_qsys_0|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.d_byteenable_0(\nios2_qsys_0|d_byteenable[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.ien_AE(\jtag_uart_0|ien_AE~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.ien_AF(\jtag_uart_0|ien_AF~q ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~q ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux|src_data[28]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux|src_data[24]~combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux|src_data[26]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[21]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux|src_data[29]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[31]~combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux|src_data[27]~combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux|src_data[25]~combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux|src_data[30]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~combout ),
	.b_full1(\jtag_uart_0|the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~q ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.read_0(\jtag_uart_0|read_0~q ),
	.src_data_51(\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ),
	.src_data_33(\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ),
	.src_data_47(\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ),
	.src_data_210(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.src_data_281(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_301(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_311(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_data_271(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_291(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.src_data_231(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_251(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_261(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.src_data_221(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.src_data_241(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_171(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.src_data_161(\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ),
	.src_data_151(\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ),
	.src_data_131(\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ),
	.src_data_141(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.src_data_121(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_471(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_382(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_392(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_402(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_412(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_422(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_432(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_442(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_452(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_462(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_472(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.src_data_481(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_491(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_322(\mm_interconnect_0|cmd_mux_006|src_data[32]~combout ),
	.d_writedata_20(\nios2_qsys_0|d_writedata[20]~q ),
	.src_payload6(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.d_byteenable_2(\nios2_qsys_0|d_byteenable[2]~q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_006|src_data[34]~combout ),
	.d_writedata_12(\nios2_qsys_0|d_writedata[12]~q ),
	.src_payload8(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.d_byteenable_1(\nios2_qsys_0|d_byteenable[1]~q ),
	.src_data_331(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_data_332(\mm_interconnect_0|cmd_mux_006|src_data[33]~combout ),
	.d_writedata_28(\nios2_qsys_0|d_writedata[28]~q ),
	.src_payload10(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.d_byteenable_3(\nios2_qsys_0|d_byteenable[3]~q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_006|src_data[35]~combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.readdata_0(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[0]~q ),
	.readdata_01(\pio_key|readdata[0]~q ),
	.readdata_02(\pio_led|readdata[0]~combout ),
	.d_writedata_16(\nios2_qsys_0|d_writedata[16]~q ),
	.src_payload14(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.d_writedata_8(\nios2_qsys_0|d_writedata[8]~q ),
	.src_payload16(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.d_writedata_24(\nios2_qsys_0|d_writedata[24]~q ),
	.src_payload18(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_data_81(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~q ),
	.src_payload20(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.d_writedata_18(\nios2_qsys_0|d_writedata[18]~q ),
	.src_payload22(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~q ),
	.src_payload24(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.ac(\jtag_uart_0|ac~q ),
	.d_writedata_26(\nios2_qsys_0|d_writedata[26]~q ),
	.src_payload26(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~q ),
	.src_payload28(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.d_writedata_21(\nios2_qsys_0|d_writedata[21]~q ),
	.src_payload30(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.d_writedata_13(\nios2_qsys_0|d_writedata[13]~q ),
	.src_payload32(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.d_writedata_29(\nios2_qsys_0|d_writedata[29]~q ),
	.src_payload34(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_data_181(\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.d_writedata_23(\nios2_qsys_0|d_writedata[23]~q ),
	.src_payload38(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.d_writedata_15(\nios2_qsys_0|d_writedata[15]~q ),
	.src_payload40(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.rvalid(\jtag_uart_0|rvalid~q ),
	.d_writedata_31(\nios2_qsys_0|d_writedata[31]~q ),
	.src_payload42(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_data_172(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.d_writedata_11(\nios2_qsys_0|d_writedata[11]~q ),
	.src_payload44(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.d_writedata_27(\nios2_qsys_0|d_writedata[27]~q ),
	.src_payload46(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.d_writedata_9(\nios2_qsys_0|d_writedata[9]~q ),
	.src_payload48(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.d_writedata_25(\nios2_qsys_0|d_writedata[25]~q ),
	.src_payload50(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.d_writedata_22(\nios2_qsys_0|d_writedata[22]~q ),
	.src_payload54(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.d_writedata_14(\nios2_qsys_0|d_writedata[14]~q ),
	.src_payload56(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.woverflow(\jtag_uart_0|woverflow~q ),
	.d_writedata_30(\nios2_qsys_0|d_writedata[30]~q ),
	.src_payload58(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ),
	.src_data_61(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_201(\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ),
	.src_data_191(\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.d_writedata_19(\nios2_qsys_0|d_writedata[19]~q ),
	.src_payload62(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.readdata_1(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|readdata[1]~q ),
	.src_payload65(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.d_writedata_17(\nios2_qsys_0|d_writedata[17]~q ),
	.src_payload67(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_342(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_data_352(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload75(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload76(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload79(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_data_333(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload82(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload83(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload87(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload88(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload89(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload90(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload91(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload92(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload93(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload94(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload95(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload96(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

Qsys_system_Qsys_system_pio_led pio_led(
	.data_out1(\pio_led|data_out~q ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.m0_write(\mm_interconnect_0|pio_led_s1_agent|m0_write~0_combout ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_led_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.readdata_0(\pio_led|readdata[0]~combout ),
	.clk(\clk_clk~input_o ));

Qsys_system_Qsys_system_pio_key pio_key(
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.rst1(\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_write(\nios2_qsys_0|d_write~q ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.Equal4(\mm_interconnect_0|router|Equal4~0_combout ),
	.mem_used_1(\mm_interconnect_0|pio_key_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_key_s1_translator|wait_latency_counter[0]~q ),
	.irq_mask1(\pio_key|irq_mask~q ),
	.edge_capture1(\pio_key|edge_capture~q ),
	.readdata_0(\pio_key|readdata[0]~q ),
	.clk(\clk_clk~input_o ),
	.in_port(\pio_key_export~input_o ));

Qsys_system_Qsys_system_onchip_rom onchip_rom(
	.q_a_4(\onchip_rom|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_rom|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_12(\onchip_rom|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\onchip_rom|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_0(\onchip_rom|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_rom|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\onchip_rom|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\onchip_rom|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_2(\onchip_rom|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_18(\onchip_rom|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_10(\onchip_rom|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\onchip_rom|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_5(\onchip_rom|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_rom|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\onchip_rom|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\onchip_rom|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_7(\onchip_rom|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_rom|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_rom|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_rom|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\onchip_rom|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\onchip_rom|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_9(\onchip_rom|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_25(\onchip_rom|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_6(\onchip_rom|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\onchip_rom|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\onchip_rom|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\onchip_rom|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_3(\onchip_rom|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_rom|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_1(\onchip_rom|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_rom|the_altsyncram|auto_generated|q_a[17] ),
	.d_write(\nios2_qsys_0|d_write~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_rom_s1_agent_rsp_fifo|mem_used[1]~q ),
	.src2_valid(\mm_interconnect_0|cmd_demux_001|src2_valid~0_combout ),
	.src6_valid(\mm_interconnect_0|cmd_demux|src6_valid~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.hbreak_enabled(\nios2_qsys_0|hbreak_enabled~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_006|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_006|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_006|src_data[33]~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_006|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

Qsys_system_Qsys_system_onchip_ram onchip_ram(
	.q_a_4(\onchip_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_12(\onchip_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\onchip_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_0(\onchip_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\onchip_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\onchip_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_2(\onchip_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_18(\onchip_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_10(\onchip_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\onchip_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_5(\onchip_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\onchip_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\onchip_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_7(\onchip_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\onchip_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\onchip_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_9(\onchip_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_25(\onchip_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_6(\onchip_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\onchip_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\onchip_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\onchip_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_3(\onchip_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_1(\onchip_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_ram|the_altsyncram|auto_generated|q_a[17] ),
	.d_write(\nios2_qsys_0|d_write~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.src3_valid(\mm_interconnect_0|cmd_demux|src3_valid~1_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

Qsys_system_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.resetrequest(\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .lut_mask = 64'hFFFFEFFFFFFFFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .shared_arith = "off";

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \pio_key_export~input_o  = pio_key_export;

assign pio_led0_export = \pio_led|data_out~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\~GND~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDDFFFFFDFFDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'hEFDFDFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hF7FFFFF7FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|tdo~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFAAAAFFAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hFBFEFEFBFEFBFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hAAFFFFAAAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFFFDF8FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\jtag_uart_0|Qsys_system_jtag_uart_0_alt_jtag_atlantic|tdo~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.dataf(!\nios2_qsys_0|the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(gnd),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'hCCCCCCCCFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(gnd),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h3C3C3C3CFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(gnd),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'hC33CC33CFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'h69966996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'hFF9FFF6FFF9FFF6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFFFFBFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module Qsys_system_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	resetrequest,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
input 	resetrequest;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \merged_reset~0_combout ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


Qsys_system_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

Qsys_system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(\merged_reset~0_combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \merged_reset~0 (
	.dataa(!reset_reset_n),
	.datab(!resetrequest),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\merged_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_reset~0 .extended_lut = "off";
defparam \merged_reset~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \merged_reset~0 .shared_arith = "off";

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Qsys_system_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	merged_reset,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_jtag_uart_0 (
	q_b_4,
	Add1,
	q_b_0,
	Add11,
	q_b_2,
	Add12,
	q_b_5,
	Add13,
	q_b_7,
	q_b_6,
	Add14,
	q_b_3,
	Add15,
	q_b_1,
	Add16,
	tdo,
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	rst1,
	d_write,
	always2,
	d_address_line_field_0,
	Equal3,
	Equal31,
	d_address_offset_field_1,
	r_sync_rst,
	suppress_change_dest_id,
	av_waitrequest1,
	av_waitrequest2,
	mem_used_1,
	cp_valid,
	last_channel_0,
	read_latency_shift_reg,
	b_full,
	d_writedata_7,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	ien_AE1,
	av_readdata_9,
	ien_AF1,
	av_readdata_8,
	d_writedata_3,
	b_full1,
	d_writedata_1,
	read_01,
	d_writedata_4,
	d_writedata_2,
	d_writedata_10,
	ac1,
	d_writedata_5,
	rvalid1,
	d_writedata_6,
	woverflow1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	Add1;
output 	q_b_0;
output 	Add11;
output 	q_b_2;
output 	Add12;
output 	q_b_5;
output 	Add13;
output 	q_b_7;
output 	q_b_6;
output 	Add14;
output 	q_b_3;
output 	Add15;
output 	q_b_1;
output 	Add16;
output 	tdo;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
output 	rst1;
input 	d_write;
output 	always2;
input 	d_address_line_field_0;
input 	Equal3;
input 	Equal31;
input 	d_address_offset_field_1;
input 	r_sync_rst;
input 	suppress_change_dest_id;
output 	av_waitrequest1;
output 	av_waitrequest2;
input 	mem_used_1;
input 	cp_valid;
input 	last_channel_0;
input 	read_latency_shift_reg;
output 	b_full;
input 	d_writedata_7;
output 	b_non_empty;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	ien_AE1;
output 	av_readdata_9;
output 	ien_AF1;
output 	av_readdata_8;
input 	d_writedata_3;
output 	b_full1;
input 	d_writedata_1;
output 	read_01;
input 	d_writedata_4;
input 	d_writedata_2;
input 	d_writedata_10;
output 	ac1;
input 	d_writedata_5;
output 	rvalid1;
input 	d_writedata_6;
output 	woverflow1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \r_val~q ;
wire \fifo_wr~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|rvalid0~1_combout ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_rd~1_combout ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_ena~q ;
wire \fifo_wr~0_combout ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \wr_rfifo~combout ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_pause~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ;
wire \Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ;
wire \Add1~2 ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~22 ;
wire \Add1~26 ;
wire \av_waitrequest~1_combout ;
wire \ien_AE~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~0_combout ;
wire \fifo_rd~2_combout ;
wire \ac~0_combout ;
wire \rvalid~0_combout ;
wire \always2~1_combout ;
wire \woverflow~0_combout ;


Qsys_system_Qsys_system_jtag_uart_0_scfifo_r the_Qsys_system_jtag_uart_0_scfifo_r(
	.q_b_4(q_b_4),
	.q_b_0(q_b_0),
	.q_b_2(q_b_2),
	.q_b_5(q_b_5),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_1(q_b_1),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(\fifo_rd~0_combout ),
	.fifo_rd1(\fifo_rd~1_combout ),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_4(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_0(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_2(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_5(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_7(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_3(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_1(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_jtag_uart_0_scfifo_w the_Qsys_system_jtag_uart_0_scfifo_w(
	.q_b_7(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.fifo_wr(\fifo_wr~q ),
	.rvalid0(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|rvalid0~1_combout ),
	.b_non_empty(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.d_writedata_7(d_writedata_7),
	.d_writedata_3(d_writedata_3),
	.b_full(b_full1),
	.counter_reg_bit_3(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_5(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.d_writedata_1(d_writedata_1),
	.d_writedata_4(d_writedata_4),
	.d_writedata_2(d_writedata_2),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.clk_clk(clk_clk));

Qsys_system_alt_jtag_atlantic Qsys_system_jtag_uart_0_alt_jtag_atlantic(
	.r_dat({\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.tdo1(tdo),
	.rst11(rst1),
	.rst_n(r_sync_rst),
	.t_dav(\t_dav~q ),
	.r_val(\r_val~q ),
	.rvalid01(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|rvalid0~1_combout ),
	.t_ena1(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.t_pause1(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.wdata_4(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_0(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_2(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_5(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_7(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_3(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_1(\Qsys_system_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \r_val~0 (
	.dataa(!\Qsys_system_jtag_uart_0_alt_jtag_atlantic|rvalid0~1_combout ),
	.datab(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_val~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_val~0 .extended_lut = "off";
defparam \r_val~0 .lut_mask = 64'h7777777777777777;
defparam \r_val~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~1 (
	.dataa(!av_waitrequest1),
	.datab(!read_latency_shift_reg),
	.datac(!b_non_empty),
	.datad(!\fifo_rd~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~1 .extended_lut = "off";
defparam \fifo_rd~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \fifo_rd~1 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!b_full1),
	.datac(!\always2~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr~0 .extended_lut = "off";
defparam \fifo_wr~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \fifo_wr~0 .shared_arith = "off";

cyclonev_lcell_comb wr_rfifo(
	.dataa(!b_full),
	.datab(!\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_rfifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wr_rfifo.extended_lut = "off";
defparam wr_rfifo.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam wr_rfifo.shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add1),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add11),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add12),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add13),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add14),
	.cout(),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add15),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add16),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always2),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h7777777777777777;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_2),
	.datac(!d_address_line_field_0),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \av_waitrequest~0 .shared_arith = "off";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest2),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AE1),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclonev_lcell_comb \av_readdata[9] (
	.dataa(!\fifo_AE~q ),
	.datab(!ien_AE1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[9] .extended_lut = "off";
defparam \av_readdata[9] .lut_mask = 64'h7777777777777777;
defparam \av_readdata[9] .shared_arith = "off";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AF1),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cyclonev_lcell_comb \av_readdata[8]~0 (
	.dataa(!ien_AF1),
	.datab(!\pause_irq~q ),
	.datac(!\fifo_AF~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[8]~0 .extended_lut = "off";
defparam \av_readdata[8]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_readdata[8]~0 .shared_arith = "off";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!av_waitrequest1),
	.datab(!av_waitrequest2),
	.datac(!mem_used_1),
	.datad(!suppress_change_dest_id),
	.datae(!cp_valid),
	.dataf(!last_channel_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \ien_AE~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!always2),
	.datac(!av_waitrequest1),
	.datad(!av_waitrequest2),
	.datae(!mem_used_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ien_AE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ien_AE~0 .extended_lut = "off";
defparam \ien_AE~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \ien_AE~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datab(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datac(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datad(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!b_full1),
	.datab(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datac(!\the_Qsys_system_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datad(!\LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cyclonev_lcell_comb \pause_irq~0 (
	.dataa(!b_non_empty),
	.datab(!\pause_irq~q ),
	.datac(!\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.datad(!read_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pause_irq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pause_irq~0 .extended_lut = "off";
defparam \pause_irq~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \pause_irq~0 .shared_arith = "off";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(!counter_reg_bit_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000000000000000;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add0~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add0~9_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan1~1 .shared_arith = "off";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclonev_lcell_comb \fifo_rd~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!av_waitrequest2),
	.datac(!mem_used_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~0 .extended_lut = "off";
defparam \fifo_rd~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \fifo_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~2 (
	.dataa(!av_waitrequest1),
	.datab(!read_latency_shift_reg),
	.datac(!\fifo_rd~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~2 .extended_lut = "off";
defparam \fifo_rd~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \fifo_rd~2 .shared_arith = "off";

cyclonev_lcell_comb \ac~0 (
	.dataa(!\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.datab(!\ien_AE~0_combout ),
	.datac(!\Qsys_system_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.datad(!ac1),
	.datae(!d_writedata_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac~0 .extended_lut = "off";
defparam \ac~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \ac~0 .shared_arith = "off";

cyclonev_lcell_comb \rvalid~0 (
	.dataa(!b_non_empty),
	.datab(!\fifo_rd~2_combout ),
	.datac(!rvalid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~0 .extended_lut = "off";
defparam \rvalid~0 .lut_mask = 64'h4747474747474747;
defparam \rvalid~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~1 (
	.dataa(!always2),
	.datab(!av_waitrequest1),
	.datac(!av_waitrequest2),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \woverflow~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!b_full1),
	.datac(!\always2~1_combout ),
	.datad(!woverflow1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~0 .extended_lut = "off";
defparam \woverflow~0 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \woverflow~0 .shared_arith = "off";

endmodule

module Qsys_system_alt_jtag_atlantic (
	r_dat,
	tdo1,
	rst11,
	rst_n,
	t_dav,
	r_val,
	rvalid01,
	t_ena1,
	t_pause1,
	wdata_4,
	wdata_0,
	wdata_2,
	wdata_5,
	wdata_7,
	wdata_6,
	wdata_3,
	wdata_1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
output 	rst11;
input 	rst_n;
input 	t_dav;
input 	r_val;
output 	rvalid01;
output 	t_ena1;
output 	t_pause1;
output 	wdata_4;
output 	wdata_0;
output 	wdata_2;
output 	wdata_5;
output 	wdata_7;
output 	wdata_6;
output 	wdata_3;
output 	wdata_1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state~1_combout ;
wire \state~q ;
wire \td_shift[0]~2_combout ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[4]~q ;
wire \count[5]~q ;
wire \count[6]~q ;
wire \count[7]~q ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count[9]~_wirecell_combout ;
wire \count[0]~q ;
wire \count[1]~q ;
wire \state~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift[10]~q ;
wire \r_ena1~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~3_combout ;
wire \td_shift[9]~q ;
wire \td_shift~0_combout ;
wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~q ;
wire \td_shift~4_combout ;
wire \rdata[0]~q ;
wire \rdata[3]~q ;
wire \rdata[4]~q ;
wire \rdata[6]~q ;
wire \td_shift~12_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~11_combout ;
wire \td_shift[7]~q ;
wire \td_shift~10_combout ;
wire \td_shift[6]~q ;
wire \td_shift~9_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~8_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~7_combout ;
wire \td_shift[3]~q ;
wire \td_shift~6_combout ;
wire \td_shift[2]~q ;
wire \td_shift~5_combout ;
wire \td_shift[1]~q ;
wire \read_req~q ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \always2~0_combout ;
wire \rst2~q ;
wire \rvalid0~0_combout ;
wire \rvalid0~q ;
wire \rvalid~q ;
wire \td_shift~1_combout ;
wire \td_shift[0]~q ;
wire \write~1_combout ;
wire \write~0_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~1_combout ;
wire \write_valid~q ;
wire \t_ena~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \always2~2_combout ;
wire \t_pause~0_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

cyclonev_lcell_comb \rvalid0~1 (
	.dataa(!\rvalid0~q ),
	.datab(!\r_ena~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rvalid01),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~1 .extended_lut = "off";
defparam \rvalid0~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \rvalid0~1 .shared_arith = "off";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

cyclonev_lcell_comb \state~1 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!state_4),
	.datae(!\state~q ),
	.dataf(!altera_internal_jtag1),
	.datag(!irf_reg_0_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~1 .extended_lut = "on";
defparam \state~1 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \state~1 .shared_arith = "off";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclonev_lcell_comb \td_shift[0]~2 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift[0]~2 .extended_lut = "off";
defparam \td_shift[0]~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \td_shift[0]~2 .shared_arith = "off";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclonev_lcell_comb \count[9]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!altera_internal_jtag1),
	.datad(!state_4),
	.datae(!\count[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~0 .extended_lut = "off";
defparam \count[9]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \count[9]~0 .shared_arith = "off";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclonev_lcell_comb \count[9]~_wirecell (
	.dataa(!\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~_wirecell .extended_lut = "off";
defparam \count[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count[9]~_wirecell .shared_arith = "off";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count[9]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \state~0 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \state~0 .shared_arith = "off";

cyclonev_lcell_comb \user_saw_rvalid~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\td_shift[0]~q ),
	.datac(!\state~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\state~0_combout ),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_saw_rvalid~0 .extended_lut = "off";
defparam \user_saw_rvalid~0 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \user_saw_rvalid~0 .shared_arith = "off";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_ena1~q ),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

cyclonev_lcell_comb \r_ena~0 (
	.dataa(!r_val),
	.datab(!\r_ena1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_ena~0 .extended_lut = "off";
defparam \r_ena~0 .lut_mask = 64'h7777777777777777;
defparam \r_ena~0 .shared_arith = "off";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~3 (
	.dataa(!\count[9]~q ),
	.datab(!\td_shift[10]~q ),
	.datac(!\rdata[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~3 .extended_lut = "off";
defparam \td_shift~3 .lut_mask = 64'h2727272727272727;
defparam \td_shift~3 .shared_arith = "off";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclonev_lcell_comb \td_shift~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~0 .extended_lut = "off";
defparam \td_shift~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \td_shift~0 .shared_arith = "off";

cyclonev_lcell_comb \tck_t_dav~0 (
	.dataa(!t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tck_t_dav~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tck_t_dav~0 .extended_lut = "off";
defparam \tck_t_dav~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \tck_t_dav~0 .shared_arith = "off";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclonev_lcell_comb \write_stalled~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\tck_t_dav~q ),
	.datac(!\td_shift[10]~q ),
	.datad(!\write_stalled~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~0 .extended_lut = "off";
defparam \write_stalled~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \write_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \write_stalled~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!state_4),
	.datae(!splitter_nodes_receive_0_3),
	.dataf(!virtual_ir_scan_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~1 .extended_lut = "off";
defparam \write_stalled~1 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \write_stalled~1 .shared_arith = "off";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclonev_lcell_comb \td_shift~4 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~4 .extended_lut = "off";
defparam \td_shift~4 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \td_shift~4 .shared_arith = "off";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~12 (
	.dataa(!\td_shift[9]~q ),
	.datab(!\count[9]~q ),
	.datac(!\rdata[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~12 .extended_lut = "off";
defparam \td_shift~12 .lut_mask = 64'h4747474747474747;
defparam \td_shift~12 .shared_arith = "off";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclonev_lcell_comb \td_shift~11 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[8]~q ),
	.datae(!\rdata[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~11 .extended_lut = "off";
defparam \td_shift~11 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~11 .shared_arith = "off";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~10 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[4]~q ),
	.dataf(!\td_shift[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~10 .extended_lut = "off";
defparam \td_shift~10 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~10 .shared_arith = "off";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~9 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[3]~q ),
	.dataf(!\td_shift[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~9 .extended_lut = "off";
defparam \td_shift~9 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~9 .shared_arith = "off";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~8 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[5]~q ),
	.datae(!\rdata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~8 .extended_lut = "off";
defparam \td_shift~8 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~8 .shared_arith = "off";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclonev_lcell_comb \td_shift~7 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[4]~q ),
	.datae(!\rdata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~7 .extended_lut = "off";
defparam \td_shift~7 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~7 .shared_arith = "off";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~6 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[0]~q ),
	.dataf(!\td_shift[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~6 .extended_lut = "off";
defparam \td_shift~6 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~6 .shared_arith = "off";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~5 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\write_stalled~q ),
	.datae(!\td_shift~4_combout ),
	.dataf(!\td_shift[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~5 .extended_lut = "off";
defparam \td_shift~5 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \td_shift~5 .shared_arith = "off";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \read~0 .shared_arith = "off";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\read1~q ),
	.datab(!\read2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h6666666666666666;
defparam \always2~0 .shared_arith = "off";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclonev_lcell_comb \rvalid0~0 (
	.dataa(!\user_saw_rvalid~q ),
	.datab(!\rvalid0~q ),
	.datac(!\r_ena~0_combout ),
	.datad(!\read_req~q ),
	.datae(!\always2~0_combout ),
	.dataf(!\rst2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~0 .extended_lut = "off";
defparam \rvalid0~0 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \rvalid0~0 .shared_arith = "off";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid0~q ),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(\rvalid0~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \td_shift~1 (
	.dataa(!\state~q ),
	.datab(!\td_shift~0_combout ),
	.datac(!\tck_t_dav~q ),
	.datad(!\td_shift[1]~q ),
	.datae(!\count[9]~q ),
	.dataf(!\rvalid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~1 .extended_lut = "off";
defparam \td_shift~1 .lut_mask = 64'hBFFFEFFFFFFFFFFF;
defparam \td_shift~1 .shared_arith = "off";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclonev_lcell_comb \write~1 (
	.dataa(!\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!state_4),
	.datad(!splitter_nodes_receive_0_3),
	.datae(!virtual_ir_scan_reg),
	.dataf(!\count[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \write~0 .shared_arith = "off";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\write1~q ),
	.datab(!\write2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h6666666666666666;
defparam \always2~1 .shared_arith = "off";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclonev_lcell_comb \t_ena~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!t_ena1),
	.datae(!\always2~1_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_ena~0 .extended_lut = "off";
defparam \t_ena~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \t_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \jupdate~0 (
	.dataa(!irf_reg_0_1),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!\jupdate~q ),
	.datae(!state_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jupdate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jupdate~0 .extended_lut = "off";
defparam \jupdate~0 .lut_mask = 64'h9669699696696996;
defparam \jupdate~0 .shared_arith = "off";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclonev_lcell_comb \always2~2 (
	.dataa(!\jupdate1~q ),
	.datab(!\jupdate2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~2 .extended_lut = "off";
defparam \always2~2 .lut_mask = 64'h6666666666666666;
defparam \always2~2 .shared_arith = "off";

cyclonev_lcell_comb \t_pause~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!\always2~1_combout ),
	.datae(!\write_valid~q ),
	.dataf(!\always2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_pause~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_pause~0 .extended_lut = "off";
defparam \t_pause~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \t_pause~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_jtag_uart_0_scfifo_r (
	q_b_4,
	q_b_0,
	q_b_2,
	q_b_5,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_1,
	r_sync_rst,
	av_waitrequest,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	wdata_4,
	wdata_0,
	wdata_2,
	wdata_5,
	wdata_7,
	wdata_6,
	wdata_3,
	wdata_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_0;
output 	q_b_2;
output 	q_b_5;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_1;
input 	r_sync_rst;
input 	av_waitrequest;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	wdata_4;
input 	wdata_0;
input 	wdata_2;
input 	wdata_5;
input 	wdata_7;
input 	wdata_6;
input 	wdata_3;
input 	wdata_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module Qsys_system_scfifo_1 (
	q,
	r_sync_rst,
	av_waitrequest,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_scfifo_3291 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module Qsys_system_scfifo_3291 (
	q,
	r_sync_rst,
	av_waitrequest,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_a_dpfifo_5771 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module Qsys_system_a_dpfifo_5771 (
	q,
	r_sync_rst,
	av_waitrequest,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


Qsys_system_cntr_jgb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

Qsys_system_cntr_jgb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd1),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

Qsys_system_altsyncram_7pu1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd1),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

Qsys_system_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wreq),
	.clock(clock));

endmodule

module Qsys_system_a_fefifo_7cf (
	r_sync_rst,
	av_waitrequest,
	read_latency_shift_reg,
	b_full1,
	b_non_empty1,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	av_waitrequest;
input 	read_latency_shift_reg;
output 	b_full1;
output 	b_non_empty1;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \b_non_empty~0_combout ;


Qsys_system_cntr_vg7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wr_rfifo),
	._(\_~2_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~2 (
	.dataa(!av_waitrequest),
	.datab(!read_latency_shift_reg),
	.datac(!b_non_empty1),
	.datad(!fifo_rd),
	.datae(!wr_rfifo),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h9669699696696996;
defparam \_~2 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!b_non_empty1),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!counter_reg_bit_3),
	.datae(!counter_reg_bit_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!fifo_rd1),
	.datac(!counter_reg_bit_1),
	.datad(!counter_reg_bit_0),
	.datae(!t_ena),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \_~0 (
	.dataa(!counter_reg_bit_5),
	.datab(!counter_reg_bit_4),
	.datac(!counter_reg_bit_3),
	.datad(!wr_rfifo),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \_~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_0),
	.datad(!\_~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!b_full1),
	.datab(!b_non_empty1),
	.datac(!fifo_rd1),
	.datad(!t_ena),
	.datae(!\_~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hF7FFD5FFF7FFD5FF;
defparam \b_non_empty~0 .shared_arith = "off";

endmodule

module Qsys_system_cntr_vg7 (
	r_sync_rst,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_altsyncram_7pu1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_r:the_Qsys_system_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module Qsys_system_cntr_jgb (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_cntr_jgb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_jtag_uart_0_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	fifo_wr,
	rvalid0,
	b_non_empty,
	r_val,
	d_writedata_7,
	d_writedata_3,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	d_writedata_1,
	d_writedata_4,
	d_writedata_2,
	d_writedata_5,
	d_writedata_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	fifo_wr;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
input 	d_writedata_7;
input 	d_writedata_3;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	d_writedata_1;
input 	d_writedata_4;
input 	d_writedata_2;
input 	d_writedata_5;
input 	d_writedata_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.wrreq(fifo_wr),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clk_clk));

endmodule

module Qsys_system_scfifo_2 (
	q,
	data,
	r_sync_rst,
	wrreq,
	rvalid0,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wrreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_scfifo_3291_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.wrreq(wrreq),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module Qsys_system_scfifo_3291_1 (
	q,
	data,
	r_sync_rst,
	wrreq,
	rvalid0,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wrreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_a_dpfifo_5771_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.wreq(wrreq),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module Qsys_system_a_dpfifo_5771_1 (
	q,
	data,
	r_sync_rst,
	wreq,
	rvalid0,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


Qsys_system_cntr_jgb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

Qsys_system_cntr_jgb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

Qsys_system_altsyncram_7pu1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.clocken1(r_val),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

Qsys_system_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.rvalid0(rvalid0),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.b_full1(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module Qsys_system_a_fefifo_7cf_1 (
	r_sync_rst,
	fifo_wr,
	rvalid0,
	b_non_empty1,
	r_val,
	b_full1,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
input 	rvalid0;
output 	b_non_empty1;
input 	r_val;
output 	b_full1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;


Qsys_system_cntr_vg7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(fifo_wr),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!rvalid0),
	.datab(!fifo_wr),
	.datac(!b_non_empty1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h9696969696969696;
defparam \_~0 .shared_arith = "off";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \b_non_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~1 (
	.dataa(!r_val),
	.datab(!counter_reg_bit_3),
	.datac(!counter_reg_bit_0),
	.datad(!\b_non_empty~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~1 .extended_lut = "off";
defparam \b_non_empty~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \b_non_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~2 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!b_full1),
	.datad(!\b_non_empty~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~2 .extended_lut = "off";
defparam \b_non_empty~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \b_non_empty~2 .shared_arith = "off";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_5),
	.datae(!counter_reg_bit_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!r_val),
	.datab(!b_full1),
	.datac(!counter_reg_bit_0),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_1),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

endmodule

module Qsys_system_cntr_vg7_1 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_altsyncram_7pu1_1 (
	q_b,
	data_a,
	wren_a,
	clocken1,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	wren_a;
input 	clocken1;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Qsys_system_jtag_uart_0:jtag_uart_0|Qsys_system_jtag_uart_0_scfifo_w:the_Qsys_system_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module Qsys_system_cntr_jgb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_cntr_jgb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0 (
	q_a_4,
	q_a_41,
	q_a_20,
	q_a_201,
	q_a_12,
	q_a_121,
	q_a_28,
	q_a_281,
	q_a_0,
	q_a_01,
	q_a_16,
	q_a_161,
	q_a_8,
	q_a_81,
	q_a_24,
	q_a_241,
	q_a_2,
	q_a_21,
	q_a_18,
	q_a_181,
	q_a_10,
	q_a_101,
	q_a_26,
	q_a_261,
	q_a_5,
	q_a_51,
	q_a_211,
	q_a_212,
	q_a_13,
	q_a_131,
	q_a_29,
	q_a_291,
	q_a_7,
	q_a_71,
	q_a_23,
	q_a_231,
	q_a_15,
	q_a_151,
	q_a_31,
	q_a_311,
	q_a_11,
	q_a_111,
	q_a_27,
	q_a_271,
	q_a_9,
	q_a_91,
	q_a_25,
	q_a_251,
	q_a_6,
	q_a_61,
	q_a_22,
	q_a_221,
	q_a_14,
	q_a_141,
	q_a_30,
	q_a_301,
	q_a_3,
	q_a_32,
	q_a_19,
	q_a_191,
	q_a_1,
	q_a_17,
	q_a_171,
	q_a_172,
	q_b_4,
	readdata_4,
	Add1,
	readdata_20,
	readdata_12,
	readdata_28,
	q_b_0,
	Add11,
	readdata_16,
	readdata_8,
	readdata_24,
	q_b_2,
	readdata_2,
	Add12,
	readdata_18,
	readdata_10,
	readdata_26,
	q_b_5,
	readdata_5,
	Add13,
	readdata_21,
	readdata_13,
	readdata_29,
	q_b_7,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_11,
	readdata_27,
	readdata_9,
	readdata_25,
	q_b_6,
	readdata_6,
	Add14,
	readdata_22,
	readdata_14,
	readdata_30,
	q_b_3,
	readdata_3,
	Add15,
	readdata_19,
	q_b_1,
	Add16,
	readdata_17,
	WideOr0,
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	rst1,
	d_write,
	always2,
	d_address_line_field_0,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	Equal3,
	d_address_line_field_1,
	d_address_tag_field_5,
	d_address_tag_field_4,
	d_address_tag_field_3,
	d_address_tag_field_2,
	Equal31,
	m0_write,
	d_address_offset_field_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	r_sync_rst,
	d_read,
	av_begintransfer,
	suppress_change_dest_id,
	av_waitrequest,
	Equal4,
	suppress_change_dest_id1,
	mem_used_1,
	wait_latency_counter_11,
	wait_latency_counter_01,
	saved_grant_0,
	mem_used_11,
	av_waitrequest1,
	mem_used_12,
	saved_grant_01,
	waitrequest,
	mem_used_13,
	saved_grant_02,
	mem_used_14,
	WideOr01,
	av_waitrequest2,
	cp_valid,
	WideOr1,
	has_pending_responses,
	i_read,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	src1_valid,
	src3_valid,
	saved_grant_1,
	last_channel_0,
	read_latency_shift_reg,
	WideOr11,
	rf_source_valid,
	src2_valid,
	src6_valid,
	saved_grant_11,
	hbreak_enabled,
	save_dest_id,
	nonposted_cmd_accepted,
	suppress_change_dest_id2,
	ic_fill_line_5,
	src_data_46,
	b_full,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	d_writedata_7,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_payload1,
	d_byteenable_0,
	src_data_32,
	WideOr12,
	ien_AE,
	av_readdata_9,
	ien_AF,
	av_readdata_8,
	d_writedata_3,
	src_payload2,
	src_data_4,
	src_data_20,
	src_data_12,
	src_data_28,
	src_data_0,
	src_data_16,
	src_data_8,
	src_data_24,
	src_data_2,
	src_data_18,
	src_data_10,
	src_data_26,
	src_data_5,
	src_data_21,
	src_data_13,
	src_data_29,
	src_data_7,
	src_data_23,
	src_data_15,
	src_data_31,
	src_data_11,
	src_data_27,
	src_data_9,
	src_data_25,
	src_data_6,
	src_data_22,
	src_data_14,
	src_data_30,
	src_data_3,
	src_data_19,
	b_full1,
	d_writedata_1,
	src_payload3,
	read_0,
	src_data_51,
	src_data_33,
	src_data_1,
	src_data_47,
	src_data_210,
	src_data_281,
	src_data_301,
	src_data_311,
	src_data_271,
	src_data_291,
	src_data_01,
	src_data_231,
	src_data_251,
	src_data_261,
	src_data_221,
	src_data_241,
	src_data_17,
	src_data_171,
	src_data_161,
	src_data_151,
	src_data_131,
	src_data_141,
	src_data_121,
	src_data_111,
	src_data_101,
	d_writedata_4,
	src_payload4,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_461,
	src_data_471,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_321,
	src_payload5,
	src_data_382,
	src_data_392,
	src_data_402,
	src_data_412,
	src_data_422,
	src_data_432,
	src_data_442,
	src_data_452,
	src_data_462,
	src_data_472,
	src_data_481,
	src_data_491,
	src_data_322,
	d_writedata_20,
	src_payload6,
	d_byteenable_2,
	src_data_34,
	src_payload7,
	src_data_341,
	d_writedata_12,
	src_payload8,
	d_byteenable_1,
	src_data_331,
	src_payload9,
	src_data_332,
	d_writedata_28,
	src_payload10,
	d_byteenable_3,
	src_data_35,
	src_payload11,
	src_data_351,
	src_payload12,
	src_payload13,
	readdata_0,
	readdata_01,
	readdata_02,
	d_writedata_16,
	src_payload14,
	src_payload15,
	d_writedata_8,
	src_payload16,
	src_payload17,
	d_writedata_24,
	src_payload18,
	src_payload19,
	src_data_81,
	d_writedata_2,
	src_payload20,
	src_payload21,
	d_writedata_18,
	src_payload22,
	src_payload23,
	d_writedata_10,
	src_payload24,
	src_payload25,
	ac,
	d_writedata_26,
	src_payload26,
	src_payload27,
	d_writedata_5,
	src_payload28,
	src_payload29,
	d_writedata_21,
	src_payload30,
	src_payload31,
	d_writedata_13,
	src_payload32,
	src_payload33,
	d_writedata_29,
	src_payload34,
	src_payload35,
	src_data_181,
	src_payload36,
	src_payload37,
	d_writedata_23,
	src_payload38,
	src_payload39,
	d_writedata_15,
	src_payload40,
	src_payload41,
	rvalid,
	d_writedata_31,
	src_payload42,
	src_payload43,
	src_data_172,
	d_writedata_11,
	src_payload44,
	src_payload45,
	d_writedata_27,
	src_payload46,
	src_payload47,
	d_writedata_9,
	src_payload48,
	src_payload49,
	d_writedata_25,
	src_payload50,
	src_payload51,
	d_writedata_6,
	src_payload52,
	src_payload53,
	d_writedata_22,
	src_payload54,
	src_payload55,
	d_writedata_14,
	src_payload56,
	src_payload57,
	woverflow,
	d_writedata_30,
	src_payload58,
	src_payload59,
	src_data_211,
	src_data_61,
	src_data_201,
	src_data_191,
	src_data_91,
	src_payload60,
	src_payload61,
	d_writedata_19,
	src_payload62,
	src_payload63,
	src_payload64,
	readdata_1,
	src_payload65,
	src_payload66,
	src_data_71,
	d_writedata_17,
	src_payload67,
	src_payload68,
	src_payload69,
	src_data_342,
	src_payload70,
	src_payload71,
	src_payload72,
	src_data_352,
	src_payload73,
	src_payload74,
	src_payload75,
	src_payload76,
	src_payload77,
	src_payload78,
	src_payload79,
	src_payload80,
	src_data_333,
	src_payload81,
	src_payload82,
	src_payload83,
	src_payload84,
	src_payload85,
	src_payload86,
	src_payload87,
	src_payload88,
	src_payload89,
	src_payload90,
	src_payload91,
	src_payload92,
	src_payload93,
	src_payload94,
	src_payload95,
	src_payload96,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	q_a_4;
input 	q_a_41;
input 	q_a_20;
input 	q_a_201;
input 	q_a_12;
input 	q_a_121;
input 	q_a_28;
input 	q_a_281;
input 	q_a_0;
input 	q_a_01;
input 	q_a_16;
input 	q_a_161;
input 	q_a_8;
input 	q_a_81;
input 	q_a_24;
input 	q_a_241;
input 	q_a_2;
input 	q_a_21;
input 	q_a_18;
input 	q_a_181;
input 	q_a_10;
input 	q_a_101;
input 	q_a_26;
input 	q_a_261;
input 	q_a_5;
input 	q_a_51;
input 	q_a_211;
input 	q_a_212;
input 	q_a_13;
input 	q_a_131;
input 	q_a_29;
input 	q_a_291;
input 	q_a_7;
input 	q_a_71;
input 	q_a_23;
input 	q_a_231;
input 	q_a_15;
input 	q_a_151;
input 	q_a_31;
input 	q_a_311;
input 	q_a_11;
input 	q_a_111;
input 	q_a_27;
input 	q_a_271;
input 	q_a_9;
input 	q_a_91;
input 	q_a_25;
input 	q_a_251;
input 	q_a_6;
input 	q_a_61;
input 	q_a_22;
input 	q_a_221;
input 	q_a_14;
input 	q_a_141;
input 	q_a_30;
input 	q_a_301;
input 	q_a_3;
input 	q_a_32;
input 	q_a_19;
input 	q_a_191;
input 	q_a_1;
input 	q_a_17;
input 	q_a_171;
input 	q_a_172;
input 	q_b_4;
input 	readdata_4;
input 	Add1;
input 	readdata_20;
input 	readdata_12;
input 	readdata_28;
input 	q_b_0;
input 	Add11;
input 	readdata_16;
input 	readdata_8;
input 	readdata_24;
input 	q_b_2;
input 	readdata_2;
input 	Add12;
input 	readdata_18;
input 	readdata_10;
input 	readdata_26;
input 	q_b_5;
input 	readdata_5;
input 	Add13;
input 	readdata_21;
input 	readdata_13;
input 	readdata_29;
input 	q_b_7;
input 	readdata_7;
input 	readdata_23;
input 	readdata_15;
input 	readdata_31;
input 	readdata_11;
input 	readdata_27;
input 	readdata_9;
input 	readdata_25;
input 	q_b_6;
input 	readdata_6;
input 	Add14;
input 	readdata_22;
input 	readdata_14;
input 	readdata_30;
input 	q_b_3;
input 	readdata_3;
input 	Add15;
input 	readdata_19;
input 	q_b_1;
input 	Add16;
input 	readdata_17;
output 	WideOr0;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	rst1;
input 	d_write;
input 	always2;
input 	d_address_line_field_0;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
output 	Equal3;
input 	d_address_line_field_1;
input 	d_address_tag_field_5;
input 	d_address_tag_field_4;
input 	d_address_tag_field_3;
input 	d_address_tag_field_2;
output 	Equal31;
output 	m0_write;
input 	d_address_offset_field_1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	r_sync_rst;
input 	d_read;
output 	av_begintransfer;
output 	suppress_change_dest_id;
input 	av_waitrequest;
output 	Equal4;
output 	suppress_change_dest_id1;
output 	mem_used_1;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
output 	saved_grant_0;
output 	mem_used_11;
input 	av_waitrequest1;
output 	mem_used_12;
output 	saved_grant_01;
input 	waitrequest;
output 	mem_used_13;
output 	saved_grant_02;
output 	mem_used_14;
output 	WideOr01;
output 	av_waitrequest2;
output 	cp_valid;
output 	WideOr1;
output 	has_pending_responses;
input 	i_read;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
output 	src1_valid;
output 	src3_valid;
output 	saved_grant_1;
output 	last_channel_0;
output 	read_latency_shift_reg;
output 	WideOr11;
output 	rf_source_valid;
output 	src2_valid;
output 	src6_valid;
output 	saved_grant_11;
input 	hbreak_enabled;
output 	save_dest_id;
output 	nonposted_cmd_accepted;
output 	suppress_change_dest_id2;
input 	ic_fill_line_5;
output 	src_data_46;
input 	b_full;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_0;
input 	d_writedata_7;
input 	b_non_empty;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
output 	src_data_45;
output 	src_data_44;
output 	src_data_43;
output 	src_data_42;
output 	src_payload1;
input 	d_byteenable_0;
output 	src_data_32;
output 	WideOr12;
input 	ien_AE;
input 	av_readdata_9;
input 	ien_AF;
input 	av_readdata_8;
input 	d_writedata_3;
output 	src_payload2;
output 	src_data_4;
output 	src_data_20;
output 	src_data_12;
output 	src_data_28;
output 	src_data_0;
output 	src_data_16;
output 	src_data_8;
output 	src_data_24;
output 	src_data_2;
output 	src_data_18;
output 	src_data_10;
output 	src_data_26;
output 	src_data_5;
output 	src_data_21;
output 	src_data_13;
output 	src_data_29;
output 	src_data_7;
output 	src_data_23;
output 	src_data_15;
output 	src_data_31;
output 	src_data_11;
output 	src_data_27;
output 	src_data_9;
output 	src_data_25;
output 	src_data_6;
output 	src_data_22;
output 	src_data_14;
output 	src_data_30;
output 	src_data_3;
output 	src_data_19;
input 	b_full1;
input 	d_writedata_1;
output 	src_payload3;
input 	read_0;
output 	src_data_51;
output 	src_data_33;
output 	src_data_1;
output 	src_data_47;
output 	src_data_210;
output 	src_data_281;
output 	src_data_301;
output 	src_data_311;
output 	src_data_271;
output 	src_data_291;
output 	src_data_01;
output 	src_data_231;
output 	src_data_251;
output 	src_data_261;
output 	src_data_221;
output 	src_data_241;
output 	src_data_17;
output 	src_data_171;
output 	src_data_161;
output 	src_data_151;
output 	src_data_131;
output 	src_data_141;
output 	src_data_121;
output 	src_data_111;
output 	src_data_101;
input 	d_writedata_4;
output 	src_payload4;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_461;
output 	src_data_471;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_321;
output 	src_payload5;
output 	src_data_382;
output 	src_data_392;
output 	src_data_402;
output 	src_data_412;
output 	src_data_422;
output 	src_data_432;
output 	src_data_442;
output 	src_data_452;
output 	src_data_462;
output 	src_data_472;
output 	src_data_481;
output 	src_data_491;
output 	src_data_322;
input 	d_writedata_20;
output 	src_payload6;
input 	d_byteenable_2;
output 	src_data_34;
output 	src_payload7;
output 	src_data_341;
input 	d_writedata_12;
output 	src_payload8;
input 	d_byteenable_1;
output 	src_data_331;
output 	src_payload9;
output 	src_data_332;
input 	d_writedata_28;
output 	src_payload10;
input 	d_byteenable_3;
output 	src_data_35;
output 	src_payload11;
output 	src_data_351;
output 	src_payload12;
output 	src_payload13;
input 	readdata_0;
input 	readdata_01;
input 	readdata_02;
input 	d_writedata_16;
output 	src_payload14;
output 	src_payload15;
input 	d_writedata_8;
output 	src_payload16;
output 	src_payload17;
input 	d_writedata_24;
output 	src_payload18;
output 	src_payload19;
output 	src_data_81;
input 	d_writedata_2;
output 	src_payload20;
output 	src_payload21;
input 	d_writedata_18;
output 	src_payload22;
output 	src_payload23;
input 	d_writedata_10;
output 	src_payload24;
output 	src_payload25;
input 	ac;
input 	d_writedata_26;
output 	src_payload26;
output 	src_payload27;
input 	d_writedata_5;
output 	src_payload28;
output 	src_payload29;
input 	d_writedata_21;
output 	src_payload30;
output 	src_payload31;
input 	d_writedata_13;
output 	src_payload32;
output 	src_payload33;
input 	d_writedata_29;
output 	src_payload34;
output 	src_payload35;
output 	src_data_181;
output 	src_payload36;
output 	src_payload37;
input 	d_writedata_23;
output 	src_payload38;
output 	src_payload39;
input 	d_writedata_15;
output 	src_payload40;
output 	src_payload41;
input 	rvalid;
input 	d_writedata_31;
output 	src_payload42;
output 	src_payload43;
output 	src_data_172;
input 	d_writedata_11;
output 	src_payload44;
output 	src_payload45;
input 	d_writedata_27;
output 	src_payload46;
output 	src_payload47;
input 	d_writedata_9;
output 	src_payload48;
output 	src_payload49;
input 	d_writedata_25;
output 	src_payload50;
output 	src_payload51;
input 	d_writedata_6;
output 	src_payload52;
output 	src_payload53;
input 	d_writedata_22;
output 	src_payload54;
output 	src_payload55;
input 	d_writedata_14;
output 	src_payload56;
output 	src_payload57;
input 	woverflow;
input 	d_writedata_30;
output 	src_payload58;
output 	src_payload59;
output 	src_data_211;
output 	src_data_61;
output 	src_data_201;
output 	src_data_191;
output 	src_data_91;
output 	src_payload60;
output 	src_payload61;
input 	d_writedata_19;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
input 	readdata_1;
output 	src_payload65;
output 	src_payload66;
output 	src_data_71;
input 	d_writedata_17;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_data_342;
output 	src_payload70;
output 	src_payload71;
output 	src_payload72;
output 	src_data_352;
output 	src_payload73;
output 	src_payload74;
output 	src_payload75;
output 	src_payload76;
output 	src_payload77;
output 	src_payload78;
output 	src_payload79;
output 	src_payload80;
output 	src_data_333;
output 	src_payload81;
output 	src_payload82;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_payload86;
output 	src_payload87;
output 	src_payload88;
output 	src_payload89;
output 	src_payload90;
output 	src_payload91;
output 	src_payload92;
output 	src_payload93;
output 	src_payload94;
output 	src_payload95;
output 	src_payload96;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \pio_led_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \nios2_qsys_0_data_master_limiter|has_pending_responses~q ;
wire \router|always1~0_combout ;
wire \router|Equal2~0_combout ;
wire \router|src_data[77]~0_combout ;
wire \router|Equal1~0_combout ;
wire \router|src_data[77]~1_combout ;
wire \router|src_data[79]~2_combout ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ;
wire \sysid_qsys_0_control_slave_translator|wait_latency_counter[0]~q ;
wire \router|src_channel[3]~0_combout ;
wire \router|Equal3~2_combout ;
wire \cmd_demux_001|sink_ready~0_combout ;
wire \onchip_rom_s1_translator|read_latency_shift_reg~0_combout ;
wire \pio_led_s1_translator|read_latency_shift_reg[0]~q ;
wire \nios2_qsys_0_data_master_limiter|last_channel[4]~q ;
wire \pio_led_s1_translator|read_latency_shift_reg~1_combout ;
wire \onchip_ram_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_ram_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_ram_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_003|src0_valid~0_combout ;
wire \onchip_rom_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_rom_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_rom_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_006|src0_valid~0_combout ;
wire \onchip_ram_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \onchip_rom_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_002|src0_valid~0_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \pio_key_s1_translator|read_latency_shift_reg[0]~q ;
wire \pio_led_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][61]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][61]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ;
wire \pio_key_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \router|src_data[78]~3_combout ;
wire \sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ;
wire \nios2_qsys_0_data_master_limiter|last_channel[1]~q ;
wire \sysid_qsys_0_control_slave_agent|m0_write~0_combout ;
wire \nios2_qsys_0_data_master_limiter|last_channel[5]~q ;
wire \pio_key_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \nios2_qsys_0_instruction_master_limiter|last_channel[1]~q ;
wire \router_001|src_channel[1]~0_combout ;
wire \nios2_qsys_0_data_master_limiter|last_channel[3]~q ;
wire \onchip_ram_s1_translator|read_latency_shift_reg~0_combout ;
wire \onchip_ram_s1_agent|rf_source_valid~0_combout ;
wire \router_001|Equal2~0_combout ;
wire \nios2_qsys_0_instruction_master_limiter|last_channel[0]~q ;
wire \cmd_demux_001|src0_valid~1_combout ;
wire \cmd_demux_001|src0_valid~2_combout ;
wire \nios2_qsys_0_data_master_limiter|last_channel[2]~q ;
wire \cmd_demux|src2_valid~0_combout ;
wire \cmd_demux|src2_valid~1_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \router_001|Equal1~0_combout ;
wire \nios2_qsys_0_instruction_master_limiter|last_channel[2]~q ;
wire \nios2_qsys_0_data_master_limiter|last_channel[6]~q ;
wire \onchip_rom_s1_agent|rf_source_valid~0_combout ;
wire \onchip_ram_s1_translator|read_latency_shift_reg~1_combout ;
wire \onchip_rom_s1_translator|read_latency_shift_reg~1_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ;
wire \pio_key_s1_translator|read_latency_shift_reg~1_combout ;
wire \onchip_rom_s1_agent_rsp_fifo|mem~3_combout ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \rsp_demux_003|src1_valid~0_combout ;
wire \rsp_demux_006|src1_valid~0_combout ;
wire \sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ;
wire \pio_key_s1_translator|av_readdata_pre[0]~q ;
wire \pio_led_s1_translator|av_readdata_pre[0]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ;


Qsys_system_altera_merlin_master_agent nios2_qsys_0_data_master_agent(
	.rst1(rst1),
	.d_write(d_write),
	.d_read(d_read),
	.suppress_change_dest_id(suppress_change_dest_id1),
	.WideOr0(WideOr01),
	.av_waitrequest1(av_waitrequest2),
	.cp_valid(cp_valid));

Qsys_system_altera_merlin_slave_translator_3 onchip_rom_s1_translator(
	.rst1(rst1),
	.reset(r_sync_rst),
	.mem_used_1(mem_used_14),
	.read_latency_shift_reg(\onchip_rom_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(\onchip_rom_s1_translator|read_latency_shift_reg[0]~q ),
	.rf_source_valid(\onchip_rom_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg1(\onchip_rom_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator_4 pio_key_s1_translator(
	.rst1(rst1),
	.d_write(d_write),
	.reset(r_sync_rst),
	.d_read(d_read),
	.av_begintransfer(av_begintransfer),
	.suppress_change_dest_id(suppress_change_dest_id),
	.Equal4(Equal4),
	.mem_used_1(mem_used_1),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(\pio_key_s1_translator|read_latency_shift_reg[0]~q ),
	.last_channel_5(\nios2_qsys_0_data_master_limiter|last_channel[5]~q ),
	.read_latency_shift_reg(\pio_key_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg1(\pio_key_s1_translator|read_latency_shift_reg~1_combout ),
	.av_readdata_pre_0(\pio_key_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_01}),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator_5 pio_led_s1_translator(
	.rst1(rst1),
	.always2(always2),
	.mem_used_1(\pio_led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(m0_write),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.reset(r_sync_rst),
	.d_read(d_read),
	.suppress_change_dest_id(suppress_change_dest_id),
	.Equal3(\router|Equal3~2_combout ),
	.read_latency_shift_reg_0(\pio_led_s1_translator|read_latency_shift_reg[0]~q ),
	.last_channel_4(\nios2_qsys_0_data_master_limiter|last_channel[4]~q ),
	.read_latency_shift_reg(\pio_led_s1_translator|read_latency_shift_reg~1_combout ),
	.cp_valid(cp_valid),
	.av_readdata_pre_0(\pio_led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_02}),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator_2 onchip_ram_s1_translator(
	.rst1(rst1),
	.reset(r_sync_rst),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\onchip_ram_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~0_combout ),
	.rf_source_valid(\onchip_ram_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg1(\onchip_ram_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator_1 nios2_qsys_0_jtag_debug_module_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.rst1(rst1),
	.reset(r_sync_rst),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.rf_source_valid(rf_source_valid),
	.av_readdata_pre_4(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_12(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_0(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_8(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_2(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_10(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_5(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_13(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_7(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_9(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_6(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_14(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_30(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_3(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_1(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator_6 sysid_qsys_0_control_slave_translator(
	.av_readdata({gnd,d_address_offset_field_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rst1(rst1),
	.d_write(d_write),
	.reset(r_sync_rst),
	.d_read(d_read),
	.av_begintransfer(av_begintransfer),
	.suppress_change_dest_id(suppress_change_dest_id),
	.always1(\router|always1~0_combout ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sysid_qsys_0_control_slave_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.av_waitrequest_generated(\sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ),
	.last_channel_1(\nios2_qsys_0_data_master_limiter|last_channel[1]~q ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_30(\sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_translator jtag_uart_0_avalon_jtag_slave_translator(
	.av_readdata_pre_4(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_2(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_5(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_7(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_3(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_1(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.q_b_4(q_b_4),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Add14,Add13,Add1,Add15,Add12,Add16,Add11,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,GND_port,GND_port,GND_port,GND_port,GND_port,GND_port,ien_AE,ien_AF}),
	.q_b_0(q_b_0),
	.q_b_2(q_b_2),
	.q_b_5(q_b_5),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_1(q_b_1),
	.rst1(rst1),
	.reset(r_sync_rst),
	.d_read(d_read),
	.suppress_change_dest_id(suppress_change_dest_id),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.last_channel_0(last_channel_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg1(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ),
	.b_full(b_full),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.av_readdata_pre_12(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_8(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_10(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_13(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_15(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_9(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_14(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.b_full1(b_full1),
	.read_0(read_0),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_agent_2 onchip_ram_s1_agent(
	.d_read(d_read),
	.saved_grant_0(saved_grant_0),
	.i_read(i_read),
	.src1_valid(src1_valid),
	.src3_valid(src3_valid),
	.saved_grant_1(saved_grant_1),
	.rf_source_valid(\onchip_ram_s1_agent|rf_source_valid~0_combout ));

Qsys_system_altera_avalon_sc_fifo_1 nios2_qsys_0_jtag_debug_module_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_read(d_read),
	.saved_grant_0(saved_grant_01),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ),
	.mem_61_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ),
	.i_read(i_read),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.rf_source_valid(rf_source_valid),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_agent_1 nios2_qsys_0_jtag_debug_module_agent(
	.d_read(d_read),
	.saved_grant_0(saved_grant_01),
	.i_read(i_read),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.WideOr1(WideOr11),
	.rf_source_valid(rf_source_valid));

Qsys_system_altera_avalon_sc_fifo_6 sysid_qsys_0_control_slave_agent_rsp_fifo(
	.rst1(rst1),
	.reset(r_sync_rst),
	.suppress_change_dest_id(suppress_change_dest_id),
	.always1(\router|always1~0_combout ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_61_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][61]~q ),
	.av_waitrequest_generated(\sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ),
	.last_channel_1(\nios2_qsys_0_data_master_limiter|last_channel[1]~q ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_agent_6 sysid_qsys_0_control_slave_agent(
	.rst1(rst1),
	.always1(\router|always1~0_combout ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ));

Qsys_system_altera_avalon_sc_fifo jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_61_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][61]~q ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg1(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

Qsys_system_Qsys_system_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_4(q_a_4),
	.q_a_41(q_a_41),
	.q_a_20(q_a_20),
	.q_a_201(q_a_201),
	.q_a_12(q_a_12),
	.q_a_121(q_a_121),
	.q_a_28(q_a_28),
	.q_a_281(q_a_281),
	.q_a_0(q_a_0),
	.q_a_01(q_a_01),
	.q_a_16(q_a_16),
	.q_a_161(q_a_161),
	.q_a_8(q_a_8),
	.q_a_81(q_a_81),
	.q_a_24(q_a_24),
	.q_a_241(q_a_241),
	.q_a_2(q_a_2),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.q_a_181(q_a_181),
	.q_a_10(q_a_10),
	.q_a_101(q_a_101),
	.q_a_26(q_a_26),
	.q_a_261(q_a_261),
	.q_a_5(q_a_5),
	.q_a_51(q_a_51),
	.q_a_211(q_a_211),
	.q_a_212(q_a_212),
	.q_a_13(q_a_13),
	.q_a_131(q_a_131),
	.q_a_29(q_a_29),
	.q_a_291(q_a_291),
	.q_a_7(q_a_7),
	.q_a_71(q_a_71),
	.q_a_23(q_a_23),
	.q_a_231(q_a_231),
	.q_a_15(q_a_15),
	.q_a_151(q_a_151),
	.q_a_31(q_a_31),
	.q_a_311(q_a_311),
	.q_a_11(q_a_11),
	.q_a_111(q_a_111),
	.q_a_27(q_a_27),
	.q_a_271(q_a_271),
	.q_a_9(q_a_9),
	.q_a_91(q_a_91),
	.q_a_25(q_a_25),
	.q_a_251(q_a_251),
	.q_a_6(q_a_6),
	.q_a_61(q_a_61),
	.q_a_22(q_a_22),
	.q_a_221(q_a_221),
	.q_a_14(q_a_14),
	.q_a_141(q_a_141),
	.q_a_30(q_a_30),
	.q_a_301(q_a_301),
	.q_a_3(q_a_3),
	.q_a_32(q_a_32),
	.q_a_19(q_a_19),
	.q_a_191(q_a_191),
	.q_a_1(q_a_1),
	.q_a_17(q_a_17),
	.q_a_171(q_a_171),
	.q_a_172(q_a_172),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.src1_valid2(\rsp_demux_006|src1_valid~0_combout ),
	.WideOr11(WideOr12),
	.av_readdata_pre_4(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_12(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_0(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_8(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_2(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_10(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_5(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_13(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_7(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_9(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_6(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_14(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_30(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_3(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.src_data_5(src_data_51),
	.src_data_3(src_data_33),
	.av_readdata_pre_1(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.src_data_4(src_data_47),
	.src_data_2(src_data_210),
	.src_data_28(src_data_281),
	.src_data_30(src_data_301),
	.src_data_31(src_data_311),
	.src_data_27(src_data_271),
	.src_data_29(src_data_291),
	.src_data_0(src_data_01),
	.src_data_23(src_data_231),
	.src_data_25(src_data_251),
	.src_data_26(src_data_261),
	.src_data_22(src_data_221),
	.src_data_24(src_data_241),
	.av_readdata_pre_17(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.src_data_16(src_data_161),
	.src_data_15(src_data_151),
	.src_data_13(src_data_131),
	.src_data_14(src_data_141),
	.src_data_12(src_data_121),
	.src_data_11(src_data_111),
	.src_data_10(src_data_101),
	.src_data_8(src_data_81),
	.src_data_18(src_data_181),
	.src_data_17(src_data_172),
	.src_data_21(src_data_211),
	.src_data_6(src_data_61),
	.src_data_20(src_data_201),
	.src_data_19(src_data_191),
	.src_data_9(src_data_91),
	.src_data_7(src_data_71));

Qsys_system_Qsys_system_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_4(q_a_4),
	.q_a_41(q_a_41),
	.av_readdata_pre_4(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.q_a_20(q_a_20),
	.q_a_201(q_a_201),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_12(q_a_12),
	.q_a_121(q_a_121),
	.q_a_28(q_a_28),
	.q_a_281(q_a_281),
	.q_a_0(q_a_0),
	.q_a_01(q_a_01),
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.q_a_16(q_a_16),
	.q_a_161(q_a_161),
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_a_8(q_a_8),
	.q_a_81(q_a_81),
	.q_a_24(q_a_24),
	.q_a_241(q_a_241),
	.q_a_2(q_a_2),
	.q_a_21(q_a_21),
	.av_readdata_pre_2(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.q_a_18(q_a_18),
	.q_a_181(q_a_181),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.q_a_10(q_a_10),
	.q_a_101(q_a_101),
	.q_a_26(q_a_26),
	.q_a_261(q_a_261),
	.q_a_5(q_a_5),
	.q_a_51(q_a_51),
	.av_readdata_pre_5(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.q_a_211(q_a_211),
	.q_a_212(q_a_212),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.q_a_13(q_a_13),
	.q_a_131(q_a_131),
	.q_a_29(q_a_29),
	.q_a_291(q_a_291),
	.q_a_7(q_a_7),
	.q_a_71(q_a_71),
	.av_readdata_pre_7(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.q_a_23(q_a_23),
	.q_a_231(q_a_231),
	.q_a_15(q_a_15),
	.q_a_151(q_a_151),
	.q_a_31(q_a_31),
	.q_a_311(q_a_311),
	.q_a_11(q_a_11),
	.q_a_111(q_a_111),
	.q_a_27(q_a_27),
	.q_a_271(q_a_271),
	.q_a_9(q_a_9),
	.q_a_91(q_a_91),
	.q_a_25(q_a_25),
	.q_a_251(q_a_251),
	.q_a_6(q_a_6),
	.q_a_61(q_a_61),
	.av_readdata_pre_6(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.q_a_22(q_a_22),
	.q_a_221(q_a_221),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_14(q_a_14),
	.q_a_141(q_a_141),
	.q_a_30(q_a_30),
	.q_a_301(q_a_301),
	.q_a_3(q_a_3),
	.q_a_32(q_a_32),
	.av_readdata_pre_3(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.q_a_19(q_a_19),
	.q_a_191(q_a_191),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_1(q_a_1),
	.q_a_17(q_a_17),
	.av_readdata_pre_1(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.q_a_171(q_a_171),
	.q_a_172(q_a_172),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.read_latency_shift_reg_0(\pio_led_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid(\rsp_demux_003|src0_valid~0_combout ),
	.src0_valid1(\rsp_demux_006|src0_valid~0_combout ),
	.src0_valid2(\rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\pio_key_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr11(WideOr1),
	.av_readdata_pre_30(\sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_41(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_201(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.src_data_20(src_data_20),
	.av_readdata_pre_12(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_121(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.src_data_28(src_data_28),
	.av_readdata_pre_01(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\pio_key_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\pio_led_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_161(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.src_data_16(src_data_16),
	.av_readdata_pre_8(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_81(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.src_data_24(src_data_24),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_181(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.src_data_18(src_data_18),
	.av_readdata_pre_10(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_101(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.src_data_10(src_data_10),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.src_data_26(src_data_26),
	.av_readdata_pre_51(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_211(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.src_data_21(src_data_21),
	.av_readdata_pre_13(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_131(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.src_data_13(src_data_13),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.src_data_29(src_data_29),
	.av_readdata_pre_71(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_231(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.src_data_23(src_data_23),
	.av_readdata_pre_15(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_151(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.src_data_15(src_data_15),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.src_data_31(src_data_31),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.src_data_11(src_data_11),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.src_data_27(src_data_27),
	.av_readdata_pre_9(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_91(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.src_data_25(src_data_25),
	.av_readdata_pre_61(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_221(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.src_data_22(src_data_22),
	.av_readdata_pre_14(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_141(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_301(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.src_data_30(src_data_30),
	.av_readdata_pre_32(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_191(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.src_data_19(src_data_19),
	.av_readdata_pre_110(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_17),
	.av_readdata_pre_171(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.src_data_17(src_data_171));

Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002_2 rsp_demux_006(
	.read_latency_shift_reg_0(\onchip_rom_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_rom_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_rom_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_006|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_006|src1_valid~0_combout ));

Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002_1 rsp_demux_003(
	.read_latency_shift_reg_0(\onchip_ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_003|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_003|src1_valid~0_combout ));

Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002 rsp_demux_002(
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_002|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ));

Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002_2 cmd_mux_006(
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_writedata_0(d_writedata_0),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_tag_field_2(d_address_tag_field_2),
	.d_address_offset_field_1(d_address_offset_field_1),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_02),
	.read_latency_shift_reg(\onchip_rom_s1_translator|read_latency_shift_reg~0_combout ),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.ic_fill_line_6(ic_fill_line_6),
	.src2_valid(src2_valid),
	.src6_valid(src6_valid),
	.saved_grant_1(saved_grant_11),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_0(ic_fill_line_0),
	.d_writedata_7(d_writedata_7),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_3(d_writedata_3),
	.d_writedata_1(d_writedata_1),
	.d_writedata_4(d_writedata_4),
	.src_payload(src_payload5),
	.src_data_38(src_data_382),
	.src_data_39(src_data_392),
	.src_data_40(src_data_402),
	.src_data_41(src_data_412),
	.src_data_42(src_data_422),
	.src_data_43(src_data_432),
	.src_data_44(src_data_442),
	.src_data_45(src_data_452),
	.src_data_46(src_data_462),
	.src_data_47(src_data_472),
	.src_data_48(src_data_481),
	.src_data_49(src_data_491),
	.src_data_32(src_data_322),
	.d_writedata_20(d_writedata_20),
	.d_byteenable_2(d_byteenable_2),
	.src_payload1(src_payload7),
	.src_data_34(src_data_341),
	.d_writedata_12(d_writedata_12),
	.d_byteenable_1(d_byteenable_1),
	.src_payload2(src_payload9),
	.src_data_33(src_data_332),
	.d_writedata_28(d_writedata_28),
	.d_byteenable_3(d_byteenable_3),
	.src_payload3(src_payload11),
	.src_data_35(src_data_351),
	.src_payload4(src_payload13),
	.d_writedata_16(d_writedata_16),
	.src_payload5(src_payload15),
	.d_writedata_8(d_writedata_8),
	.src_payload6(src_payload17),
	.d_writedata_24(d_writedata_24),
	.src_payload7(src_payload19),
	.d_writedata_2(d_writedata_2),
	.src_payload8(src_payload21),
	.d_writedata_18(d_writedata_18),
	.src_payload9(src_payload23),
	.d_writedata_10(d_writedata_10),
	.src_payload10(src_payload25),
	.d_writedata_26(d_writedata_26),
	.src_payload11(src_payload27),
	.d_writedata_5(d_writedata_5),
	.src_payload12(src_payload29),
	.d_writedata_21(d_writedata_21),
	.src_payload13(src_payload31),
	.d_writedata_13(d_writedata_13),
	.src_payload14(src_payload33),
	.d_writedata_29(d_writedata_29),
	.src_payload15(src_payload35),
	.src_payload16(src_payload37),
	.d_writedata_23(d_writedata_23),
	.src_payload17(src_payload39),
	.d_writedata_15(d_writedata_15),
	.src_payload18(src_payload41),
	.d_writedata_31(d_writedata_31),
	.src_payload19(src_payload43),
	.d_writedata_11(d_writedata_11),
	.src_payload20(src_payload45),
	.d_writedata_27(d_writedata_27),
	.src_payload21(src_payload47),
	.d_writedata_9(d_writedata_9),
	.src_payload22(src_payload49),
	.d_writedata_25(d_writedata_25),
	.src_payload23(src_payload51),
	.d_writedata_6(d_writedata_6),
	.src_payload24(src_payload53),
	.d_writedata_22(d_writedata_22),
	.src_payload25(src_payload55),
	.d_writedata_14(d_writedata_14),
	.src_payload26(src_payload57),
	.d_writedata_30(d_writedata_30),
	.src_payload27(src_payload59),
	.src_payload28(src_payload61),
	.d_writedata_19(d_writedata_19),
	.src_payload29(src_payload63),
	.src_payload30(src_payload66),
	.d_writedata_17(d_writedata_17),
	.src_payload31(src_payload68),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002_1 cmd_mux_003(
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_writedata_0(d_writedata_0),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_tag_field_3(d_address_tag_field_3),
	.d_address_tag_field_2(d_address_tag_field_2),
	.d_address_offset_field_1(d_address_offset_field_1),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.ic_fill_line_6(ic_fill_line_6),
	.src1_valid(src1_valid),
	.src3_valid(src3_valid),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_1(saved_grant_1),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_0(ic_fill_line_0),
	.d_writedata_7(d_writedata_7),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_3(d_writedata_3),
	.d_writedata_1(d_writedata_1),
	.d_writedata_4(d_writedata_4),
	.src_payload(src_payload4),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_46(src_data_461),
	.src_data_47(src_data_471),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.src_data_32(src_data_321),
	.d_writedata_20(d_writedata_20),
	.src_payload1(src_payload6),
	.d_byteenable_2(d_byteenable_2),
	.src_data_34(src_data_34),
	.d_writedata_12(d_writedata_12),
	.src_payload2(src_payload8),
	.d_byteenable_1(d_byteenable_1),
	.src_data_33(src_data_331),
	.d_writedata_28(d_writedata_28),
	.src_payload3(src_payload10),
	.d_byteenable_3(d_byteenable_3),
	.src_data_35(src_data_35),
	.src_payload4(src_payload12),
	.d_writedata_16(d_writedata_16),
	.src_payload5(src_payload14),
	.d_writedata_8(d_writedata_8),
	.src_payload6(src_payload16),
	.d_writedata_24(d_writedata_24),
	.src_payload7(src_payload18),
	.d_writedata_2(d_writedata_2),
	.src_payload8(src_payload20),
	.d_writedata_18(d_writedata_18),
	.src_payload9(src_payload22),
	.d_writedata_10(d_writedata_10),
	.src_payload10(src_payload24),
	.d_writedata_26(d_writedata_26),
	.src_payload11(src_payload26),
	.d_writedata_5(d_writedata_5),
	.src_payload12(src_payload28),
	.d_writedata_21(d_writedata_21),
	.src_payload13(src_payload30),
	.d_writedata_13(d_writedata_13),
	.src_payload14(src_payload32),
	.d_writedata_29(d_writedata_29),
	.src_payload15(src_payload34),
	.src_payload16(src_payload36),
	.d_writedata_23(d_writedata_23),
	.src_payload17(src_payload38),
	.d_writedata_15(d_writedata_15),
	.src_payload18(src_payload40),
	.d_writedata_31(d_writedata_31),
	.src_payload19(src_payload42),
	.d_writedata_11(d_writedata_11),
	.src_payload20(src_payload44),
	.d_writedata_27(d_writedata_27),
	.src_payload21(src_payload46),
	.d_writedata_9(d_writedata_9),
	.src_payload22(src_payload48),
	.d_writedata_25(d_writedata_25),
	.src_payload23(src_payload50),
	.d_writedata_6(d_writedata_6),
	.src_payload24(src_payload52),
	.d_writedata_22(d_writedata_22),
	.src_payload25(src_payload54),
	.d_writedata_14(d_writedata_14),
	.src_payload26(src_payload56),
	.d_writedata_30(d_writedata_30),
	.src_payload27(src_payload58),
	.src_payload28(src_payload60),
	.d_writedata_19(d_writedata_19),
	.src_payload29(src_payload62),
	.src_payload30(src_payload65),
	.d_writedata_17(d_writedata_17),
	.src_payload31(src_payload67),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002 cmd_mux_002(
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_writedata_0(d_writedata_0),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_offset_field_1(d_address_offset_field_1),
	.r_sync_rst(r_sync_rst),
	.Equal2(\router|Equal2~0_combout ),
	.saved_grant_0(saved_grant_01),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.Equal21(\router_001|Equal2~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~1_combout ),
	.src0_valid1(\cmd_demux_001|src0_valid~2_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux|src2_valid~1_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.WideOr11(WideOr11),
	.hbreak_enabled(hbreak_enabled),
	.ic_fill_line_5(ic_fill_line_5),
	.src_data_46(src_data_46),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_0(ic_fill_line_0),
	.d_writedata_7(d_writedata_7),
	.src_payload(src_payload),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.src_data_38(src_data_38),
	.src_data_41(src_data_41),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.src_data_40(src_data_40),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.src_data_39(src_data_39),
	.src_data_45(src_data_45),
	.src_data_44(src_data_44),
	.src_data_43(src_data_43),
	.src_data_42(src_data_42),
	.src_payload1(src_payload1),
	.d_byteenable_0(d_byteenable_0),
	.src_data_32(src_data_32),
	.d_writedata_3(d_writedata_3),
	.src_payload2(src_payload2),
	.d_writedata_1(d_writedata_1),
	.src_payload3(src_payload3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_20(d_writedata_20),
	.d_byteenable_2(d_byteenable_2),
	.d_writedata_12(d_writedata_12),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_28(d_writedata_28),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_16(d_writedata_16),
	.d_writedata_8(d_writedata_8),
	.d_writedata_24(d_writedata_24),
	.d_writedata_2(d_writedata_2),
	.d_writedata_18(d_writedata_18),
	.d_writedata_10(d_writedata_10),
	.d_writedata_26(d_writedata_26),
	.d_writedata_5(d_writedata_5),
	.d_writedata_21(d_writedata_21),
	.d_writedata_13(d_writedata_13),
	.d_writedata_29(d_writedata_29),
	.d_writedata_23(d_writedata_23),
	.d_writedata_15(d_writedata_15),
	.d_writedata_31(d_writedata_31),
	.d_writedata_11(d_writedata_11),
	.d_writedata_27(d_writedata_27),
	.d_writedata_9(d_writedata_9),
	.d_writedata_25(d_writedata_25),
	.d_writedata_6(d_writedata_6),
	.d_writedata_22(d_writedata_22),
	.d_writedata_14(d_writedata_14),
	.d_writedata_30(d_writedata_30),
	.d_writedata_19(d_writedata_19),
	.src_payload4(src_payload64),
	.d_writedata_17(d_writedata_17),
	.src_payload5(src_payload69),
	.src_data_34(src_data_342),
	.src_payload6(src_payload70),
	.src_payload7(src_payload71),
	.src_payload8(src_payload72),
	.src_data_35(src_data_352),
	.src_payload9(src_payload73),
	.src_payload10(src_payload74),
	.src_payload11(src_payload75),
	.src_payload12(src_payload76),
	.src_payload13(src_payload77),
	.src_payload14(src_payload78),
	.src_payload15(src_payload79),
	.src_payload16(src_payload80),
	.src_data_33(src_data_333),
	.src_payload17(src_payload81),
	.src_payload18(src_payload82),
	.src_payload19(src_payload83),
	.src_payload20(src_payload84),
	.src_payload21(src_payload85),
	.src_payload22(src_payload86),
	.src_payload23(src_payload87),
	.src_payload24(src_payload88),
	.src_payload25(src_payload89),
	.src_payload26(src_payload90),
	.src_payload27(src_payload91),
	.src_payload28(src_payload92),
	.src_payload29(src_payload93),
	.src_payload30(src_payload94),
	.src_payload31(src_payload95),
	.src_payload32(src_payload96),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.WideOr0(WideOr0),
	.rst1(rst1),
	.mem_used_1(mem_used_11),
	.waitrequest(waitrequest),
	.mem_used_11(mem_used_13),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.has_pending_responses(has_pending_responses),
	.i_read(i_read),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.last_channel_1(\nios2_qsys_0_instruction_master_limiter|last_channel[1]~q ),
	.src_channel_1(\router_001|src_channel[1]~0_combout ),
	.src1_valid(src1_valid),
	.saved_grant_1(saved_grant_1),
	.Equal2(\router_001|Equal2~0_combout ),
	.last_channel_0(\nios2_qsys_0_instruction_master_limiter|last_channel[0]~q ),
	.src0_valid1(\cmd_demux_001|src0_valid~1_combout ),
	.src0_valid2(\cmd_demux_001|src0_valid~2_combout ),
	.saved_grant_11(\cmd_mux_002|saved_grant[1]~q ),
	.Equal1(\router_001|Equal1~0_combout ),
	.last_channel_2(\nios2_qsys_0_instruction_master_limiter|last_channel[2]~q ),
	.src2_valid(src2_valid),
	.mem(\onchip_rom_s1_agent_rsp_fifo|mem~3_combout ));

Qsys_system_Qsys_system_mm_interconnect_0_cmd_demux cmd_demux(
	.rst1(rst1),
	.d_write(d_write),
	.mem_used_1(\pio_led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.d_read(d_read),
	.has_pending_responses(\nios2_qsys_0_data_master_limiter|has_pending_responses~q ),
	.suppress_change_dest_id(suppress_change_dest_id),
	.av_waitrequest(av_waitrequest),
	.always1(\router|always1~0_combout ),
	.Equal4(Equal4),
	.Equal2(\router|Equal2~0_combout ),
	.src_data_77(\router|src_data[77]~0_combout ),
	.Equal1(\router|Equal1~0_combout ),
	.mem_used_11(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_11(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\sysid_qsys_0_control_slave_translator|wait_latency_counter[0]~q ),
	.src_channel_3(\router|src_channel[3]~0_combout ),
	.Equal3(\router|Equal3~2_combout ),
	.mem_used_12(mem_used_1),
	.wait_latency_counter_12(wait_latency_counter_11),
	.wait_latency_counter_02(wait_latency_counter_01),
	.saved_grant_0(saved_grant_0),
	.mem_used_13(mem_used_11),
	.av_waitrequest1(av_waitrequest1),
	.mem_used_14(mem_used_12),
	.saved_grant_01(saved_grant_01),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.saved_grant_02(saved_grant_02),
	.read_latency_shift_reg(\onchip_rom_s1_translator|read_latency_shift_reg~0_combout ),
	.WideOr01(WideOr01),
	.cp_valid(cp_valid),
	.last_channel_3(\nios2_qsys_0_data_master_limiter|last_channel[3]~q ),
	.src3_valid(src3_valid),
	.last_channel_2(\nios2_qsys_0_data_master_limiter|last_channel[2]~q ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux|src2_valid~1_combout ),
	.last_channel_6(\nios2_qsys_0_data_master_limiter|last_channel[6]~q ),
	.src6_valid(src6_valid));

Qsys_system_altera_merlin_traffic_limiter_1 nios2_qsys_0_instruction_master_limiter(
	.WideOr0(WideOr0),
	.reset(r_sync_rst),
	.mem_61_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_01(\onchip_rom_s1_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_02(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ),
	.has_pending_responses1(has_pending_responses),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.last_channel_1(\nios2_qsys_0_instruction_master_limiter|last_channel[1]~q ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router_001|src_channel[1]~0_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_sink_channel({gnd,gnd,gnd,gnd,\router_001|Equal1~0_combout ,gnd,\router_001|Equal2~0_combout }),
	.last_channel_0(\nios2_qsys_0_instruction_master_limiter|last_channel[0]~q ),
	.last_channel_2(\nios2_qsys_0_instruction_master_limiter|last_channel[2]~q ),
	.save_dest_id(save_dest_id),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.src1_valid2(\rsp_demux_006|src1_valid~0_combout ),
	.suppress_change_dest_id(suppress_change_dest_id2),
	.clk(clk_clk));

Qsys_system_altera_merlin_traffic_limiter nios2_qsys_0_data_master_limiter(
	.d_write(d_write),
	.reset(r_sync_rst),
	.has_pending_responses1(\nios2_qsys_0_data_master_limiter|has_pending_responses~q ),
	.suppress_change_dest_id(suppress_change_dest_id),
	.cmd_sink_channel({\router|Equal1~0_combout ,Equal4,\router|Equal3~2_combout ,\router|src_channel[3]~0_combout ,\router|Equal2~0_combout ,\router|always1~0_combout ,av_waitrequest}),
	.src_data_77(\router|src_data[77]~0_combout ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router|src_data[79]~2_combout ,\router|src_data[78]~3_combout ,\router|src_data[77]~1_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.suppress_change_dest_id1(suppress_change_dest_id1),
	.WideOr0(WideOr01),
	.read_latency_shift_reg_0(\pio_led_s1_translator|read_latency_shift_reg[0]~q ),
	.last_channel_4(\nios2_qsys_0_data_master_limiter|last_channel[4]~q ),
	.cp_valid(cp_valid),
	.src0_valid(\rsp_demux_003|src0_valid~0_combout ),
	.src0_valid1(\rsp_demux_006|src0_valid~0_combout ),
	.mem_61_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_01(\onchip_rom_s1_agent_rsp_fifo|mem[0][61]~q ),
	.src0_valid2(\rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\pio_key_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(WideOr1),
	.mem_61_02(\pio_led_s1_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_03(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_04(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_05(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_06(\pio_key_s1_agent_rsp_fifo|mem[0][61]~q ),
	.last_channel_1(\nios2_qsys_0_data_master_limiter|last_channel[1]~q ),
	.last_channel_5(\nios2_qsys_0_data_master_limiter|last_channel[5]~q ),
	.last_channel_3(\nios2_qsys_0_data_master_limiter|last_channel[3]~q ),
	.last_channel_0(last_channel_0),
	.last_channel_2(\nios2_qsys_0_data_master_limiter|last_channel[2]~q ),
	.last_channel_6(\nios2_qsys_0_data_master_limiter|last_channel[6]~q ),
	.clk(clk_clk));

Qsys_system_Qsys_system_mm_interconnect_0_router_001 router_001(
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.ic_fill_line_6(ic_fill_line_6),
	.src_channel_1(\router_001|src_channel[1]~0_combout ),
	.Equal2(\router_001|Equal2~0_combout ),
	.Equal1(\router_001|Equal1~0_combout ));

Qsys_system_Qsys_system_mm_interconnect_0_router router(
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.Equal3(Equal3),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_tag_field_5(d_address_tag_field_5),
	.d_address_tag_field_4(d_address_tag_field_4),
	.d_address_tag_field_3(d_address_tag_field_3),
	.d_address_tag_field_2(d_address_tag_field_2),
	.Equal31(Equal31),
	.d_address_offset_field_1(d_address_offset_field_1),
	.d_read(d_read),
	.av_waitrequest(av_waitrequest),
	.always1(\router|always1~0_combout ),
	.Equal4(Equal4),
	.Equal2(\router|Equal2~0_combout ),
	.src_data_77(\router|src_data[77]~0_combout ),
	.Equal1(\router|Equal1~0_combout ),
	.src_data_771(\router|src_data[77]~1_combout ),
	.src_data_79(\router|src_data[79]~2_combout ),
	.src_channel_3(\router|src_channel[3]~0_combout ),
	.Equal32(\router|Equal3~2_combout ),
	.src_data_78(\router|src_data[78]~3_combout ));

Qsys_system_altera_avalon_sc_fifo_3 onchip_rom_s1_agent_rsp_fifo(
	.rst1(rst1),
	.reset(r_sync_rst),
	.d_read(d_read),
	.saved_grant_0(saved_grant_02),
	.mem_used_1(mem_used_14),
	.read_latency_shift_reg_0(\onchip_rom_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_rom_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_rom_s1_agent_rsp_fifo|mem[0][56]~q ),
	.mem_61_0(\onchip_rom_s1_agent_rsp_fifo|mem[0][61]~q ),
	.i_read(i_read),
	.saved_grant_1(saved_grant_11),
	.rf_source_valid(\onchip_rom_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg(\onchip_rom_s1_translator|read_latency_shift_reg~1_combout ),
	.mem(\onchip_rom_s1_agent_rsp_fifo|mem~3_combout ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_agent_3 onchip_rom_s1_agent(
	.d_read(d_read),
	.saved_grant_0(saved_grant_02),
	.i_read(i_read),
	.src2_valid(src2_valid),
	.src6_valid(src6_valid),
	.saved_grant_1(saved_grant_11),
	.rf_source_valid(\onchip_rom_s1_agent|rf_source_valid~0_combout ));

Qsys_system_altera_avalon_sc_fifo_4 pio_key_s1_agent_rsp_fifo(
	.rst1(rst1),
	.reset(r_sync_rst),
	.Equal4(Equal4),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg_0(\pio_key_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_61_0(\pio_key_s1_agent_rsp_fifo|mem[0][61]~q ),
	.read_latency_shift_reg(\pio_key_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg1(\pio_key_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

Qsys_system_altera_avalon_sc_fifo_5 pio_led_s1_agent_rsp_fifo(
	.mem_used_1(\pio_led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\pio_led_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\pio_led_s1_translator|read_latency_shift_reg~1_combout ),
	.mem_61_0(\pio_led_s1_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

Qsys_system_altera_merlin_slave_agent_5 pio_led_s1_agent(
	.always2(always2),
	.mem_used_1(\pio_led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.d_address_line_field_0(d_address_line_field_0),
	.Equal3(Equal3),
	.Equal31(Equal31),
	.m0_write(m0_write));

Qsys_system_altera_avalon_sc_fifo_2 onchip_ram_s1_agent_rsp_fifo(
	.rst1(rst1),
	.reset(r_sync_rst),
	.d_read(d_read),
	.saved_grant_0(saved_grant_0),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\onchip_ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][56]~q ),
	.mem_61_0(\onchip_ram_s1_agent_rsp_fifo|mem[0][61]~q ),
	.i_read(i_read),
	.saved_grant_1(saved_grant_1),
	.rf_source_valid(\onchip_ram_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

endmodule

module Qsys_system_altera_avalon_sc_fifo (
	reset,
	av_waitrequest,
	av_waitrequest1,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_61_0,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_61_0;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][94]~q ;
wire \mem~0_combout ;
wire \mem[0][61]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem[0][61]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!av_waitrequest),
	.datab(!av_waitrequest1),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFFFFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][61]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(!mem_61_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][61]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][61]~1 .extended_lut = "off";
defparam \mem[0][61]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \mem[0][61]~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_1 (
	reset,
	d_read,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	mem_61_0,
	i_read,
	saved_grant_1,
	rf_source_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_read;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	mem_61_0;
input 	i_read;
input 	saved_grant_1;
input 	rf_source_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem[1][94]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hBF8FFFFFBF8FFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBFBFFF3FBFBFFF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][56]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][94]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_2 (
	rst1,
	reset,
	d_read,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	mem_61_0,
	i_read,
	saved_grant_1,
	rf_source_valid,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	d_read;
input 	saved_grant_0;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	mem_61_0;
input 	i_read;
input 	saved_grant_1;
input 	rf_source_valid;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem[1][94]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][56]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][94]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_3 (
	rst1,
	reset,
	d_read,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	mem_61_0,
	i_read,
	saved_grant_1,
	rf_source_valid,
	read_latency_shift_reg,
	mem,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	d_read;
input 	saved_grant_0;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	mem_61_0;
input 	i_read;
input 	saved_grant_1;
input 	rf_source_valid;
input 	read_latency_shift_reg;
output 	mem;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem[1][94]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~3 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][56]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][94]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_4 (
	rst1,
	reset,
	Equal4,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_61_0,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	Equal4;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_61_0;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][94]~q ;
wire \mem~0_combout ;
wire \mem[0][61]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem[0][61]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!rst1),
	.datab(!Equal4),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFFFFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][61]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(!mem_61_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][61]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][61]~1 .extended_lut = "off";
defparam \mem[0][61]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \mem[0][61]~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_5 (
	mem_used_1,
	reset,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	mem_61_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	mem_used_1;
input 	reset;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;
output 	mem_61_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][94]~q ;
wire \mem~0_combout ;
wire \mem[0][61]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem[0][61]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][61]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(!mem_61_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][61]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][61]~1 .extended_lut = "off";
defparam \mem[0][61]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \mem[0][61]~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_avalon_sc_fifo_6 (
	rst1,
	reset,
	suppress_change_dest_id,
	always1,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_61_0,
	av_waitrequest_generated,
	last_channel_1,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	suppress_change_dest_id;
input 	always1;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_61_0;
input 	av_waitrequest_generated;
input 	last_channel_1;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][94]~q ;
wire \mem~0_combout ;
wire \mem[0][61]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem[0][61]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~3 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~3 .extended_lut = "off";
defparam \mem_used[0]~3 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~3 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!suppress_change_dest_id),
	.datab(!last_channel_1),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!rst1),
	.datab(!always1),
	.datac(!av_waitrequest_generated),
	.datad(!\mem_used[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!\mem_used[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \mem_used[1]~2 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][61]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(!mem_61_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][61]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][61]~1 .extended_lut = "off";
defparam \mem[0][61]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \mem[0][61]~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_master_agent (
	rst1,
	d_write,
	d_read,
	suppress_change_dest_id,
	WideOr0,
	av_waitrequest1,
	cp_valid)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	d_write;
input 	d_read;
input 	suppress_change_dest_id;
input 	WideOr0;
output 	av_waitrequest1;
output 	cp_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb av_waitrequest(
	.dataa(!rst1),
	.datab(!suppress_change_dest_id),
	.datac(!WideOr0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam av_waitrequest.extended_lut = "off";
defparam av_waitrequest.lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam av_waitrequest.shared_arith = "off";

cyclonev_lcell_comb \cp_valid~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!d_read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_valid~0 .extended_lut = "off";
defparam \cp_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \cp_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_agent_1 (
	d_read,
	saved_grant_0,
	i_read,
	saved_grant_1,
	WideOr1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	saved_grant_0;
input 	i_read;
input 	saved_grant_1;
input 	WideOr1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!saved_grant_1),
	.datae(!WideOr1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_agent_2 (
	d_read,
	saved_grant_0,
	i_read,
	src1_valid,
	src3_valid,
	saved_grant_1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	saved_grant_0;
input 	i_read;
input 	src1_valid;
input 	src3_valid;
input 	saved_grant_1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!src1_valid),
	.datae(!src3_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_agent_3 (
	d_read,
	saved_grant_0,
	i_read,
	src2_valid,
	src6_valid,
	saved_grant_1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	saved_grant_0;
input 	i_read;
input 	src2_valid;
input 	src6_valid;
input 	saved_grant_1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!src2_valid),
	.datae(!src6_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_agent_5 (
	always2,
	mem_used_1,
	d_address_line_field_0,
	Equal3,
	Equal31,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	always2;
input 	mem_used_1;
input 	d_address_line_field_0;
input 	Equal3;
input 	Equal31;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!always2),
	.datab(!mem_used_1),
	.datac(!d_address_line_field_0),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_agent_6 (
	rst1,
	always1,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	always1;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(!always1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator (
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_1,
	av_readdata_pre_17,
	q_b_4,
	av_readdata,
	q_b_0,
	q_b_2,
	q_b_5,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_1,
	rst1,
	reset,
	d_read,
	suppress_change_dest_id,
	av_waitrequest,
	av_waitrequest1,
	mem_used_1,
	read_latency_shift_reg_0,
	last_channel_0,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	b_full,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	av_readdata_pre_12,
	av_readdata_pre_8,
	av_readdata_pre_10,
	av_readdata_pre_13,
	av_readdata_pre_15,
	av_readdata_pre_9,
	av_readdata_pre_14,
	b_full1,
	read_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_4;
output 	av_readdata_pre_20;
output 	av_readdata_pre_0;
output 	av_readdata_pre_16;
output 	av_readdata_pre_2;
output 	av_readdata_pre_18;
output 	av_readdata_pre_5;
output 	av_readdata_pre_21;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_22;
output 	av_readdata_pre_3;
output 	av_readdata_pre_19;
output 	av_readdata_pre_1;
output 	av_readdata_pre_17;
input 	q_b_4;
input 	[31:0] av_readdata;
input 	q_b_0;
input 	q_b_2;
input 	q_b_5;
input 	q_b_7;
input 	q_b_6;
input 	q_b_3;
input 	q_b_1;
input 	rst1;
input 	reset;
input 	d_read;
input 	suppress_change_dest_id;
input 	av_waitrequest;
input 	av_waitrequest1;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
input 	last_channel_0;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg1;
input 	b_full;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
output 	av_readdata_pre_12;
output 	av_readdata_pre_8;
output 	av_readdata_pre_10;
output 	av_readdata_pre_13;
output 	av_readdata_pre_15;
output 	av_readdata_pre_9;
output 	av_readdata_pre_14;
input 	b_full1;
input 	read_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[13]~0_combout ;


dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(q_b_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_7),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_6),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(q_b_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(q_b_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!d_read),
	.datac(!suppress_change_dest_id),
	.datad(!last_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!av_waitrequest),
	.datab(!av_waitrequest1),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

cyclonev_lcell_comb \av_readdata_pre[13]~0 (
	.dataa(!b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_readdata_pre[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata_pre[13]~0 .extended_lut = "off";
defparam \av_readdata_pre[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \av_readdata_pre[13]~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_1 (
	av_readdata,
	rst1,
	reset,
	sink_ready,
	read_latency_shift_reg_0,
	rf_source_valid,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_12,
	av_readdata_pre_28,
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_8,
	av_readdata_pre_24,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_10,
	av_readdata_pre_26,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_13,
	av_readdata_pre_29,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_11,
	av_readdata_pre_27,
	av_readdata_pre_9,
	av_readdata_pre_25,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_14,
	av_readdata_pre_30,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_1,
	av_readdata_pre_17,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	rst1;
input 	reset;
input 	sink_ready;
output 	read_latency_shift_reg_0;
input 	rf_source_valid;
output 	av_readdata_pre_4;
output 	av_readdata_pre_20;
output 	av_readdata_pre_12;
output 	av_readdata_pre_28;
output 	av_readdata_pre_0;
output 	av_readdata_pre_16;
output 	av_readdata_pre_8;
output 	av_readdata_pre_24;
output 	av_readdata_pre_2;
output 	av_readdata_pre_18;
output 	av_readdata_pre_10;
output 	av_readdata_pre_26;
output 	av_readdata_pre_5;
output 	av_readdata_pre_21;
output 	av_readdata_pre_13;
output 	av_readdata_pre_29;
output 	av_readdata_pre_7;
output 	av_readdata_pre_23;
output 	av_readdata_pre_15;
output 	av_readdata_pre_31;
output 	av_readdata_pre_11;
output 	av_readdata_pre_27;
output 	av_readdata_pre_9;
output 	av_readdata_pre_25;
output 	av_readdata_pre_6;
output 	av_readdata_pre_22;
output 	av_readdata_pre_14;
output 	av_readdata_pre_30;
output 	av_readdata_pre_3;
output 	av_readdata_pre_19;
output 	av_readdata_pre_1;
output 	av_readdata_pre_17;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!sink_ready),
	.datac(!rf_source_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_2 (
	rst1,
	reset,
	mem_used_1,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	rf_source_valid,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	rf_source_valid;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!read_latency_shift_reg),
	.datab(!rf_source_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_3 (
	rst1,
	reset,
	mem_used_1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	rf_source_valid,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	reset;
input 	mem_used_1;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	rf_source_valid;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!read_latency_shift_reg),
	.datab(!rf_source_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_4 (
	rst1,
	d_write,
	reset,
	d_read,
	av_begintransfer,
	suppress_change_dest_id,
	Equal4,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	last_channel_5,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	av_readdata_pre_0,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	d_write;
input 	reset;
input 	d_read;
input 	av_begintransfer;
input 	suppress_change_dest_id;
input 	Equal4;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	last_channel_5;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg1;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_waitrequest_generated~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!d_read),
	.datab(!\av_waitrequest_generated~0_combout ),
	.datac(!suppress_change_dest_id),
	.datad(!last_channel_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!rst1),
	.datab(!Equal4),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!Equal4),
	.datad(!mem_used_1),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest_generated~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hFFFF9669FFFF6996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!av_begintransfer),
	.datab(!suppress_change_dest_id),
	.datac(!last_channel_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(!rst1),
	.datab(!Equal4),
	.datac(!mem_used_1),
	.datad(!\av_waitrequest_generated~0_combout ),
	.datae(!\wait_latency_counter[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~1 .extended_lut = "off";
defparam \wait_latency_counter[1]~1 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \wait_latency_counter[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~3 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~3 .extended_lut = "off";
defparam \wait_latency_counter~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \wait_latency_counter~3 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_5 (
	rst1,
	always2,
	mem_used_1,
	m0_write,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset,
	d_read,
	suppress_change_dest_id,
	Equal3,
	read_latency_shift_reg_0,
	last_channel_4,
	read_latency_shift_reg,
	cp_valid,
	av_readdata_pre_0,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	always2;
input 	mem_used_1;
input 	m0_write;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	reset;
input 	d_read;
input 	suppress_change_dest_id;
input 	Equal3;
output 	read_latency_shift_reg_0;
input 	last_channel_4;
output 	read_latency_shift_reg;
input 	cp_valid;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \read_latency_shift_reg~2_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!d_read),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(!suppress_change_dest_id),
	.datad(!last_channel_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!suppress_change_dest_id),
	.datab(!last_channel_4),
	.datac(!cp_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!always2),
	.datad(!mem_used_1),
	.datae(!Equal3),
	.dataf(!\wait_latency_counter[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~1 .extended_lut = "off";
defparam \wait_latency_counter[0]~1 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \wait_latency_counter[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~3 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~3 .extended_lut = "off";
defparam \wait_latency_counter~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \wait_latency_counter~3 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~2 .extended_lut = "off";
defparam \read_latency_shift_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \read_latency_shift_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!rst1),
	.datad(!Equal3),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hBFFFEFFFBFFFEFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_slave_translator_6 (
	av_readdata,
	rst1,
	d_write,
	reset,
	d_read,
	av_begintransfer,
	suppress_change_dest_id,
	always1,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_waitrequest_generated,
	last_channel_1,
	m0_write,
	read_latency_shift_reg,
	av_readdata_pre_30,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	rst1;
input 	d_write;
input 	reset;
input 	d_read;
output 	av_begintransfer;
input 	suppress_change_dest_id;
input 	always1;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_waitrequest_generated;
input 	last_channel_1;
input 	m0_write;
output 	read_latency_shift_reg;
output 	av_readdata_pre_30;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;


cyclonev_lcell_comb \av_begintransfer~0 (
	.dataa(!d_write),
	.datab(!d_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_begintransfer),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_begintransfer~0 .extended_lut = "off";
defparam \av_begintransfer~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \av_begintransfer~0 .shared_arith = "off";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!mem_used_1),
	.datad(!always1),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hFFFF9669FFFF6996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!m0_write),
	.datab(!av_waitrequest_generated),
	.datac(!suppress_change_dest_id),
	.datad(!last_channel_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!m0_write),
	.datab(!av_waitrequest_generated),
	.datac(!suppress_change_dest_id),
	.datad(!last_channel_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \wait_latency_counter~2 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_traffic_limiter (
	d_write,
	reset,
	has_pending_responses1,
	suppress_change_dest_id,
	cmd_sink_channel,
	src_data_77,
	cmd_sink_data,
	suppress_change_dest_id1,
	WideOr0,
	read_latency_shift_reg_0,
	last_channel_4,
	cp_valid,
	src0_valid,
	src0_valid1,
	mem_61_0,
	mem_61_01,
	src0_valid2,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	WideOr1,
	mem_61_02,
	mem_61_03,
	mem_61_04,
	mem_61_05,
	mem_61_06,
	last_channel_1,
	last_channel_5,
	last_channel_3,
	last_channel_0,
	last_channel_2,
	last_channel_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	reset;
output 	has_pending_responses1;
output 	suppress_change_dest_id;
input 	[6:0] cmd_sink_channel;
input 	src_data_77;
input 	[92:0] cmd_sink_data;
output 	suppress_change_dest_id1;
input 	WideOr0;
input 	read_latency_shift_reg_0;
output 	last_channel_4;
input 	cp_valid;
input 	src0_valid;
input 	src0_valid1;
input 	mem_61_0;
input 	mem_61_01;
input 	src0_valid2;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	WideOr1;
input 	mem_61_02;
input 	mem_61_03;
input 	mem_61_04;
input 	mem_61_05;
input 	mem_61_06;
output 	last_channel_1;
output 	last_channel_5;
output 	last_channel_3;
output 	last_channel_0;
output 	last_channel_2;
output 	last_channel_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_dest_id[0]~q ;
wire \last_dest_id[1]~q ;
wire \Equal0~0_combout ;
wire \last_dest_id[2]~q ;
wire \Equal0~1_combout ;
wire \save_dest_id~0_combout ;
wire \save_dest_id~1_combout ;
wire \nonposted_cmd_accepted~combout ;
wire \response_sink_accepted~0_combout ;
wire \response_sink_accepted~1_combout ;
wire \response_sink_accepted~2_combout ;
wire \response_sink_accepted~3_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!d_write),
	.datab(!has_pending_responses1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \suppress_change_dest_id~1 (
	.dataa(!suppress_change_dest_id),
	.datab(!\last_dest_id[0]~q ),
	.datac(!cmd_sink_data[77]),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id1),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~1 .extended_lut = "off";
defparam \suppress_change_dest_id~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \suppress_change_dest_id~1 .shared_arith = "off";

dffeas \last_channel[4] (
	.clk(clk),
	.d(cmd_sink_channel[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_4),
	.prn(vcc));
defparam \last_channel[4] .is_wysiwyg = "true";
defparam \last_channel[4] .power_up = "low";

dffeas \last_channel[1] (
	.clk(clk),
	.d(cmd_sink_channel[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas \last_channel[5] (
	.clk(clk),
	.d(cmd_sink_channel[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_5),
	.prn(vcc));
defparam \last_channel[5] .is_wysiwyg = "true";
defparam \last_channel[5] .power_up = "low";

dffeas \last_channel[3] (
	.clk(clk),
	.d(cmd_sink_channel[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_3),
	.prn(vcc));
defparam \last_channel[3] .is_wysiwyg = "true";
defparam \last_channel[3] .power_up = "low";

dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

dffeas \last_channel[6] (
	.clk(clk),
	.d(cmd_sink_channel[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(last_channel_6),
	.prn(vcc));
defparam \last_channel[6] .is_wysiwyg = "true";
defparam \last_channel[6] .power_up = "low";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[77]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(cmd_sink_data[78]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(\last_dest_id[1]~q ),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!cmd_sink_channel[0]),
	.datab(!cmd_sink_channel[1]),
	.datac(!cmd_sink_channel[5]),
	.datad(!src_data_77),
	.datae(!\last_dest_id[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h9669699696696996;
defparam \Equal0~0 .shared_arith = "off";

dffeas \last_dest_id[2] (
	.clk(clk),
	.d(cmd_sink_data[79]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~1_combout ),
	.q(\last_dest_id[2]~q ),
	.prn(vcc));
defparam \last_dest_id[2] .is_wysiwyg = "true";
defparam \last_dest_id[2] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\last_dest_id[2]~q ),
	.datab(!cmd_sink_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h6666666666666666;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~1 (
	.dataa(!suppress_change_dest_id),
	.datab(!\last_dest_id[0]~q ),
	.datac(!cmd_sink_data[77]),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(!\save_dest_id~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~1 .extended_lut = "off";
defparam \save_dest_id~1 .lut_mask = 64'hFFFFFFBEFFFFFFFF;
defparam \save_dest_id~1 .shared_arith = "off";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!WideOr0),
	.datab(!\save_dest_id~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nonposted_cmd_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_02),
	.datac(!mem_61_03),
	.datad(!mem_61_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~1 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!src0_valid2),
	.datac(!mem_61_05),
	.datad(!mem_61_06),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~1 .extended_lut = "off";
defparam \response_sink_accepted~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \response_sink_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_61_02),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(!\response_sink_accepted~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~2 .extended_lut = "off";
defparam \response_sink_accepted~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \response_sink_accepted~2 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~3 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_61_0),
	.datad(!mem_61_01),
	.datae(!WideOr1),
	.dataf(!\response_sink_accepted~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~3 .extended_lut = "off";
defparam \response_sink_accepted~3 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \response_sink_accepted~3 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!\nonposted_cmd_accepted~combout ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h9696969696969696;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!\nonposted_cmd_accepted~combout ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \has_pending_responses~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_traffic_limiter_1 (
	WideOr0,
	reset,
	mem_61_0,
	mem_61_01,
	mem_61_02,
	has_pending_responses1,
	src0_valid,
	last_channel_1,
	cmd_sink_data,
	cmd_sink_channel,
	last_channel_0,
	last_channel_2,
	save_dest_id,
	nonposted_cmd_accepted1,
	src1_valid,
	src1_valid1,
	src1_valid2,
	suppress_change_dest_id,
	clk)/* synthesis synthesis_greybox=1 */;
input 	WideOr0;
input 	reset;
input 	mem_61_0;
input 	mem_61_01;
input 	mem_61_02;
output 	has_pending_responses1;
input 	src0_valid;
output 	last_channel_1;
input 	[92:0] cmd_sink_data;
input 	[6:0] cmd_sink_channel;
output 	last_channel_0;
output 	last_channel_2;
output 	save_dest_id;
output 	nonposted_cmd_accepted1;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
output 	suppress_change_dest_id;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \response_sink_accepted~0_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;
wire \last_channel[1]~0_combout ;
wire \last_dest_id[0]~q ;
wire \last_dest_id[1]~0_combout ;
wire \last_dest_id[1]~q ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_channel[1] (
	.clk(clk),
	.d(\last_channel[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!has_pending_responses1),
	.datab(!src0_valid),
	.datac(!cmd_sink_channel[0]),
	.datad(!cmd_sink_channel[2]),
	.datae(!\last_dest_id[0]~q ),
	.dataf(!\last_dest_id[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(save_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hBFFBFBBFFBBFBFFB;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!save_dest_id),
	.datab(!WideOr0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'h7777777777777777;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!cmd_sink_channel[0]),
	.datab(!cmd_sink_channel[2]),
	.datac(!\last_dest_id[0]~q ),
	.datad(!\last_dest_id[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'h6996699669966996;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!mem_61_02),
	.datab(!mem_61_0),
	.datac(!mem_61_01),
	.datad(!src1_valid),
	.datae(!src1_valid1),
	.dataf(!src1_valid2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!nonposted_cmd_accepted1),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h9696969696969696;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!nonposted_cmd_accepted1),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \last_channel[1]~0 (
	.dataa(!cmd_sink_data[77]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[1]~0 .extended_lut = "off";
defparam \last_channel[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_channel[1]~0 .shared_arith = "off";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[77]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

cyclonev_lcell_comb \last_dest_id[1]~0 (
	.dataa(!cmd_sink_channel[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_dest_id[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_dest_id[1]~0 .extended_lut = "off";
defparam \last_dest_id[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_dest_id[1]~0 .shared_arith = "off";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(\last_dest_id[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(\last_dest_id[1]~q ),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_cmd_demux (
	rst1,
	d_write,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_read,
	has_pending_responses,
	suppress_change_dest_id,
	av_waitrequest,
	always1,
	Equal4,
	Equal2,
	src_data_77,
	Equal1,
	mem_used_11,
	wait_latency_counter_11,
	wait_latency_counter_01,
	src_channel_3,
	Equal3,
	mem_used_12,
	wait_latency_counter_12,
	wait_latency_counter_02,
	saved_grant_0,
	mem_used_13,
	av_waitrequest1,
	mem_used_14,
	saved_grant_01,
	sink_ready,
	saved_grant_02,
	read_latency_shift_reg,
	WideOr01,
	cp_valid,
	last_channel_3,
	src3_valid,
	last_channel_2,
	src2_valid,
	src2_valid1,
	last_channel_6,
	src6_valid)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	d_write;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	d_read;
input 	has_pending_responses;
input 	suppress_change_dest_id;
input 	av_waitrequest;
input 	always1;
input 	Equal4;
input 	Equal2;
input 	src_data_77;
input 	Equal1;
input 	mem_used_11;
input 	wait_latency_counter_11;
input 	wait_latency_counter_01;
input 	src_channel_3;
input 	Equal3;
input 	mem_used_12;
input 	wait_latency_counter_12;
input 	wait_latency_counter_02;
input 	saved_grant_0;
input 	mem_used_13;
input 	av_waitrequest1;
input 	mem_used_14;
input 	saved_grant_01;
input 	sink_ready;
input 	saved_grant_02;
input 	read_latency_shift_reg;
output 	WideOr01;
input 	cp_valid;
input 	last_channel_3;
output 	src3_valid;
input 	last_channel_2;
output 	src2_valid;
output 	src2_valid1;
input 	last_channel_6;
output 	src6_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \sink_ready~1_combout ;
wire \sink_ready~2_combout ;
wire \sink_ready~3_combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \src3_valid~0_combout ;


cyclonev_lcell_comb WideOr0(
	.dataa(!\sink_ready~0_combout ),
	.datab(!src_channel_3),
	.datac(!\sink_ready~1_combout ),
	.datad(!\sink_ready~2_combout ),
	.datae(!\sink_ready~3_combout ),
	.dataf(!\WideOr0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \src3_valid~1 (
	.dataa(!av_waitrequest),
	.datab(!always1),
	.datac(!Equal4),
	.datad(!src_data_77),
	.datae(!Equal1),
	.dataf(!\src3_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~1 .extended_lut = "off";
defparam \src3_valid~1 .lut_mask = 64'hFFFF6996FFFFFFFF;
defparam \src3_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!has_pending_responses),
	.datae(!last_channel_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!Equal2),
	.datab(!src2_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'h7777777777777777;
defparam \src2_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~0 (
	.dataa(!Equal1),
	.datab(!suppress_change_dest_id),
	.datac(!cp_valid),
	.datad(!last_channel_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~0 .extended_lut = "off";
defparam \src6_valid~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \src6_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!mem_used_11),
	.datad(!always1),
	.datae(!wait_latency_counter_11),
	.dataf(!wait_latency_counter_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFFFFF7FFFFFFFDFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!rst1),
	.datad(!d_write),
	.datae(!mem_used_1),
	.dataf(!Equal3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hFFFFBFEFFFFFFFFF;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!Equal4),
	.datad(!mem_used_12),
	.datae(!wait_latency_counter_12),
	.dataf(!wait_latency_counter_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'hFFFFFF7FFFFFFFDF;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!rst1),
	.datab(!saved_grant_0),
	.datac(!mem_used_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!saved_grant_01),
	.datab(!sink_ready),
	.datac(!Equal2),
	.datad(!Equal1),
	.datae(!saved_grant_02),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!av_waitrequest),
	.datab(!av_waitrequest1),
	.datac(!mem_used_14),
	.datad(!\WideOr0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \src3_valid~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!has_pending_responses),
	.datae(!last_channel_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src3_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~0 .extended_lut = "off";
defparam \src3_valid~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \src3_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_cmd_demux_001 (
	WideOr0,
	rst1,
	mem_used_1,
	waitrequest,
	mem_used_11,
	sink_ready,
	has_pending_responses,
	i_read,
	src0_valid,
	last_channel_1,
	src_channel_1,
	src1_valid,
	saved_grant_1,
	Equal2,
	last_channel_0,
	src0_valid1,
	src0_valid2,
	saved_grant_11,
	Equal1,
	last_channel_2,
	src2_valid,
	mem)/* synthesis synthesis_greybox=1 */;
output 	WideOr0;
input 	rst1;
input 	mem_used_1;
input 	waitrequest;
input 	mem_used_11;
output 	sink_ready;
input 	has_pending_responses;
input 	i_read;
output 	src0_valid;
input 	last_channel_1;
input 	src_channel_1;
output 	src1_valid;
input 	saved_grant_1;
input 	Equal2;
input 	last_channel_0;
output 	src0_valid1;
output 	src0_valid2;
input 	saved_grant_11;
input 	Equal1;
input 	last_channel_2;
output 	src2_valid;
input 	mem;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~1_combout ;


cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!mem_used_1),
	.datab(!\sink_ready~1_combout ),
	.datac(!mem),
	.datad(!Equal2),
	.datae(!Equal1),
	.dataf(!rst1),
	.datag(!saved_grant_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "on";
defparam \WideOr0~0 .lut_mask = 64'hDDF5DDF5DDF5DDF5;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h7777777777777777;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!src0_valid),
	.datac(!last_channel_1),
	.datad(!src_channel_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!rst1),
	.datab(!last_channel_0),
	.datac(!has_pending_responses),
	.datad(!i_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \src0_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~2 (
	.dataa(!Equal2),
	.datab(!src0_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~2 .extended_lut = "off";
defparam \src0_valid~2 .lut_mask = 64'h7777777777777777;
defparam \src0_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!src0_valid),
	.datac(!Equal1),
	.datad(!last_channel_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!waitrequest),
	.datab(!mem_used_11),
	.datac(!saved_grant_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \sink_ready~1 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002 (
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	d_address_line_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_offset_field_1,
	r_sync_rst,
	Equal2,
	saved_grant_0,
	sink_ready,
	Equal21,
	src0_valid,
	src0_valid1,
	src2_valid,
	src2_valid1,
	saved_grant_1,
	WideOr11,
	hbreak_enabled,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	d_writedata_7,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_payload1,
	d_byteenable_0,
	src_data_32,
	d_writedata_3,
	src_payload2,
	d_writedata_1,
	src_payload3,
	d_writedata_4,
	d_writedata_20,
	d_byteenable_2,
	d_writedata_12,
	d_byteenable_1,
	d_writedata_28,
	d_byteenable_3,
	d_writedata_16,
	d_writedata_8,
	d_writedata_24,
	d_writedata_2,
	d_writedata_18,
	d_writedata_10,
	d_writedata_26,
	d_writedata_5,
	d_writedata_21,
	d_writedata_13,
	d_writedata_29,
	d_writedata_23,
	d_writedata_15,
	d_writedata_31,
	d_writedata_11,
	d_writedata_27,
	d_writedata_9,
	d_writedata_25,
	d_writedata_6,
	d_writedata_22,
	d_writedata_14,
	d_writedata_30,
	d_writedata_19,
	src_payload4,
	d_writedata_17,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_35,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_33,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	d_address_line_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_offset_field_1;
input 	r_sync_rst;
input 	Equal2;
output 	saved_grant_0;
input 	sink_ready;
input 	Equal21;
input 	src0_valid;
input 	src0_valid1;
input 	src2_valid;
input 	src2_valid1;
output 	saved_grant_1;
output 	WideOr11;
input 	hbreak_enabled;
input 	ic_fill_line_5;
output 	src_data_46;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_0;
input 	d_writedata_7;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
output 	src_data_45;
output 	src_data_44;
output 	src_data_43;
output 	src_data_42;
output 	src_payload1;
input 	d_byteenable_0;
output 	src_data_32;
input 	d_writedata_3;
output 	src_payload2;
input 	d_writedata_1;
output 	src_payload3;
input 	d_writedata_4;
input 	d_writedata_20;
input 	d_byteenable_2;
input 	d_writedata_12;
input 	d_byteenable_1;
input 	d_writedata_28;
input 	d_byteenable_3;
input 	d_writedata_16;
input 	d_writedata_8;
input 	d_writedata_24;
input 	d_writedata_2;
input 	d_writedata_18;
input 	d_writedata_10;
input 	d_writedata_26;
input 	d_writedata_5;
input 	d_writedata_21;
input 	d_writedata_13;
input 	d_writedata_29;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_31;
input 	d_writedata_11;
input 	d_writedata_27;
input 	d_writedata_9;
input 	d_writedata_25;
input 	d_writedata_6;
input 	d_writedata_22;
input 	d_writedata_14;
input 	d_writedata_30;
input 	d_writedata_19;
output 	src_payload4;
input 	d_writedata_17;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_data_35;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_data_33;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


Qsys_system_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.sink_ready(sink_ready),
	.src0_valid(src0_valid1),
	.src2_valid(src2_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_0),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(!src0_valid),
	.datae(!src2_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!d_address_line_field_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!d_address_offset_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!d_address_line_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!d_address_offset_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!d_address_offset_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!d_address_line_field_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!d_address_line_field_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!d_address_line_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!d_address_line_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!sink_ready),
	.datac(!\packet_in_progress~q ),
	.datad(!saved_grant_1),
	.datae(!WideOr11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF3FF77FFF3FF77FF;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	sink_ready,
	src0_valid,
	src2_valid,
	grant_0,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	sink_ready;
input 	src0_valid;
input 	src2_valid;
output 	grant_0;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src0_valid),
	.datad(!src2_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src0_valid),
	.datad(!src2_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!sink_ready),
	.datac(!src0_valid),
	.datad(!src2_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002_1 (
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	d_address_line_field_0,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_tag_field_3,
	d_address_tag_field_2,
	d_address_offset_field_1,
	r_sync_rst,
	saved_grant_0,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	src1_valid,
	src3_valid,
	read_latency_shift_reg,
	saved_grant_1,
	ic_fill_line_5,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	d_writedata_7,
	ic_fill_ap_offset_0,
	ic_fill_ap_offset_2,
	ic_fill_ap_offset_1,
	d_byteenable_0,
	d_writedata_3,
	d_writedata_1,
	d_writedata_4,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	d_writedata_20,
	src_payload1,
	d_byteenable_2,
	src_data_34,
	d_writedata_12,
	src_payload2,
	d_byteenable_1,
	src_data_33,
	d_writedata_28,
	src_payload3,
	d_byteenable_3,
	src_data_35,
	src_payload4,
	d_writedata_16,
	src_payload5,
	d_writedata_8,
	src_payload6,
	d_writedata_24,
	src_payload7,
	d_writedata_2,
	src_payload8,
	d_writedata_18,
	src_payload9,
	d_writedata_10,
	src_payload10,
	d_writedata_26,
	src_payload11,
	d_writedata_5,
	src_payload12,
	d_writedata_21,
	src_payload13,
	d_writedata_13,
	src_payload14,
	d_writedata_29,
	src_payload15,
	src_payload16,
	d_writedata_23,
	src_payload17,
	d_writedata_15,
	src_payload18,
	d_writedata_31,
	src_payload19,
	d_writedata_11,
	src_payload20,
	d_writedata_27,
	src_payload21,
	d_writedata_9,
	src_payload22,
	d_writedata_25,
	src_payload23,
	d_writedata_6,
	src_payload24,
	d_writedata_22,
	src_payload25,
	d_writedata_14,
	src_payload26,
	d_writedata_30,
	src_payload27,
	src_payload28,
	d_writedata_19,
	src_payload29,
	src_payload30,
	d_writedata_17,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	d_address_line_field_0;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_tag_field_3;
input 	d_address_tag_field_2;
input 	d_address_offset_field_1;
input 	r_sync_rst;
output 	saved_grant_0;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
input 	src1_valid;
input 	src3_valid;
input 	read_latency_shift_reg;
output 	saved_grant_1;
input 	ic_fill_line_5;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_0;
input 	d_writedata_7;
input 	ic_fill_ap_offset_0;
input 	ic_fill_ap_offset_2;
input 	ic_fill_ap_offset_1;
input 	d_byteenable_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	d_writedata_4;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_32;
input 	d_writedata_20;
output 	src_payload1;
input 	d_byteenable_2;
output 	src_data_34;
input 	d_writedata_12;
output 	src_payload2;
input 	d_byteenable_1;
output 	src_data_33;
input 	d_writedata_28;
output 	src_payload3;
input 	d_byteenable_3;
output 	src_data_35;
output 	src_payload4;
input 	d_writedata_16;
output 	src_payload5;
input 	d_writedata_8;
output 	src_payload6;
input 	d_writedata_24;
output 	src_payload7;
input 	d_writedata_2;
output 	src_payload8;
input 	d_writedata_18;
output 	src_payload9;
input 	d_writedata_10;
output 	src_payload10;
input 	d_writedata_26;
output 	src_payload11;
input 	d_writedata_5;
output 	src_payload12;
input 	d_writedata_21;
output 	src_payload13;
input 	d_writedata_13;
output 	src_payload14;
input 	d_writedata_29;
output 	src_payload15;
output 	src_payload16;
input 	d_writedata_23;
output 	src_payload17;
input 	d_writedata_15;
output 	src_payload18;
input 	d_writedata_31;
output 	src_payload19;
input 	d_writedata_11;
output 	src_payload20;
input 	d_writedata_27;
output 	src_payload21;
input 	d_writedata_9;
output 	src_payload22;
input 	d_writedata_25;
output 	src_payload23;
input 	d_writedata_6;
output 	src_payload24;
input 	d_writedata_22;
output 	src_payload25;
input 	d_writedata_14;
output 	src_payload26;
input 	d_writedata_30;
output 	src_payload27;
output 	src_payload28;
input 	d_writedata_19;
output 	src_payload29;
output 	src_payload30;
input 	d_writedata_17;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


Qsys_system_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.src1_valid(src1_valid),
	.src3_valid(src3_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!d_address_offset_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!d_address_offset_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!d_address_offset_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!d_address_line_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!d_address_line_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!d_address_line_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!d_address_line_field_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!d_address_line_field_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!d_address_line_field_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!d_address_tag_field_0),
	.datab(!saved_grant_0),
	.datac(!ic_fill_line_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!d_address_tag_field_1),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!d_address_tag_field_2),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!d_address_tag_field_3),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src1_valid),
	.datad(!src3_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	src1_valid,
	src3_valid,
	grant_0,
	read_latency_shift_reg,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	src1_valid;
input 	src3_valid;
output 	grant_0;
input 	read_latency_shift_reg;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src1_valid),
	.datad(!src3_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src1_valid),
	.datad(!src3_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src1_valid),
	.datad(!src3_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_cmd_mux_002_2 (
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	d_address_line_field_0,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_tag_field_2,
	d_address_offset_field_1,
	r_sync_rst,
	saved_grant_0,
	read_latency_shift_reg,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	src2_valid,
	src6_valid,
	saved_grant_1,
	ic_fill_line_5,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	d_writedata_7,
	ic_fill_ap_offset_0,
	ic_fill_ap_offset_2,
	ic_fill_ap_offset_1,
	d_byteenable_0,
	d_writedata_3,
	d_writedata_1,
	d_writedata_4,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_32,
	d_writedata_20,
	d_byteenable_2,
	src_payload1,
	src_data_34,
	d_writedata_12,
	d_byteenable_1,
	src_payload2,
	src_data_33,
	d_writedata_28,
	d_byteenable_3,
	src_payload3,
	src_data_35,
	src_payload4,
	d_writedata_16,
	src_payload5,
	d_writedata_8,
	src_payload6,
	d_writedata_24,
	src_payload7,
	d_writedata_2,
	src_payload8,
	d_writedata_18,
	src_payload9,
	d_writedata_10,
	src_payload10,
	d_writedata_26,
	src_payload11,
	d_writedata_5,
	src_payload12,
	d_writedata_21,
	src_payload13,
	d_writedata_13,
	src_payload14,
	d_writedata_29,
	src_payload15,
	src_payload16,
	d_writedata_23,
	src_payload17,
	d_writedata_15,
	src_payload18,
	d_writedata_31,
	src_payload19,
	d_writedata_11,
	src_payload20,
	d_writedata_27,
	src_payload21,
	d_writedata_9,
	src_payload22,
	d_writedata_25,
	src_payload23,
	d_writedata_6,
	src_payload24,
	d_writedata_22,
	src_payload25,
	d_writedata_14,
	src_payload26,
	d_writedata_30,
	src_payload27,
	src_payload28,
	d_writedata_19,
	src_payload29,
	src_payload30,
	d_writedata_17,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	d_address_line_field_0;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_tag_field_2;
input 	d_address_offset_field_1;
input 	r_sync_rst;
output 	saved_grant_0;
input 	read_latency_shift_reg;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
input 	src2_valid;
input 	src6_valid;
output 	saved_grant_1;
input 	ic_fill_line_5;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_0;
input 	d_writedata_7;
input 	ic_fill_ap_offset_0;
input 	ic_fill_ap_offset_2;
input 	ic_fill_ap_offset_1;
input 	d_byteenable_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	d_writedata_4;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_32;
input 	d_writedata_20;
input 	d_byteenable_2;
output 	src_payload1;
output 	src_data_34;
input 	d_writedata_12;
input 	d_byteenable_1;
output 	src_payload2;
output 	src_data_33;
input 	d_writedata_28;
input 	d_byteenable_3;
output 	src_payload3;
output 	src_data_35;
output 	src_payload4;
input 	d_writedata_16;
output 	src_payload5;
input 	d_writedata_8;
output 	src_payload6;
input 	d_writedata_24;
output 	src_payload7;
input 	d_writedata_2;
output 	src_payload8;
input 	d_writedata_18;
output 	src_payload9;
input 	d_writedata_10;
output 	src_payload10;
input 	d_writedata_26;
output 	src_payload11;
input 	d_writedata_5;
output 	src_payload12;
input 	d_writedata_21;
output 	src_payload13;
input 	d_writedata_13;
output 	src_payload14;
input 	d_writedata_29;
output 	src_payload15;
output 	src_payload16;
input 	d_writedata_23;
output 	src_payload17;
input 	d_writedata_15;
output 	src_payload18;
input 	d_writedata_31;
output 	src_payload19;
input 	d_writedata_11;
output 	src_payload20;
input 	d_writedata_27;
output 	src_payload21;
input 	d_writedata_9;
output 	src_payload22;
input 	d_writedata_25;
output 	src_payload23;
input 	d_writedata_6;
output 	src_payload24;
input 	d_writedata_22;
output 	src_payload25;
input 	d_writedata_14;
output 	src_payload26;
input 	d_writedata_30;
output 	src_payload27;
output 	src_payload28;
input 	d_writedata_19;
output 	src_payload29;
output 	src_payload30;
input 	d_writedata_17;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


Qsys_system_altera_merlin_arbitrator_2 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.src2_valid(src2_valid),
	.src6_valid(src6_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!d_address_offset_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!d_address_offset_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!d_address_offset_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!d_address_line_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!d_address_line_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!d_address_line_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!d_address_line_field_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!d_address_line_field_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!d_address_line_field_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!d_address_tag_field_0),
	.datab(!saved_grant_0),
	.datac(!ic_fill_line_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!d_address_tag_field_1),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!d_address_tag_field_2),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src2_valid),
	.datad(!src6_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_merlin_arbitrator_2 (
	reset,
	saved_grant_0,
	read_latency_shift_reg,
	src2_valid,
	src6_valid,
	grant_0,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	read_latency_shift_reg;
input 	src2_valid;
input 	src6_valid;
output 	grant_0;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src2_valid),
	.datad(!src6_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src2_valid),
	.datad(!src6_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src2_valid),
	.datad(!src6_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_router (
	d_address_offset_field_2,
	d_address_line_field_0,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	Equal3,
	d_address_line_field_1,
	d_address_tag_field_5,
	d_address_tag_field_4,
	d_address_tag_field_3,
	d_address_tag_field_2,
	Equal31,
	d_address_offset_field_1,
	d_read,
	av_waitrequest,
	always1,
	Equal4,
	Equal2,
	src_data_77,
	Equal1,
	src_data_771,
	src_data_79,
	src_channel_3,
	Equal32,
	src_data_78)/* synthesis synthesis_greybox=1 */;
input 	d_address_offset_field_2;
input 	d_address_line_field_0;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
output 	Equal3;
input 	d_address_line_field_1;
input 	d_address_tag_field_5;
input 	d_address_tag_field_4;
input 	d_address_tag_field_3;
input 	d_address_tag_field_2;
output 	Equal31;
input 	d_address_offset_field_1;
input 	d_read;
input 	av_waitrequest;
output 	always1;
output 	Equal4;
output 	Equal2;
output 	src_data_77;
output 	Equal1;
output 	src_data_771;
output 	src_data_79;
output 	src_channel_3;
output 	Equal32;
output 	src_data_78;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal3~0 (
	.dataa(!d_address_tag_field_1),
	.datab(!d_address_tag_field_0),
	.datac(!d_address_line_field_5),
	.datad(!d_address_line_field_4),
	.datae(!d_address_line_field_3),
	.dataf(!d_address_line_field_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!d_address_line_field_1),
	.datab(!d_address_tag_field_5),
	.datac(!d_address_tag_field_4),
	.datad(!d_address_tag_field_3),
	.datae(!d_address_tag_field_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_2),
	.datac(!d_address_line_field_0),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(!d_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!d_address_offset_field_2),
	.datab(!d_address_line_field_0),
	.datac(!Equal3),
	.datad(!Equal31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!d_address_tag_field_1),
	.datab(!d_address_tag_field_0),
	.datac(!d_address_tag_field_5),
	.datad(!d_address_tag_field_4),
	.datae(!d_address_tag_field_3),
	.dataf(!d_address_tag_field_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[77]~0 (
	.dataa(!d_address_line_field_0),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(!Equal2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77]~0 .extended_lut = "off";
defparam \src_data[77]~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \src_data[77]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!d_address_tag_field_5),
	.datab(!d_address_tag_field_4),
	.datac(!d_address_tag_field_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[77]~1 (
	.dataa(!av_waitrequest),
	.datab(!always1),
	.datac(!Equal4),
	.datad(!src_data_77),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_771),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77]~1 .extended_lut = "off";
defparam \src_data[77]~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[77]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[79]~2 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_2),
	.datac(!d_address_line_field_0),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(!d_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79]~2 .extended_lut = "off";
defparam \src_data[79]~2 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \src_data[79]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[3]~0 (
	.dataa(!av_waitrequest),
	.datab(!always1),
	.datac(!Equal4),
	.datad(!src_data_77),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[3]~0 .extended_lut = "off";
defparam \src_channel[3]~0 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \src_channel[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!d_address_line_field_0),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Equal3~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[78]~3 (
	.dataa(!av_waitrequest),
	.datab(!always1),
	.datac(!Equal4),
	.datad(!src_data_77),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78]~3 .extended_lut = "off";
defparam \src_data[78]~3 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \src_data[78]~3 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_router_001 (
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	src_channel_1,
	Equal2,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
output 	src_channel_1;
output 	Equal2;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src_channel[1]~0 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!ic_fill_tag_2),
	.datad(!ic_fill_tag_1),
	.datae(!ic_fill_tag_0),
	.dataf(!ic_fill_line_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[1]~0 .extended_lut = "off";
defparam \src_channel[1]~0 .lut_mask = 64'hFFFFFF7DFFFFFFFF;
defparam \src_channel[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!ic_fill_tag_2),
	.datad(!ic_fill_tag_1),
	.datae(!ic_fill_tag_0),
	.dataf(!ic_fill_line_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFF7FFFFFFFF;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!ic_fill_tag_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002_1 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_rsp_demux_002_2 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_rsp_mux (
	q_a_4,
	q_a_41,
	av_readdata_pre_4,
	q_a_20,
	q_a_201,
	av_readdata_pre_20,
	q_a_12,
	q_a_121,
	q_a_28,
	q_a_281,
	q_a_0,
	q_a_01,
	av_readdata_pre_0,
	q_a_16,
	q_a_161,
	av_readdata_pre_16,
	q_a_8,
	q_a_81,
	q_a_24,
	q_a_241,
	q_a_2,
	q_a_21,
	av_readdata_pre_2,
	q_a_18,
	q_a_181,
	av_readdata_pre_18,
	q_a_10,
	q_a_101,
	q_a_26,
	q_a_261,
	q_a_5,
	q_a_51,
	av_readdata_pre_5,
	q_a_211,
	q_a_212,
	av_readdata_pre_21,
	q_a_13,
	q_a_131,
	q_a_29,
	q_a_291,
	q_a_7,
	q_a_71,
	av_readdata_pre_7,
	q_a_23,
	q_a_231,
	q_a_15,
	q_a_151,
	q_a_31,
	q_a_311,
	q_a_11,
	q_a_111,
	q_a_27,
	q_a_271,
	q_a_9,
	q_a_91,
	q_a_25,
	q_a_251,
	q_a_6,
	q_a_61,
	av_readdata_pre_6,
	q_a_22,
	q_a_221,
	av_readdata_pre_22,
	q_a_14,
	q_a_141,
	q_a_30,
	q_a_301,
	q_a_3,
	q_a_32,
	av_readdata_pre_3,
	q_a_19,
	q_a_191,
	av_readdata_pre_19,
	q_a_1,
	q_a_17,
	av_readdata_pre_1,
	q_a_171,
	q_a_172,
	av_readdata_pre_17,
	read_latency_shift_reg_0,
	src0_valid,
	src0_valid1,
	src0_valid2,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	WideOr11,
	av_readdata_pre_30,
	av_readdata_pre_41,
	src_data_4,
	av_readdata_pre_201,
	src_data_20,
	av_readdata_pre_12,
	av_readdata_pre_121,
	src_data_12,
	av_readdata_pre_28,
	src_data_28,
	av_readdata_pre_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	src_data_0,
	av_readdata_pre_161,
	src_data_16,
	av_readdata_pre_8,
	av_readdata_pre_81,
	src_data_8,
	av_readdata_pre_24,
	src_data_24,
	av_readdata_pre_23,
	src_data_2,
	av_readdata_pre_181,
	src_data_18,
	av_readdata_pre_10,
	av_readdata_pre_101,
	src_data_10,
	av_readdata_pre_26,
	src_data_26,
	av_readdata_pre_51,
	src_data_5,
	av_readdata_pre_211,
	src_data_21,
	av_readdata_pre_13,
	av_readdata_pre_131,
	src_data_13,
	av_readdata_pre_29,
	src_data_29,
	av_readdata_pre_71,
	src_data_7,
	av_readdata_pre_231,
	src_data_23,
	av_readdata_pre_15,
	av_readdata_pre_151,
	src_data_15,
	av_readdata_pre_31,
	src_data_31,
	av_readdata_pre_11,
	src_data_11,
	av_readdata_pre_27,
	src_data_27,
	av_readdata_pre_9,
	av_readdata_pre_91,
	src_data_9,
	av_readdata_pre_25,
	src_data_25,
	av_readdata_pre_61,
	src_data_6,
	av_readdata_pre_221,
	src_data_22,
	av_readdata_pre_14,
	av_readdata_pre_141,
	src_data_14,
	av_readdata_pre_301,
	src_data_30,
	av_readdata_pre_32,
	src_data_3,
	av_readdata_pre_191,
	src_data_19,
	av_readdata_pre_110,
	src_data_1,
	av_readdata_pre_171,
	src_data_17)/* synthesis synthesis_greybox=1 */;
input 	q_a_4;
input 	q_a_41;
input 	av_readdata_pre_4;
input 	q_a_20;
input 	q_a_201;
input 	av_readdata_pre_20;
input 	q_a_12;
input 	q_a_121;
input 	q_a_28;
input 	q_a_281;
input 	q_a_0;
input 	q_a_01;
input 	av_readdata_pre_0;
input 	q_a_16;
input 	q_a_161;
input 	av_readdata_pre_16;
input 	q_a_8;
input 	q_a_81;
input 	q_a_24;
input 	q_a_241;
input 	q_a_2;
input 	q_a_21;
input 	av_readdata_pre_2;
input 	q_a_18;
input 	q_a_181;
input 	av_readdata_pre_18;
input 	q_a_10;
input 	q_a_101;
input 	q_a_26;
input 	q_a_261;
input 	q_a_5;
input 	q_a_51;
input 	av_readdata_pre_5;
input 	q_a_211;
input 	q_a_212;
input 	av_readdata_pre_21;
input 	q_a_13;
input 	q_a_131;
input 	q_a_29;
input 	q_a_291;
input 	q_a_7;
input 	q_a_71;
input 	av_readdata_pre_7;
input 	q_a_23;
input 	q_a_231;
input 	q_a_15;
input 	q_a_151;
input 	q_a_31;
input 	q_a_311;
input 	q_a_11;
input 	q_a_111;
input 	q_a_27;
input 	q_a_271;
input 	q_a_9;
input 	q_a_91;
input 	q_a_25;
input 	q_a_251;
input 	q_a_6;
input 	q_a_61;
input 	av_readdata_pre_6;
input 	q_a_22;
input 	q_a_221;
input 	av_readdata_pre_22;
input 	q_a_14;
input 	q_a_141;
input 	q_a_30;
input 	q_a_301;
input 	q_a_3;
input 	q_a_32;
input 	av_readdata_pre_3;
input 	q_a_19;
input 	q_a_191;
input 	av_readdata_pre_19;
input 	q_a_1;
input 	q_a_17;
input 	av_readdata_pre_1;
input 	q_a_171;
input 	q_a_172;
input 	av_readdata_pre_17;
input 	read_latency_shift_reg_0;
input 	src0_valid;
input 	src0_valid1;
input 	src0_valid2;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
output 	WideOr11;
input 	av_readdata_pre_30;
input 	av_readdata_pre_41;
output 	src_data_4;
input 	av_readdata_pre_201;
output 	src_data_20;
input 	av_readdata_pre_12;
input 	av_readdata_pre_121;
output 	src_data_12;
input 	av_readdata_pre_28;
output 	src_data_28;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
output 	src_data_0;
input 	av_readdata_pre_161;
output 	src_data_16;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
output 	src_data_8;
input 	av_readdata_pre_24;
output 	src_data_24;
input 	av_readdata_pre_23;
output 	src_data_2;
input 	av_readdata_pre_181;
output 	src_data_18;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
output 	src_data_10;
input 	av_readdata_pre_26;
output 	src_data_26;
input 	av_readdata_pre_51;
output 	src_data_5;
input 	av_readdata_pre_211;
output 	src_data_21;
input 	av_readdata_pre_13;
input 	av_readdata_pre_131;
output 	src_data_13;
input 	av_readdata_pre_29;
output 	src_data_29;
input 	av_readdata_pre_71;
output 	src_data_7;
input 	av_readdata_pre_231;
output 	src_data_23;
input 	av_readdata_pre_15;
input 	av_readdata_pre_151;
output 	src_data_15;
input 	av_readdata_pre_31;
output 	src_data_31;
input 	av_readdata_pre_11;
output 	src_data_11;
input 	av_readdata_pre_27;
output 	src_data_27;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
output 	src_data_9;
input 	av_readdata_pre_25;
output 	src_data_25;
input 	av_readdata_pre_61;
output 	src_data_6;
input 	av_readdata_pre_221;
output 	src_data_22;
input 	av_readdata_pre_14;
input 	av_readdata_pre_141;
output 	src_data_14;
input 	av_readdata_pre_301;
output 	src_data_30;
input 	av_readdata_pre_32;
output 	src_data_3;
input 	av_readdata_pre_191;
output 	src_data_19;
input 	av_readdata_pre_110;
output 	src_data_1;
input 	av_readdata_pre_171;
output 	src_data_17;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \src_payload~0_combout ;
wire \src_data[4]~0_combout ;
wire \src_data[20]~1_combout ;
wire \src_data[12]~2_combout ;
wire \src_data[28]~3_combout ;
wire \src_data[0]~4_combout ;
wire \src_data[0]~5_combout ;
wire \src_data[16]~6_combout ;
wire \src_data[8]~7_combout ;
wire \src_data[24]~8_combout ;
wire \src_data[2]~9_combout ;
wire \src_data[18]~10_combout ;
wire \src_data[10]~11_combout ;
wire \src_data[5]~12_combout ;
wire \src_data[21]~13_combout ;
wire \src_data[13]~14_combout ;
wire \src_data[7]~15_combout ;
wire \src_data[23]~16_combout ;
wire \src_data[15]~17_combout ;
wire \src_data[11]~18_combout ;
wire \src_data[27]~19_combout ;
wire \src_data[9]~20_combout ;
wire \src_data[6]~21_combout ;
wire \src_data[22]~22_combout ;
wire \src_data[14]~23_combout ;
wire \src_data[30]~24_combout ;
wire \src_data[3]~25_combout ;
wire \src_data[19]~26_combout ;
wire \src_data[1]~27_combout ;
wire \src_data[17]~28_combout ;


cyclonev_lcell_comb WideOr1(
	.dataa(!src0_valid2),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!\WideOr1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_4),
	.datad(!q_a_41),
	.datae(!\src_data[4]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_20),
	.datad(!q_a_201),
	.datae(!\src_data[20]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_12),
	.datad(!q_a_121),
	.datae(!\src_data[12]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_28),
	.datad(!q_a_281),
	.datae(!\src_data[28]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_0),
	.datad(!q_a_01),
	.datae(!\src_data[0]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_16),
	.datad(!q_a_161),
	.datae(!\src_data[16]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_8),
	.datad(!q_a_81),
	.datae(!\src_data[8]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_24),
	.datad(!q_a_241),
	.datae(!\src_data[24]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_2),
	.datad(!q_a_21),
	.datae(!\src_data[2]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_18),
	.datad(!q_a_181),
	.datae(!\src_data[18]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_10),
	.datad(!q_a_101),
	.datae(!\src_data[10]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src0_valid2),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_26),
	.datae(!q_a_26),
	.dataf(!q_a_261),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_5),
	.datad(!q_a_51),
	.datae(!\src_data[5]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_211),
	.datad(!q_a_212),
	.datae(!\src_data[21]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_13),
	.datad(!q_a_131),
	.datae(!\src_data[13]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src0_valid2),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_29),
	.datae(!q_a_29),
	.dataf(!q_a_291),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_7),
	.datad(!q_a_71),
	.datae(!\src_data[7]~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_23),
	.datad(!q_a_231),
	.datae(!\src_data[23]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_15),
	.datad(!q_a_151),
	.datae(!\src_data[15]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src0_valid2),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_31),
	.datae(!q_a_31),
	.dataf(!q_a_311),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_11),
	.datad(!q_a_111),
	.datae(!\src_data[11]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_27),
	.datad(!q_a_271),
	.datae(!\src_data[27]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_9),
	.datad(!q_a_91),
	.datae(!\src_data[9]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src0_valid2),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_25),
	.datae(!q_a_25),
	.dataf(!q_a_251),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_6),
	.datad(!q_a_61),
	.datae(!\src_data[6]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_22),
	.datad(!q_a_221),
	.datae(!\src_data[22]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_14),
	.datad(!q_a_141),
	.datae(!\src_data[14]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_30),
	.datad(!q_a_301),
	.datae(!\src_data[30]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_3),
	.datad(!q_a_32),
	.datae(!\src_data[3]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_19),
	.datad(!q_a_191),
	.datae(!\src_data[19]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[19] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_1),
	.datad(!q_a_17),
	.datae(!\src_data[1]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!q_a_171),
	.datad(!q_a_172),
	.datae(!\src_data[17]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!read_latency_shift_reg_02),
	.datad(!read_latency_shift_reg_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~0 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_4),
	.datae(!av_readdata_pre_41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~0 .extended_lut = "off";
defparam \src_data[4]~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~1 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_20),
	.datae(!av_readdata_pre_201),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[20]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~1 .extended_lut = "off";
defparam \src_data[20]~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[20]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~2 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_12),
	.datad(!av_readdata_pre_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[12]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~2 .extended_lut = "off";
defparam \src_data[12]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[12]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~3 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~3 .extended_lut = "off";
defparam \src_data[28]~3 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[28]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~4 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_0),
	.datad(!av_readdata_pre_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~4 .extended_lut = "off";
defparam \src_data[0]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~5 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_01),
	.datad(!av_readdata_pre_02),
	.datae(!\src_data[0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~5 .extended_lut = "off";
defparam \src_data[0]~5 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~6 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_16),
	.datad(!av_readdata_pre_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~6 .extended_lut = "off";
defparam \src_data[16]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[16]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~7 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_8),
	.datad(!av_readdata_pre_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~7 .extended_lut = "off";
defparam \src_data[8]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~8 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~8 .extended_lut = "off";
defparam \src_data[24]~8 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[24]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~9 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_2),
	.datad(!av_readdata_pre_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~9 .extended_lut = "off";
defparam \src_data[2]~9 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_18),
	.datad(!av_readdata_pre_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~10 .extended_lut = "off";
defparam \src_data[18]~10 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[18]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~11 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_10),
	.datae(!av_readdata_pre_101),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[10]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~11 .extended_lut = "off";
defparam \src_data[10]~11 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[10]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~12 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_5),
	.datad(!av_readdata_pre_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~12 .extended_lut = "off";
defparam \src_data[5]~12 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[5]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~13 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_21),
	.datae(!av_readdata_pre_211),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~13 .extended_lut = "off";
defparam \src_data[21]~13 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[21]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~14 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_13),
	.datad(!av_readdata_pre_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~14 .extended_lut = "off";
defparam \src_data[13]~14 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[13]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~15 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_7),
	.datae(!av_readdata_pre_71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~15 .extended_lut = "off";
defparam \src_data[7]~15 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[7]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~16 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_231),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~16 .extended_lut = "off";
defparam \src_data[23]~16 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[23]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~17 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_15),
	.datae(!av_readdata_pre_151),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[15]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~17 .extended_lut = "off";
defparam \src_data[15]~17 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[15]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~18 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[11]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~18 .extended_lut = "off";
defparam \src_data[11]~18 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[11]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~19 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~19 .extended_lut = "off";
defparam \src_data[27]~19 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[27]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~20 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_9),
	.datad(!av_readdata_pre_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~20 .extended_lut = "off";
defparam \src_data[9]~20 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~21 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_6),
	.datae(!av_readdata_pre_61),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~21 .extended_lut = "off";
defparam \src_data[6]~21 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[6]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~22 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_22),
	.datae(!av_readdata_pre_221),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[22]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~22 .extended_lut = "off";
defparam \src_data[22]~22 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[22]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~23 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_14),
	.datad(!av_readdata_pre_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[14]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~23 .extended_lut = "off";
defparam \src_data[14]~23 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[14]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~24 (
	.dataa(!src0_valid2),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_301),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~24 .extended_lut = "off";
defparam \src_data[30]~24 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_data[30]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~25 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_3),
	.datad(!av_readdata_pre_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~25 .extended_lut = "off";
defparam \src_data[3]~25 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~26 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!av_readdata_pre_19),
	.datad(!av_readdata_pre_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~26 .extended_lut = "off";
defparam \src_data[19]~26 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[19]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~27 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_110),
	.datae(!av_readdata_pre_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~27 .extended_lut = "off";
defparam \src_data[1]~27 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[1]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~28 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid2),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_17),
	.datae(!av_readdata_pre_171),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[17]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~28 .extended_lut = "off";
defparam \src_data[17]~28 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[17]~28 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_mm_interconnect_0_rsp_mux_001 (
	q_a_4,
	q_a_41,
	q_a_20,
	q_a_201,
	q_a_12,
	q_a_121,
	q_a_28,
	q_a_281,
	q_a_0,
	q_a_01,
	q_a_16,
	q_a_161,
	q_a_8,
	q_a_81,
	q_a_24,
	q_a_241,
	q_a_2,
	q_a_21,
	q_a_18,
	q_a_181,
	q_a_10,
	q_a_101,
	q_a_26,
	q_a_261,
	q_a_5,
	q_a_51,
	q_a_211,
	q_a_212,
	q_a_13,
	q_a_131,
	q_a_29,
	q_a_291,
	q_a_7,
	q_a_71,
	q_a_23,
	q_a_231,
	q_a_15,
	q_a_151,
	q_a_31,
	q_a_311,
	q_a_11,
	q_a_111,
	q_a_27,
	q_a_271,
	q_a_9,
	q_a_91,
	q_a_25,
	q_a_251,
	q_a_6,
	q_a_61,
	q_a_22,
	q_a_221,
	q_a_14,
	q_a_141,
	q_a_30,
	q_a_301,
	q_a_3,
	q_a_32,
	q_a_19,
	q_a_191,
	q_a_1,
	q_a_17,
	q_a_171,
	q_a_172,
	src1_valid,
	src1_valid1,
	src1_valid2,
	WideOr11,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_12,
	av_readdata_pre_28,
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_8,
	av_readdata_pre_24,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_10,
	av_readdata_pre_26,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_13,
	av_readdata_pre_29,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_11,
	av_readdata_pre_27,
	av_readdata_pre_9,
	av_readdata_pre_25,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_14,
	av_readdata_pre_30,
	av_readdata_pre_3,
	av_readdata_pre_19,
	src_data_5,
	src_data_3,
	av_readdata_pre_1,
	src_data_1,
	src_data_4,
	src_data_2,
	src_data_28,
	src_data_30,
	src_data_31,
	src_data_27,
	src_data_29,
	src_data_0,
	src_data_23,
	src_data_25,
	src_data_26,
	src_data_22,
	src_data_24,
	av_readdata_pre_17,
	src_data_16,
	src_data_15,
	src_data_13,
	src_data_14,
	src_data_12,
	src_data_11,
	src_data_10,
	src_data_8,
	src_data_18,
	src_data_17,
	src_data_21,
	src_data_6,
	src_data_20,
	src_data_19,
	src_data_9,
	src_data_7)/* synthesis synthesis_greybox=1 */;
input 	q_a_4;
input 	q_a_41;
input 	q_a_20;
input 	q_a_201;
input 	q_a_12;
input 	q_a_121;
input 	q_a_28;
input 	q_a_281;
input 	q_a_0;
input 	q_a_01;
input 	q_a_16;
input 	q_a_161;
input 	q_a_8;
input 	q_a_81;
input 	q_a_24;
input 	q_a_241;
input 	q_a_2;
input 	q_a_21;
input 	q_a_18;
input 	q_a_181;
input 	q_a_10;
input 	q_a_101;
input 	q_a_26;
input 	q_a_261;
input 	q_a_5;
input 	q_a_51;
input 	q_a_211;
input 	q_a_212;
input 	q_a_13;
input 	q_a_131;
input 	q_a_29;
input 	q_a_291;
input 	q_a_7;
input 	q_a_71;
input 	q_a_23;
input 	q_a_231;
input 	q_a_15;
input 	q_a_151;
input 	q_a_31;
input 	q_a_311;
input 	q_a_11;
input 	q_a_111;
input 	q_a_27;
input 	q_a_271;
input 	q_a_9;
input 	q_a_91;
input 	q_a_25;
input 	q_a_251;
input 	q_a_6;
input 	q_a_61;
input 	q_a_22;
input 	q_a_221;
input 	q_a_14;
input 	q_a_141;
input 	q_a_30;
input 	q_a_301;
input 	q_a_3;
input 	q_a_32;
input 	q_a_19;
input 	q_a_191;
input 	q_a_1;
input 	q_a_17;
input 	q_a_171;
input 	q_a_172;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
output 	WideOr11;
input 	av_readdata_pre_4;
input 	av_readdata_pre_20;
input 	av_readdata_pre_12;
input 	av_readdata_pre_28;
input 	av_readdata_pre_0;
input 	av_readdata_pre_16;
input 	av_readdata_pre_8;
input 	av_readdata_pre_24;
input 	av_readdata_pre_2;
input 	av_readdata_pre_18;
input 	av_readdata_pre_10;
input 	av_readdata_pre_26;
input 	av_readdata_pre_5;
input 	av_readdata_pre_21;
input 	av_readdata_pre_13;
input 	av_readdata_pre_29;
input 	av_readdata_pre_7;
input 	av_readdata_pre_23;
input 	av_readdata_pre_15;
input 	av_readdata_pre_31;
input 	av_readdata_pre_11;
input 	av_readdata_pre_27;
input 	av_readdata_pre_9;
input 	av_readdata_pre_25;
input 	av_readdata_pre_6;
input 	av_readdata_pre_22;
input 	av_readdata_pre_14;
input 	av_readdata_pre_30;
input 	av_readdata_pre_3;
input 	av_readdata_pre_19;
output 	src_data_5;
output 	src_data_3;
input 	av_readdata_pre_1;
output 	src_data_1;
output 	src_data_4;
output 	src_data_2;
output 	src_data_28;
output 	src_data_30;
output 	src_data_31;
output 	src_data_27;
output 	src_data_29;
output 	src_data_0;
output 	src_data_23;
output 	src_data_25;
output 	src_data_26;
output 	src_data_22;
output 	src_data_24;
input 	av_readdata_pre_17;
output 	src_data_16;
output 	src_data_15;
output 	src_data_13;
output 	src_data_14;
output 	src_data_12;
output 	src_data_11;
output 	src_data_10;
output 	src_data_8;
output 	src_data_18;
output 	src_data_17;
output 	src_data_21;
output 	src_data_6;
output 	src_data_20;
output 	src_data_19;
output 	src_data_9;
output 	src_data_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_5),
	.datae(!q_a_5),
	.dataf(!q_a_51),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_3),
	.datae(!q_a_3),
	.dataf(!q_a_32),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_1),
	.datae(!q_a_1),
	.dataf(!q_a_17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_4),
	.datae(!q_a_4),
	.dataf(!q_a_41),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_2),
	.datae(!q_a_2),
	.dataf(!q_a_21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_28),
	.datae(!q_a_28),
	.dataf(!q_a_281),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_30),
	.datae(!q_a_30),
	.dataf(!q_a_301),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_31),
	.datae(!q_a_31),
	.dataf(!q_a_311),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_27),
	.datae(!q_a_27),
	.dataf(!q_a_271),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_29),
	.datae(!q_a_29),
	.dataf(!q_a_291),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_0),
	.datae(!q_a_0),
	.dataf(!q_a_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_23),
	.datae(!q_a_23),
	.dataf(!q_a_231),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_25),
	.datae(!q_a_25),
	.dataf(!q_a_251),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_26),
	.datae(!q_a_26),
	.dataf(!q_a_261),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_22),
	.datae(!q_a_22),
	.dataf(!q_a_221),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_24),
	.datae(!q_a_24),
	.dataf(!q_a_241),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_16),
	.datae(!q_a_16),
	.dataf(!q_a_161),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_15),
	.datae(!q_a_15),
	.dataf(!q_a_151),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_13),
	.datae(!q_a_13),
	.dataf(!q_a_131),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_14),
	.datae(!q_a_14),
	.dataf(!q_a_141),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_12),
	.datae(!q_a_12),
	.dataf(!q_a_121),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_11),
	.datae(!q_a_11),
	.dataf(!q_a_111),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_10),
	.datae(!q_a_10),
	.dataf(!q_a_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_8),
	.datae(!q_a_8),
	.dataf(!q_a_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_18),
	.datae(!q_a_18),
	.dataf(!q_a_181),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_17),
	.datae(!q_a_171),
	.dataf(!q_a_172),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_21),
	.datae(!q_a_211),
	.dataf(!q_a_212),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_6),
	.datae(!q_a_6),
	.dataf(!q_a_61),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_20),
	.datae(!q_a_20),
	.dataf(!q_a_201),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_19),
	.datae(!q_a_19),
	.dataf(!q_a_191),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[19] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_9),
	.datae(!q_a_9),
	.dataf(!q_a_91),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!av_readdata_pre_7),
	.datae(!q_a_7),
	.dataf(!q_a_71),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[7] .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0 (
	readdata_4,
	readdata_20,
	readdata_12,
	readdata_28,
	readdata_16,
	readdata_8,
	readdata_24,
	readdata_2,
	readdata_18,
	readdata_10,
	readdata_26,
	readdata_5,
	readdata_21,
	readdata_13,
	readdata_29,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_11,
	readdata_27,
	readdata_9,
	readdata_25,
	readdata_6,
	readdata_22,
	readdata_14,
	readdata_30,
	readdata_3,
	readdata_19,
	readdata_17,
	WideOr0,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	rst1,
	d_write1,
	d_address_line_field_0,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_tag_field_5,
	d_address_tag_field_4,
	d_address_tag_field_3,
	d_address_tag_field_2,
	d_address_offset_field_1,
	r_sync_rst,
	d_read1,
	av_begintransfer,
	suppress_change_dest_id,
	saved_grant_0,
	jtag_debug_module_waitrequest,
	mem_used_1,
	WideOr01,
	av_waitrequest,
	d_readdatavalid,
	has_pending_responses,
	i_read1,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	WideOr1,
	rf_source_valid,
	hbreak_enabled1,
	save_dest_id,
	nonposted_cmd_accepted,
	suppress_change_dest_id1,
	ic_fill_line_5,
	src_data_46,
	r_early_rst,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	d_writedata_7,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_payload1,
	d_byteenable_0,
	src_data_32,
	WideOr11,
	av_readdata_9,
	av_readdata_8,
	irq_mask,
	edge_capture,
	d_writedata_3,
	src_payload2,
	d_readdata,
	d_writedata_1,
	src_payload3,
	i_readdata,
	d_writedata_4,
	d_writedata_20,
	d_byteenable_2,
	d_writedata_12,
	d_byteenable_1,
	d_writedata_28,
	d_byteenable_3,
	readdata_0,
	d_writedata_16,
	d_writedata_8,
	d_writedata_24,
	d_writedata_2,
	d_writedata_18,
	d_writedata_10,
	d_writedata_26,
	d_writedata_5,
	d_writedata_21,
	d_writedata_13,
	d_writedata_29,
	d_writedata_23,
	d_writedata_15,
	d_writedata_31,
	d_writedata_11,
	d_writedata_27,
	d_writedata_9,
	d_writedata_25,
	d_writedata_6,
	d_writedata_22,
	d_writedata_14,
	d_writedata_30,
	d_writedata_19,
	jtag_debug_module_resetrequest,
	src_payload4,
	readdata_1,
	d_writedata_17,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_35,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_33,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_4;
output 	readdata_20;
output 	readdata_12;
output 	readdata_28;
output 	readdata_16;
output 	readdata_8;
output 	readdata_24;
output 	readdata_2;
output 	readdata_18;
output 	readdata_10;
output 	readdata_26;
output 	readdata_5;
output 	readdata_21;
output 	readdata_13;
output 	readdata_29;
output 	readdata_7;
output 	readdata_23;
output 	readdata_15;
output 	readdata_31;
output 	readdata_11;
output 	readdata_27;
output 	readdata_9;
output 	readdata_25;
output 	readdata_6;
output 	readdata_22;
output 	readdata_14;
output 	readdata_30;
output 	readdata_3;
output 	readdata_19;
output 	readdata_17;
input 	WideOr0;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	d_address_offset_field_2;
output 	d_writedata_0;
output 	d_address_offset_field_0;
input 	rst1;
output 	d_write1;
output 	d_address_line_field_0;
output 	d_address_tag_field_1;
output 	d_address_tag_field_0;
output 	d_address_line_field_5;
output 	d_address_line_field_4;
output 	d_address_line_field_3;
output 	d_address_line_field_2;
output 	d_address_line_field_1;
output 	d_address_tag_field_5;
output 	d_address_tag_field_4;
output 	d_address_tag_field_3;
output 	d_address_tag_field_2;
output 	d_address_offset_field_1;
input 	r_sync_rst;
output 	d_read1;
input 	av_begintransfer;
input 	suppress_change_dest_id;
input 	saved_grant_0;
output 	jtag_debug_module_waitrequest;
input 	mem_used_1;
input 	WideOr01;
input 	av_waitrequest;
input 	d_readdatavalid;
input 	has_pending_responses;
output 	i_read1;
output 	ic_fill_tag_4;
output 	ic_fill_tag_3;
output 	ic_fill_tag_2;
output 	ic_fill_tag_1;
output 	ic_fill_tag_0;
output 	ic_fill_line_6;
input 	WideOr1;
input 	rf_source_valid;
output 	hbreak_enabled1;
input 	save_dest_id;
input 	nonposted_cmd_accepted;
input 	suppress_change_dest_id1;
output 	ic_fill_line_5;
input 	src_data_46;
input 	r_early_rst;
output 	ic_fill_line_4;
output 	ic_fill_line_3;
output 	ic_fill_line_1;
output 	ic_fill_line_2;
output 	ic_fill_line_0;
output 	d_writedata_7;
input 	src_payload;
output 	ic_fill_ap_offset_0;
input 	src_data_38;
input 	src_data_41;
output 	ic_fill_ap_offset_2;
input 	src_data_40;
output 	ic_fill_ap_offset_1;
input 	src_data_39;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_payload1;
output 	d_byteenable_0;
input 	src_data_32;
input 	WideOr11;
input 	av_readdata_9;
input 	av_readdata_8;
input 	irq_mask;
input 	edge_capture;
output 	d_writedata_3;
input 	src_payload2;
input 	[31:0] d_readdata;
output 	d_writedata_1;
input 	src_payload3;
input 	[31:0] i_readdata;
output 	d_writedata_4;
output 	d_writedata_20;
output 	d_byteenable_2;
output 	d_writedata_12;
output 	d_byteenable_1;
output 	d_writedata_28;
output 	d_byteenable_3;
output 	readdata_0;
output 	d_writedata_16;
output 	d_writedata_8;
output 	d_writedata_24;
output 	d_writedata_2;
output 	d_writedata_18;
output 	d_writedata_10;
output 	d_writedata_26;
output 	d_writedata_5;
output 	d_writedata_21;
output 	d_writedata_13;
output 	d_writedata_29;
output 	d_writedata_23;
output 	d_writedata_15;
output 	d_writedata_31;
output 	d_writedata_11;
output 	d_writedata_27;
output 	d_writedata_9;
output 	d_writedata_25;
output 	d_writedata_6;
output 	d_writedata_22;
output 	d_writedata_14;
output 	d_writedata_30;
output 	d_writedata_19;
output 	jtag_debug_module_resetrequest;
input 	src_payload4;
output 	readdata_1;
output 	d_writedata_17;
input 	src_payload5;
input 	src_data_34;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_data_35;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_33;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \A_dc_xfer_wr_data[0]~q ;
wire \Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[7] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ;
wire \Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ;
wire \Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~1_sumout ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ;
wire \ic_fill_valid_bits[5]~q ;
wire \ic_fill_valid_bits[7]~q ;
wire \ic_fill_valid_bits[4]~q ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ;
wire \ic_fill_valid_bits[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~5_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~9_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~13_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~17_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~21_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~25_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~29_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~33_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~37_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~41_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~45_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~49_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~53_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~57_sumout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|Add0~61_sumout ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ;
wire \A_dc_xfer_wr_data[7]~q ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ;
wire \ic_fill_valid_bits[1]~q ;
wire \ic_fill_valid_bits[3]~q ;
wire \ic_fill_valid_bits[0]~q ;
wire \ic_fill_valid_bits[2]~q ;
wire \A_dc_xfer_wr_data[3]~q ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ;
wire \A_mul_src2[0]~q ;
wire \A_mul_src2[1]~q ;
wire \A_mul_src2[2]~q ;
wire \A_mul_src2[3]~q ;
wire \A_mul_src2[4]~q ;
wire \A_mul_src2[5]~q ;
wire \A_mul_src2[6]~q ;
wire \A_mul_src2[7]~q ;
wire \A_mul_src2[8]~q ;
wire \A_mul_src2[9]~q ;
wire \A_mul_src2[10]~q ;
wire \A_mul_src2[11]~q ;
wire \A_mul_src2[12]~q ;
wire \A_mul_src2[13]~q ;
wire \A_mul_src2[14]~q ;
wire \A_mul_src2[15]~q ;
wire \A_mul_src1[0]~q ;
wire \A_mul_src1[1]~q ;
wire \A_mul_src1[2]~q ;
wire \A_mul_src1[3]~q ;
wire \A_mul_src1[4]~q ;
wire \A_mul_src1[5]~q ;
wire \A_mul_src1[6]~q ;
wire \A_mul_src1[7]~q ;
wire \A_mul_src1[8]~q ;
wire \A_mul_src1[9]~q ;
wire \A_mul_src1[10]~q ;
wire \A_mul_src1[11]~q ;
wire \A_mul_src1[12]~q ;
wire \A_mul_src1[13]~q ;
wire \A_mul_src1[14]~q ;
wire \A_mul_src1[15]~q ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ;
wire \A_dc_xfer_wr_data[1]~q ;
wire \Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ;
wire \A_dc_xfer_wr_data[4]~q ;
wire \A_dc_xfer_wr_data[20]~q ;
wire \A_dc_xfer_wr_data[12]~q ;
wire \A_dc_xfer_wr_data[28]~q ;
wire \A_mul_src2[16]~q ;
wire \A_mul_src2[17]~q ;
wire \A_mul_src2[18]~q ;
wire \A_mul_src2[19]~q ;
wire \A_mul_src2[20]~q ;
wire \A_mul_src2[21]~q ;
wire \A_mul_src2[22]~q ;
wire \A_mul_src2[23]~q ;
wire \A_mul_src2[24]~q ;
wire \A_mul_src2[25]~q ;
wire \A_mul_src2[26]~q ;
wire \A_mul_src2[27]~q ;
wire \A_mul_src2[28]~q ;
wire \A_mul_src2[29]~q ;
wire \A_mul_src2[30]~q ;
wire \A_mul_src2[31]~q ;
wire \Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ;
wire \A_dc_xfer_wr_data[16]~q ;
wire \A_dc_xfer_wr_data[8]~q ;
wire \A_dc_xfer_wr_data[24]~q ;
wire \A_dc_xfer_wr_data[2]~q ;
wire \A_dc_xfer_wr_data[18]~q ;
wire \A_dc_xfer_wr_data[10]~q ;
wire \A_dc_xfer_wr_data[26]~q ;
wire \A_dc_xfer_wr_data[5]~q ;
wire \A_dc_xfer_wr_data[21]~q ;
wire \A_dc_xfer_wr_data[13]~q ;
wire \A_dc_xfer_wr_data[29]~q ;
wire \A_dc_xfer_wr_data[23]~q ;
wire \A_dc_xfer_wr_data[15]~q ;
wire \A_dc_xfer_wr_data[31]~q ;
wire \A_dc_xfer_wr_data[11]~q ;
wire \A_dc_xfer_wr_data[27]~q ;
wire \A_dc_xfer_wr_data[9]~q ;
wire \A_dc_xfer_wr_data[25]~q ;
wire \A_dc_xfer_wr_data[6]~q ;
wire \A_dc_xfer_wr_data[22]~q ;
wire \A_dc_xfer_wr_data[14]~q ;
wire \A_dc_xfer_wr_data[30]~q ;
wire \A_mul_src1[16]~q ;
wire \A_mul_src1[17]~q ;
wire \A_mul_src1[18]~q ;
wire \A_mul_src1[19]~q ;
wire \A_mul_src1[20]~q ;
wire \A_mul_src1[21]~q ;
wire \A_mul_src1[22]~q ;
wire \A_mul_src1[23]~q ;
wire \A_mul_src1[24]~q ;
wire \A_mul_src1[25]~q ;
wire \A_mul_src1[26]~q ;
wire \A_mul_src1[27]~q ;
wire \A_mul_src1[28]~q ;
wire \A_mul_src1[29]~q ;
wire \A_mul_src1[30]~q ;
wire \A_mul_src1[31]~q ;
wire \A_dc_xfer_wr_data[19]~q ;
wire \A_dc_xfer_wr_data[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ;
wire \A_dc_xfer_wr_active~q ;
wire \A_dc_wb_rd_en~0_combout ;
wire \A_dc_wb_rd_en~combout ;
wire \A_dc_xfer_wr_offset[0]~q ;
wire \A_dc_xfer_wr_offset[1]~q ;
wire \A_dc_xfer_wr_offset[2]~q ;
wire \A_dc_wb_rd_addr_offset[0]~q ;
wire \A_dc_wb_rd_addr_offset[1]~q ;
wire \A_dc_wb_rd_addr_offset[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ;
wire \A_dc_fill_starting_d1~q ;
wire \A_en_d1~q ;
wire \A_ctrl_dc_index_inv~q ;
wire \A_ctrl_dc_addr_inv~q ;
wire \A_dc_tag_dcache_management_wr_en~0_combout ;
wire \dc_tag_wr_port_data[5]~0_combout ;
wire \dc_tag_wr_port_en~combout ;
wire \dc_tag_wr_port_data[4]~1_combout ;
wire \dc_tag_wr_port_addr[0]~0_combout ;
wire \dc_tag_wr_port_addr[1]~1_combout ;
wire \dc_tag_wr_port_addr[2]~2_combout ;
wire \dc_tag_wr_port_addr[3]~3_combout ;
wire \dc_tag_wr_port_addr[4]~4_combout ;
wire \dc_tag_wr_port_addr[5]~5_combout ;
wire \dc_tag_rd_port_addr[0]~0_combout ;
wire \dc_tag_rd_port_addr[1]~1_combout ;
wire \dc_tag_rd_port_addr[2]~2_combout ;
wire \dc_tag_rd_port_addr[3]~3_combout ;
wire \dc_tag_rd_port_addr[4]~4_combout ;
wire \dc_tag_rd_port_addr[5]~5_combout ;
wire \dc_tag_wr_port_data[5]~2_combout ;
wire \dc_tag_wr_port_data[6]~3_combout ;
wire \dc_tag_wr_port_data[0]~4_combout ;
wire \dc_tag_wr_port_data[1]~5_combout ;
wire \dc_tag_wr_port_data[2]~6_combout ;
wire \dc_tag_wr_port_data[3]~7_combout ;
wire \A_dc_xfer_rd_data_active~q ;
wire \A_dc_rd_data[0]~q ;
wire \A_dc_xfer_rd_data_offset_match~q ;
wire \A_dc_xfer_wr_offset_nxt[0]~0_combout ;
wire \A_dc_xfer_wr_offset_nxt[1]~1_combout ;
wire \A_dc_xfer_wr_offset_nxt[2]~2_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[0]~0_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[1]~1_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[2]~2_combout ;
wire \M_ctrl_dc_index_inv~q ;
wire \M_ctrl_dc_addr_inv~q ;
wire \A_valid_st_writes_mem~q ;
wire \dc_tag_wr_port_data[7]~8_combout ;
wire \rf_b_rd_port_addr[0]~0_combout ;
wire \rf_b_rd_port_addr[1]~1_combout ;
wire \rf_b_rd_port_addr[2]~2_combout ;
wire \rf_b_rd_port_addr[3]~3_combout ;
wire \rf_b_rd_port_addr[4]~4_combout ;
wire \rf_a_rd_port_addr[0]~0_combout ;
wire \rf_a_rd_port_addr[1]~1_combout ;
wire \rf_a_rd_port_addr[2]~2_combout ;
wire \rf_a_rd_port_addr[3]~3_combout ;
wire \rf_a_rd_port_addr[4]~4_combout ;
wire \A_dc_valid_st_bypass_hit_wr_en~combout ;
wire \dc_data_wr_port_en~combout ;
wire \M_dc_st_data[0]~0_combout ;
wire \A_dc_st_data[0]~q ;
wire \A_ctrl_st~q ;
wire \dc_data_wr_port_data[6]~0_combout ;
wire \dc_data_wr_port_data[0]~1_combout ;
wire \dc_data_wr_port_addr[0]~0_combout ;
wire \dc_data_wr_port_addr[1]~1_combout ;
wire \dc_data_wr_port_addr[2]~2_combout ;
wire \dc_data_wr_port_addr[3]~3_combout ;
wire \dc_data_wr_port_addr[4]~4_combout ;
wire \dc_data_wr_port_addr[5]~5_combout ;
wire \dc_data_wr_port_addr[6]~6_combout ;
wire \dc_data_wr_port_addr[7]~7_combout ;
wire \dc_data_wr_port_addr[8]~8_combout ;
wire \dc_data_rd_port_addr[0]~0_combout ;
wire \dc_data_rd_port_addr[1]~1_combout ;
wire \dc_data_rd_port_addr[2]~2_combout ;
wire \dc_data_rd_port_addr[3]~3_combout ;
wire \dc_data_rd_port_addr[4]~4_combout ;
wire \dc_data_rd_port_addr[5]~5_combout ;
wire \dc_data_rd_port_addr[6]~6_combout ;
wire \dc_data_rd_port_addr[7]~7_combout ;
wire \dc_data_rd_port_addr[8]~8_combout ;
wire \A_dc_xfer_rd_addr_offset_match~0_combout ;
wire \A_dc_xfer_rd_addr_offset_match~combout ;
wire \ic_tag_clr_valid_bits~q ;
wire \ic_tag_wren~combout ;
wire \ic_tag_wraddress[0]~q ;
wire \ic_tag_wraddress[1]~q ;
wire \ic_tag_wraddress[2]~q ;
wire \ic_tag_wraddress[3]~q ;
wire \ic_tag_wraddress[4]~q ;
wire \ic_tag_wraddress[5]~q ;
wire \ic_tag_wraddress[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[1]~q ;
wire \i_readdata_d1[5]~q ;
wire \i_readdata_d1[3]~q ;
wire \i_readdata_d1[1]~q ;
wire \i_readdata_d1[4]~q ;
wire \i_readdata_d1[2]~q ;
wire \i_readdata_d1[28]~q ;
wire \i_readdata_d1[30]~q ;
wire \i_readdata_d1[31]~q ;
wire \i_readdata_d1[27]~q ;
wire \i_readdata_d1[29]~q ;
wire \i_readdata_d1[0]~q ;
wire \i_readdata_d1[23]~q ;
wire \i_readdata_d1[25]~q ;
wire \i_readdata_d1[26]~q ;
wire \i_readdata_d1[22]~q ;
wire \i_readdata_d1[24]~q ;
wire \i_readdata_d1[16]~q ;
wire \i_readdata_d1[15]~q ;
wire \i_readdata_d1[13]~q ;
wire \i_readdata_d1[14]~q ;
wire \i_readdata_d1[12]~q ;
wire \i_readdata_d1[11]~q ;
wire \E_ctrl_dc_index_inv~0_combout ;
wire \M_ctrl_st~q ;
wire \M_valid_st_writes_mem~combout ;
wire \i_readdata_d1[10]~q ;
wire \M_dc_st_data[4]~1_combout ;
wire \A_dc_st_data[4]~q ;
wire \dc_data_wr_port_data[4]~2_combout ;
wire \M_dc_st_data[20]~2_combout ;
wire \A_dc_st_data[20]~q ;
wire \dc_data_wr_port_data[18]~3_combout ;
wire \dc_data_wr_port_data[20]~4_combout ;
wire \M_dc_st_data[12]~3_combout ;
wire \A_dc_st_data[12]~q ;
wire \dc_data_wr_port_data[12]~5_combout ;
wire \dc_data_wr_port_data[12]~6_combout ;
wire \M_dc_st_data[28]~4_combout ;
wire \A_dc_st_data[28]~q ;
wire \dc_data_wr_port_data[31]~7_combout ;
wire \dc_data_wr_port_data[28]~8_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \M_ctrl_br_cond~q ;
wire \M_bht_wr_en_unfiltered~combout ;
wire \M_bht_data[1]~q ;
wire \M_bht_data[0]~q ;
wire \M_br_mispredict~q ;
wire \M_bht_wr_data_unfiltered[1]~0_combout ;
wire \M_bht_ptr_unfiltered[0]~q ;
wire \M_bht_ptr_unfiltered[1]~q ;
wire \M_bht_ptr_unfiltered[2]~q ;
wire \M_bht_ptr_unfiltered[3]~q ;
wire \M_bht_ptr_unfiltered[4]~q ;
wire \M_bht_ptr_unfiltered[5]~q ;
wire \M_bht_ptr_unfiltered[6]~q ;
wire \M_bht_ptr_unfiltered[7]~q ;
wire \M_br_cond_taken_history[0]~q ;
wire \F_bht_ptr_nxt[0]~combout ;
wire \M_br_cond_taken_history[1]~q ;
wire \F_bht_ptr_nxt[1]~combout ;
wire \M_br_cond_taken_history[2]~q ;
wire \F_bht_ptr_nxt[2]~combout ;
wire \M_br_cond_taken_history[3]~q ;
wire \F_bht_ptr_nxt[3]~combout ;
wire \M_br_cond_taken_history[4]~q ;
wire \F_bht_ptr_nxt[4]~combout ;
wire \M_br_cond_taken_history[5]~q ;
wire \F_bht_ptr_nxt[5]~combout ;
wire \M_br_cond_taken_history[6]~q ;
wire \F_bht_ptr_nxt[6]~combout ;
wire \M_br_cond_taken_history[7]~q ;
wire \F_bht_ptr_nxt[7]~combout ;
wire \M_dc_st_data[16]~5_combout ;
wire \A_dc_st_data[16]~q ;
wire \dc_data_wr_port_data[16]~9_combout ;
wire \M_dc_st_data[8]~6_combout ;
wire \A_dc_st_data[8]~q ;
wire \dc_data_wr_port_data[8]~10_combout ;
wire \M_dc_st_data[24]~7_combout ;
wire \A_dc_st_data[24]~q ;
wire \dc_data_wr_port_data[24]~11_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \i_readdata_d1[8]~q ;
wire \M_dc_st_data[2]~8_combout ;
wire \A_dc_st_data[2]~q ;
wire \dc_data_wr_port_data[2]~12_combout ;
wire \M_dc_st_data[18]~9_combout ;
wire \A_dc_st_data[18]~q ;
wire \dc_data_wr_port_data[18]~13_combout ;
wire \M_dc_st_data[10]~10_combout ;
wire \A_dc_st_data[10]~q ;
wire \dc_data_wr_port_data[10]~14_combout ;
wire \M_dc_st_data[26]~11_combout ;
wire \A_dc_st_data[26]~q ;
wire \dc_data_wr_port_data[26]~15_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \M_dc_st_data[5]~12_combout ;
wire \A_dc_st_data[5]~q ;
wire \dc_data_wr_port_data[5]~16_combout ;
wire \M_dc_st_data[21]~13_combout ;
wire \A_dc_st_data[21]~q ;
wire \dc_data_wr_port_data[21]~17_combout ;
wire \M_dc_st_data[13]~14_combout ;
wire \A_dc_st_data[13]~q ;
wire \dc_data_wr_port_data[13]~18_combout ;
wire \M_dc_st_data[29]~15_combout ;
wire \A_dc_st_data[29]~q ;
wire \dc_data_wr_port_data[29]~19_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \i_readdata_d1[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \M_dc_st_data[7]~16_combout ;
wire \A_dc_st_data[7]~q ;
wire \dc_data_wr_port_data[7]~20_combout ;
wire \M_dc_st_data[23]~17_combout ;
wire \A_dc_st_data[23]~q ;
wire \dc_data_wr_port_data[23]~21_combout ;
wire \M_dc_st_data[15]~18_combout ;
wire \A_dc_st_data[15]~q ;
wire \dc_data_wr_port_data[15]~22_combout ;
wire \M_dc_st_data[31]~19_combout ;
wire \A_dc_st_data[31]~q ;
wire \dc_data_wr_port_data[31]~23_combout ;
wire \i_readdata_d1[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \M_dc_st_data[11]~20_combout ;
wire \A_dc_st_data[11]~q ;
wire \dc_data_wr_port_data[11]~24_combout ;
wire \M_dc_st_data[27]~21_combout ;
wire \A_dc_st_data[27]~q ;
wire \dc_data_wr_port_data[27]~25_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \M_dc_st_data[9]~22_combout ;
wire \A_dc_st_data[9]~q ;
wire \dc_data_wr_port_data[9]~26_combout ;
wire \M_dc_st_data[25]~23_combout ;
wire \A_dc_st_data[25]~q ;
wire \dc_data_wr_port_data[25]~27_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \M_dc_st_data[6]~24_combout ;
wire \A_dc_st_data[6]~q ;
wire \dc_data_wr_port_data[6]~28_combout ;
wire \M_dc_st_data[22]~25_combout ;
wire \A_dc_st_data[22]~q ;
wire \dc_data_wr_port_data[22]~29_combout ;
wire \M_dc_st_data[14]~26_combout ;
wire \A_dc_st_data[14]~q ;
wire \dc_data_wr_port_data[14]~30_combout ;
wire \M_dc_st_data[30]~27_combout ;
wire \A_dc_st_data[30]~q ;
wire \dc_data_wr_port_data[30]~31_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \i_readdata_d1[21]~q ;
wire \i_readdata_d1[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \i_readdata_d1[20]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \i_readdata_d1[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \i_readdata_d1[9]~q ;
wire \M_dc_st_data[3]~28_combout ;
wire \A_dc_st_data[3]~q ;
wire \dc_data_wr_port_data[3]~32_combout ;
wire \M_dc_st_data[19]~29_combout ;
wire \A_dc_st_data[19]~q ;
wire \dc_data_wr_port_data[19]~33_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \ic_tag_clr_valid_bits_nxt~combout ;
wire \ic_tag_wraddress_nxt~7_combout ;
wire \ic_tag_wraddress_nxt[0]~8_combout ;
wire \ic_tag_wraddress_nxt[1]~9_combout ;
wire \ic_tag_wraddress_nxt[1]~10_combout ;
wire \ic_tag_wraddress_nxt[2]~11_combout ;
wire \ic_tag_wraddress_nxt[3]~12_combout ;
wire \ic_tag_wraddress_nxt[4]~13_combout ;
wire \ic_tag_wraddress_nxt[5]~14_combout ;
wire \ic_tag_wraddress_nxt[6]~15_combout ;
wire \i_readdata_d1[7]~q ;
wire \M_dc_st_data[1]~30_combout ;
wire \A_dc_st_data[1]~q ;
wire \dc_data_wr_port_data[1]~34_combout ;
wire \M_dc_st_data[17]~31_combout ;
wire \A_dc_st_data[17]~q ;
wire \dc_data_wr_port_data[17]~35_combout ;
wire \the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \E_bht_data[0]~q ;
wire \E_br_mispredict~combout ;
wire \E_bht_ptr[0]~q ;
wire \E_bht_ptr[1]~q ;
wire \E_bht_ptr[2]~q ;
wire \E_bht_ptr[3]~q ;
wire \E_bht_ptr[4]~q ;
wire \E_bht_ptr[5]~q ;
wire \E_bht_ptr[6]~q ;
wire \E_bht_ptr[7]~q ;
wire \M_br_cond_taken_history[0]~0_combout ;
wire \ic_fill_valid_bits_nxt~0_combout ;
wire \ic_fill_valid_bits_en~combout ;
wire \ic_fill_valid_bits_nxt~1_combout ;
wire \ic_fill_valid_bits_nxt~2_combout ;
wire \ic_fill_valid_bits_nxt~3_combout ;
wire \D_bht_data[0]~q ;
wire \D_bht_ptr[0]~q ;
wire \D_bht_ptr[1]~q ;
wire \D_bht_ptr[2]~q ;
wire \D_bht_ptr[3]~q ;
wire \D_bht_ptr[4]~q ;
wire \D_bht_ptr[5]~q ;
wire \D_bht_ptr[6]~q ;
wire \D_bht_ptr[7]~q ;
wire \A_dc_rd_data[7]~q ;
wire \ic_fill_valid_bits_nxt~4_combout ;
wire \ic_fill_valid_bits_nxt~5_combout ;
wire \ic_fill_valid_bits_nxt~6_combout ;
wire \ic_fill_valid_bits_nxt~7_combout ;
wire \A_dc_rd_data[3]~q ;
wire \F_bht_ptr[0]~q ;
wire \F_bht_ptr[1]~q ;
wire \F_bht_ptr[2]~q ;
wire \F_bht_ptr[3]~q ;
wire \F_bht_ptr[4]~q ;
wire \F_bht_ptr[5]~q ;
wire \F_bht_ptr[6]~q ;
wire \F_bht_ptr[7]~q ;
wire \A_dc_rd_data[1]~q ;
wire \A_dc_rd_data[4]~q ;
wire \A_dc_rd_data[20]~q ;
wire \A_dc_rd_data[12]~q ;
wire \A_dc_rd_data[28]~q ;
wire \A_dc_rd_data[16]~q ;
wire \A_dc_rd_data[8]~q ;
wire \A_dc_rd_data[24]~q ;
wire \A_dc_rd_data[2]~q ;
wire \A_dc_rd_data[18]~q ;
wire \A_dc_rd_data[10]~q ;
wire \A_dc_rd_data[26]~q ;
wire \A_dc_rd_data[5]~q ;
wire \A_dc_rd_data[21]~q ;
wire \A_dc_rd_data[13]~q ;
wire \A_dc_rd_data[29]~q ;
wire \A_dc_rd_data[23]~q ;
wire \A_dc_rd_data[15]~q ;
wire \A_dc_rd_data[31]~q ;
wire \A_dc_rd_data[11]~q ;
wire \A_dc_rd_data[27]~q ;
wire \A_dc_rd_data[9]~q ;
wire \A_dc_rd_data[25]~q ;
wire \A_dc_rd_data[6]~q ;
wire \A_dc_rd_data[22]~q ;
wire \A_dc_rd_data[14]~q ;
wire \A_dc_rd_data[30]~q ;
wire \A_dc_rd_data[19]~q ;
wire \A_dc_rd_data[17]~q ;
wire \ic_tag_clr_valid_bits~0_combout ;
wire \M_br_mispredict~_wirecell_combout ;
wire \av_addr_accepted~combout ;
wire \F_iw[14]~10_combout ;
wire \F_iw[16]~6_combout ;
wire \D_iw[16]~q ;
wire \E_iw[16]~q ;
wire \F_iw[15]~7_combout ;
wire \D_iw[15]~q ;
wire \E_iw[15]~q ;
wire \F_iw[13]~8_combout ;
wire \D_iw[13]~q ;
wire \E_iw[13]~q ;
wire \E_hbreak_req~0_combout ;
wire \E_iw[5]~q ;
wire \F_iw[3]~2_combout ;
wire \D_iw[3]~q ;
wire \E_iw[3]~q ;
wire \F_iw[1]~3_combout ;
wire \D_iw[1]~q ;
wire \E_iw[1]~q ;
wire \F_iw[4]~4_combout ;
wire \D_iw[4]~q ;
wire \E_iw[4]~q ;
wire \F_iw[2]~5_combout ;
wire \D_iw[2]~q ;
wire \E_iw[2]~q ;
wire \Equal207~0_combout ;
wire \E_iw[14]~q ;
wire \F_iw[12]~11_combout ;
wire \D_iw[12]~q ;
wire \E_iw[12]~q ;
wire \F_iw[11]~12_combout ;
wire \D_iw[11]~q ;
wire \E_iw[11]~q ;
wire \E_hbreak_req~1_combout ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \E_valid~1_combout ;
wire \M_valid_from_E~q ;
wire \A_valid~q ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_div~0_combout ;
wire \E_ctrl_div~q ;
wire \M_ctrl_div~q ;
wire \A_ctrl_div~q ;
wire \A_div_do_sub~0_combout ;
wire \A_div_do_sub~q ;
wire \A_div_accumulate_quotient_bits~q ;
wire \A_div_discover_quotient_bits~0_combout ;
wire \F_iw[6]~28_combout ;
wire \D_iw[6]~q ;
wire \F_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~q ;
wire \F_iw[23]~14_combout ;
wire \D_iw[23]~q ;
wire \F_iw[18]~25_combout ;
wire \D_iw[18]~q ;
wire \F_ctrl_implicit_dst_retaddr~0_combout ;
wire \D_ctrl_implicit_dst_retaddr~q ;
wire \F_op_slli~2_combout ;
wire \F_op_slli~0_combout ;
wire \F_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~q ;
wire \D_dst_regnum[1]~0_combout ;
wire \F_iw[25]~17_combout ;
wire \D_iw[25]~q ;
wire \F_iw[20]~29_combout ;
wire \D_iw[20]~q ;
wire \D_dst_regnum[3]~3_combout ;
wire \F_ctrl_ignore_dst~combout ;
wire \D_ctrl_ignore_dst~q ;
wire \F_iw[22]~15_combout ;
wire \D_iw[22]~q ;
wire \F_iw[17]~26_combout ;
wire \D_iw[17]~q ;
wire \D_dst_regnum[0]~1_combout ;
wire \F_iw[24]~18_combout ;
wire \D_iw[24]~q ;
wire \F_iw[19]~30_combout ;
wire \D_iw[19]~q ;
wire \D_dst_regnum[2]~2_combout ;
wire \F_iw[26]~16_combout ;
wire \D_iw[26]~q ;
wire \F_iw[21]~27_combout ;
wire \D_iw[21]~q ;
wire \D_dst_regnum[4]~4_combout ;
wire \Equal297~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \D_regnum_b_cmp_F~0_combout ;
wire \D_regnum_b_cmp_F~1_combout ;
wire \D_regnum_b_cmp_F~combout ;
wire \E_regnum_b_cmp_D~q ;
wire \E_dst_regnum[2]~q ;
wire \E_hbreak_req~combout ;
wire \D_bht_data[1]~q ;
wire \E_bht_data[1]~q ;
wire \D_ctrl_cmp~3_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \E_ctrl_alu_subtract~q ;
wire \Equal152~1_combout ;
wire \Equal152~3_combout ;
wire \D_ctrl_alu_signed_comparison~0_combout ;
wire \D_ctrl_alu_signed_comparison~1_combout ;
wire \E_ctrl_alu_signed_comparison~q ;
wire \F_op_slli~3_combout ;
wire \F_op_slli~1_combout ;
wire \F_ctrl_src2_choose_imm~combout ;
wire \D_ctrl_src2_choose_imm~q ;
wire \Equal299~0_combout ;
wire \D_src2_reg[29]~2_combout ;
wire \D_src2_reg[0]~30_combout ;
wire \Equal90~0_combout ;
wire \D_ctrl_logic~1_combout ;
wire \D_ctrl_logic~2_combout ;
wire \E_ctrl_logic~q ;
wire \Equal103~0_combout ;
wire \Equal152~0_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \E_ctrl_retaddr~q ;
wire \D_ctrl_cmp~2_combout ;
wire \D_ctrl_cmp~0_combout ;
wire \D_ctrl_cmp~1_combout ;
wire \E_ctrl_cmp~q ;
wire \E_alu_result~0_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \Equal152~2_combout ;
wire \Equal152~4_combout ;
wire \Equal152~5_combout ;
wire \D_ctrl_alu_force_xor~0_combout ;
wire \D_ctrl_alu_force_xor~1_combout ;
wire \D_ctrl_alu_force_xor~2_combout ;
wire \D_logic_op[1]~0_combout ;
wire \E_logic_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \D_logic_op[0]~1_combout ;
wire \E_logic_op[0]~q ;
wire \E_alu_result~31_combout ;
wire \E_alu_result[31]~combout ;
wire \M_alu_result[31]~q ;
wire \D_ctrl_late_result~3_combout ;
wire \D_ctrl_mul_lsw~0_combout ;
wire \E_ctrl_mul_lsw~q ;
wire \M_ctrl_mul_lsw~q ;
wire \A_ctrl_mul_lsw~q ;
wire \E_op_rdctl~0_combout ;
wire \E_op_rdctl~combout ;
wire \M_ctrl_rdctl_inst~q ;
wire \M_ctrl_mem_nxt~0_combout ;
wire \M_ctrl_mem~q ;
wire \A_inst_result[31]~q ;
wire \D_ctrl_shift_rot~0_combout ;
wire \E_ctrl_shift_rot~q ;
wire \M_ctrl_shift_rot~q ;
wire \A_ctrl_shift_rot~q ;
wire \E_dst_regnum[4]~q ;
wire \M_dst_regnum[4]~q ;
wire \M_wr_dst_reg_from_E~q ;
wire \E_dst_regnum[0]~q ;
wire \M_dst_regnum[0]~q ;
wire \E_dst_regnum[1]~q ;
wire \M_dst_regnum[1]~q ;
wire \M_regnum_b_cmp_F~0_combout ;
wire \M_dst_regnum[2]~q ;
wire \E_dst_regnum[3]~q ;
wire \M_dst_regnum[3]~q ;
wire \M_regnum_b_cmp_F~1_combout ;
wire \M_regnum_b_cmp_F~combout ;
wire \A_regnum_b_cmp_D~q ;
wire \A_dst_regnum_from_M[4]~q ;
wire \A_wr_dst_reg_from_M~q ;
wire \A_dst_regnum_from_M[0]~q ;
wire \A_dst_regnum_from_M[1]~q ;
wire \A_regnum_b_cmp_F~0_combout ;
wire \A_dst_regnum_from_M[2]~q ;
wire \A_dst_regnum_from_M[3]~q ;
wire \A_regnum_b_cmp_F~1_combout ;
wire \A_regnum_b_cmp_F~combout ;
wire \W_regnum_b_cmp_D~q ;
wire \D_src2_reg[29]~4_combout ;
wire \D_src2_reg[29]~3_combout ;
wire \D_src2_reg[3]~13_combout ;
wire \A_mul_partial_prod[15]~q ;
wire \A_mul_partial_prod[14]~q ;
wire \A_mul_partial_prod[13]~q ;
wire \A_mul_partial_prod[12]~q ;
wire \A_mul_partial_prod[11]~q ;
wire \A_mul_partial_prod[10]~q ;
wire \A_mul_partial_prod[9]~q ;
wire \A_mul_partial_prod[8]~q ;
wire \A_mul_partial_prod[7]~q ;
wire \A_mul_partial_prod[6]~q ;
wire \A_mul_partial_prod[5]~q ;
wire \A_mul_partial_prod[4]~q ;
wire \A_mul_partial_prod[3]~q ;
wire \A_mul_partial_prod[2]~q ;
wire \A_mul_partial_prod[1]~q ;
wire \A_mul_partial_prod[0]~q ;
wire \Add26~5_sumout ;
wire \E_ld_st_dcache_management_bus~0_combout ;
wire \M_ctrl_ld_st_bypass_or_dcache_management~q ;
wire \A_mem_stall_nxt~0_combout ;
wire \E_st_bus~0_combout ;
wire \M_ctrl_st_bypass~q ;
wire \A_inst_result[16]~q ;
wire \A_mul_partial_prod[16]~q ;
wire \Add26~50 ;
wire \Add26~45_sumout ;
wire \A_mul_result[16]~q ;
wire \F_iw[7]~32_combout ;
wire \D_iw[7]~q ;
wire \d_readdata_d1[1]~q ;
wire \d_readdata_d1[17]~q ;
wire \d_readdata_d1[9]~q ;
wire \d_readdata_d1[25]~q ;
wire \E_ctrl_ld8_ld16~0_combout ;
wire \Equal182~0_combout ;
wire \M_ctrl_ld8~q ;
wire \Equal185~0_combout ;
wire \M_ctrl_ld16~q ;
wire \M_ld_align_sh16~0_combout ;
wire \A_ld_align_sh16~q ;
wire \E_compare_op[0]~q ;
wire \D_src2_reg[0]~31_combout ;
wire \E_alu_result~17_combout ;
wire \E_alu_result[29]~combout ;
wire \M_alu_result[29]~q ;
wire \A_inst_result[29]~q ;
wire \A_mul_partial_prod[29]~q ;
wire \A_mul_partial_prod[28]~q ;
wire \A_mul_partial_prod[27]~q ;
wire \A_mul_partial_prod[26]~q ;
wire \A_mul_partial_prod[25]~q ;
wire \A_mul_partial_prod[24]~q ;
wire \A_mul_partial_prod[23]~q ;
wire \A_mul_partial_prod[22]~q ;
wire \A_mul_partial_prod[21]~q ;
wire \A_mul_partial_prod[20]~q ;
wire \A_mul_partial_prod[19]~q ;
wire \A_mul_partial_prod[18]~q ;
wire \A_mul_partial_prod[17]~q ;
wire \Add26~46 ;
wire \Add26~97_sumout ;
wire \A_mul_result[17]~q ;
wire \Add26~98 ;
wire \Add26~113_sumout ;
wire \A_mul_result[18]~q ;
wire \Add26~114 ;
wire \Add26~89_sumout ;
wire \A_mul_result[19]~q ;
wire \Add26~90 ;
wire \Add26~109_sumout ;
wire \A_mul_result[20]~q ;
wire \Add26~110 ;
wire \Add26~105_sumout ;
wire \A_mul_result[21]~q ;
wire \Add26~106 ;
wire \Add26~101_sumout ;
wire \A_mul_result[22]~q ;
wire \Add26~102 ;
wire \Add26~121_sumout ;
wire \A_mul_result[23]~q ;
wire \Add26~122 ;
wire \Add26~117_sumout ;
wire \A_mul_result[24]~q ;
wire \Add26~118 ;
wire \Add26~85_sumout ;
wire \A_mul_result[25]~q ;
wire \Add26~86 ;
wire \Add26~81_sumout ;
wire \A_mul_result[26]~q ;
wire \Add26~82 ;
wire \Add26~73_sumout ;
wire \A_mul_result[27]~q ;
wire \Add26~74 ;
wire \Add26~69_sumout ;
wire \A_mul_result[28]~q ;
wire \Add26~70 ;
wire \Add26~65_sumout ;
wire \A_mul_result[29]~q ;
wire \E_ctrl_ld_signed~0_combout ;
wire \M_ctrl_ld_signed~q ;
wire \A_ctrl_ld_signed~q ;
wire \D_ctrl_shift_right_arith~0_combout ;
wire \E_ctrl_shift_right_arith~q ;
wire \E_rot_fill_bit~0_combout ;
wire \M_rot_fill_bit~q ;
wire \F_iw[8]~24_combout ;
wire \D_iw[8]~q ;
wire \d_readdata_d1[2]~q ;
wire \d_readdata_d1[18]~q ;
wire \d_readdata_d1[10]~q ;
wire \d_readdata_d1[26]~q ;
wire \A_slow_inst_result_nxt[2]~2_combout ;
wire \Equal152~6_combout ;
wire \E_ctrl_div_signed_nxt~combout ;
wire \E_ctrl_div_signed~q ;
wire \E_div_negate_src2~0_combout ;
wire \E_div_negate_src1~0_combout ;
wire \E_div_negate_result~combout ;
wire \M_div_negate_result~q ;
wire \A_div_negate_result~q ;
wire \A_div_quot_bit~0_combout ;
wire \A_div_quot_bit~q ;
wire \Add14~5_sumout ;
wire \A_div_quot_en~combout ;
wire \A_div_quot[0]~q ;
wire \Add14~6 ;
wire \Add14~93_sumout ;
wire \A_div_quot[1]~q ;
wire \Add14~94 ;
wire \Add14~9_sumout ;
wire \A_div_quot[2]~q ;
wire \d_readdatavalid_d1~q ;
wire \E_ld_bus~0_combout ;
wire \M_ctrl_ld_bypass~q ;
wire \A_ctrl_ld_bypass~q ;
wire \F_iw[10]~13_combout ;
wire \D_iw[10]~q ;
wire \d_readdata_d1[4]~q ;
wire \d_readdata_d1[20]~q ;
wire \d_readdata_d1[12]~q ;
wire \d_readdata_d1[28]~q ;
wire \A_slow_inst_result_nxt[4]~0_combout ;
wire \Add14~10 ;
wire \Add14~61_sumout ;
wire \A_div_quot[3]~q ;
wire \Add14~62 ;
wire \Add14~1_sumout ;
wire \A_div_quot[4]~q ;
wire \A_slow_inst_result[4]~q ;
wire \A_inst_result[4]~q ;
wire \F_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~q ;
wire \F_ctrl_unsigned_lo_imm16~1_combout ;
wire \F_ctrl_unsigned_lo_imm16~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~q ;
wire \Equal300~0_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \E_ctrl_shift_rot_right~q ;
wire \E_rot_mask[4]~0_combout ;
wire \M_rot_mask[4]~q ;
wire \F_iw[9]~31_combout ;
wire \D_iw[9]~q ;
wire \d_readdata_d1[3]~q ;
wire \d_readdata_d1[19]~q ;
wire \d_readdata_d1[11]~q ;
wire \d_readdata_d1[27]~q ;
wire \A_slow_inst_result_nxt[3]~15_combout ;
wire \A_slow_inst_result[3]~q ;
wire \A_inst_result[3]~q ;
wire \E_rot_mask[3]~4_combout ;
wire \M_rot_mask[3]~q ;
wire \D_ctrl_shift_rot_left~0_combout ;
wire \E_ctrl_shift_rot_left~q ;
wire \E_rot_sel_fill2~0_combout ;
wire \M_rot_sel_fill2~q ;
wire \F_ctrl_a_not_src~0_combout ;
wire \D_ctrl_a_not_src~q ;
wire \E_regnum_a_cmp_F~0_combout ;
wire \E_regnum_a_cmp_F~1_combout ;
wire \E_regnum_a_cmp_F~combout ;
wire \D_regnum_a_cmp_F~0_combout ;
wire \D_regnum_a_cmp_F~1_combout ;
wire \D_regnum_a_cmp_F~combout ;
wire \E_regnum_a_cmp_D~q ;
wire \M_regnum_a_cmp_D~q ;
wire \A_regnum_a_cmp_F~0_combout ;
wire \A_regnum_a_cmp_F~1_combout ;
wire \A_regnum_a_cmp_F~combout ;
wire \M_regnum_a_cmp_F~0_combout ;
wire \M_regnum_a_cmp_F~1_combout ;
wire \M_regnum_a_cmp_F~combout ;
wire \A_regnum_a_cmp_D~q ;
wire \W_regnum_a_cmp_D~q ;
wire \E_src1[3]~0_combout ;
wire \E_src1[3]~1_combout ;
wire \D_src1_reg[15]~11_combout ;
wire \F_iw[31]~19_combout ;
wire \D_iw[31]~q ;
wire \F_iw[30]~20_combout ;
wire \D_iw[30]~q ;
wire \F_iw[29]~21_combout ;
wire \D_iw[29]~q ;
wire \F_iw[27]~22_combout ;
wire \D_iw[27]~q ;
wire \F_iw[28]~23_combout ;
wire \D_iw[28]~q ;
wire \Equal298~0_combout ;
wire \D_src1_hazard_E~combout ;
wire \E_src1[15]~q ;
wire \D_ctrl_rot~0_combout ;
wire \E_ctrl_rot~q ;
wire \E_rot_pass1~0_combout ;
wire \M_rot_pass1~q ;
wire \E_rot_sel_fill1~0_combout ;
wire \M_rot_sel_fill1~q ;
wire \E_rot_mask[6]~7_combout ;
wire \M_rot_mask[6]~q ;
wire \E_rot_mask[2]~2_combout ;
wire \M_rot_mask[2]~q ;
wire \d_readdata_d1[6]~q ;
wire \d_readdata_d1[22]~q ;
wire \d_readdata_d1[14]~q ;
wire \d_readdata_d1[30]~q ;
wire \A_slow_inst_result_nxt[6]~10_combout ;
wire \Add14~2 ;
wire \Add14~13_sumout ;
wire \A_div_quot[5]~q ;
wire \Add14~14 ;
wire \Add14~41_sumout ;
wire \A_div_quot[6]~q ;
wire \A_slow_inst_result[6]~q ;
wire \A_inst_result[6]~q ;
wire \A_inst_result[18]~q ;
wire \E_rot_mask[1]~5_combout ;
wire \M_rot_mask[1]~q ;
wire \d_readdata_d1[5]~q ;
wire \d_readdata_d1[21]~q ;
wire \d_readdata_d1[13]~q ;
wire \d_readdata_d1[29]~q ;
wire \A_slow_inst_result_nxt[5]~3_combout ;
wire \A_slow_inst_result[5]~q ;
wire \A_inst_result[5]~q ;
wire \A_inst_result[17]~q ;
wire \E_rot_mask[0]~1_combout ;
wire \M_rot_mask[0]~q ;
wire \D_src1_reg[4]~0_combout ;
wire \E_src1[4]~q ;
wire \D_src1_reg[1]~23_combout ;
wire \E_src1[1]~q ;
wire \Add7~0_combout ;
wire \E_rot_step1[4]~1_combout ;
wire \Add7~1_combout ;
wire \M_rot_prestep2[8]~q ;
wire \D_src1_reg[20]~27_combout ;
wire \E_src1[20]~q ;
wire \D_src1_reg[19]~22_combout ;
wire \E_src1[19]~q ;
wire \D_src1_reg[16]~10_combout ;
wire \E_src1[16]~q ;
wire \d_readdata_d1[7]~q ;
wire \d_readdata_d1[23]~q ;
wire \d_readdata_d1[15]~q ;
wire \d_readdata_d1[31]~q ;
wire \A_slow_inst_result_nxt[7]~9_combout ;
wire \Add14~42 ;
wire \Add14~37_sumout ;
wire \A_div_quot[7]~q ;
wire \A_slow_inst_result[7]~q ;
wire \A_inst_result[7]~q ;
wire \A_inst_result[23]~q ;
wire \A_inst_result[15]~q ;
wire \A_wr_data_unfiltered[7]~22_combout ;
wire \E_rot_pass0~0_combout ;
wire \M_rot_pass0~q ;
wire \E_rot_sel_fill0~0_combout ;
wire \M_rot_sel_fill0~q ;
wire \E_rot_mask[7]~6_combout ;
wire \M_rot_mask[7]~q ;
wire \d_readdata_d1[0]~q ;
wire \d_readdata_d1[16]~q ;
wire \d_readdata_d1[8]~q ;
wire \d_readdata_d1[24]~q ;
wire \A_slow_inst_result_nxt[0]~1_combout ;
wire \A_slow_inst_result[0]~q ;
wire \M_inst_result[0]~0_combout ;
wire \A_div_stall~0_combout ;
wire \E_iw[6]~q ;
wire \M_iw[6]~q ;
wire \E_iw[7]~q ;
wire \M_iw[7]~q ;
wire \E_iw[8]~q ;
wire \M_iw[8]~q ;
wire \E_op_wrctl~combout ;
wire \M_ctrl_wrctl_inst~q ;
wire \A_ienable_reg_irq0_nxt~0_combout ;
wire \A_ienable_reg_irq0~0_combout ;
wire \A_ienable_reg_irq0~q ;
wire \A_ipending_reg_irq0_nxt~0_combout ;
wire \A_ipending_reg_irq0~q ;
wire \D_ctrl_exception~0_combout ;
wire \E_ctrl_exception~q ;
wire \M_ctrl_exception~q ;
wire \D_ctrl_crst~0_combout ;
wire \E_ctrl_crst~q ;
wire \M_ctrl_crst~q ;
wire \M_wrctl_estatus~combout ;
wire \A_estatus_reg_pie_inst_nxt~0_combout ;
wire \A_estatus_reg_pie~q ;
wire \M_wrctl_bstatus~combout ;
wire \A_bstatus_reg_pie_inst_nxt~0_combout ;
wire \A_bstatus_reg_pie~q ;
wire \D_control_reg_rddata_muxed[0]~0_combout ;
wire \D_control_reg_rddata_muxed[0]~1_combout ;
wire \E_control_reg_rddata[0]~q ;
wire \M_control_reg_rddata[0]~q ;
wire \A_inst_result[0]~q ;
wire \A_inst_result[8]~q ;
wire \A_inst_result[24]~q ;
wire \A_wr_data_unfiltered[0]~4_combout ;
wire \E_rot_step1[20]~5_combout ;
wire \E_rot_step1[24]~2_combout ;
wire \M_rot_prestep2[24]~q ;
wire \E_rot_step1[12]~7_combout ;
wire \E_rot_step1[16]~4_combout ;
wire \M_rot_prestep2[16]~q ;
wire \Add7~2_combout ;
wire \M_rot_rn[3]~q ;
wire \Add7~3_combout ;
wire \M_rot_rn[4]~q ;
wire \M_rot[0]~1_combout ;
wire \A_shift_rot_result~1_combout ;
wire \A_shift_rot_result[0]~q ;
wire \A_wr_data_unfiltered[6]~1_combout ;
wire \A_wr_data_unfiltered[6]~2_combout ;
wire \A_wr_data_unfiltered[0]~5_combout ;
wire \W_wr_data[0]~q ;
wire \D_src1_reg[0]~21_combout ;
wire \E_src1[0]~q ;
wire \E_rot_step1[3]~27_combout ;
wire \M_rot_prestep2[7]~q ;
wire \E_rot_step1[27]~29_combout ;
wire \E_logic_result[30]~12_combout ;
wire \E_alu_result~20_combout ;
wire \D_src2_reg[30]~38_combout ;
wire \A_inst_result[30]~q ;
wire \A_mul_partial_prod[30]~q ;
wire \Add26~66 ;
wire \Add26~77_sumout ;
wire \A_mul_result[30]~q ;
wire \E_rot_pass3~0_combout ;
wire \M_rot_pass3~q ;
wire \E_rot_sel_fill3~0_combout ;
wire \M_rot_sel_fill3~q ;
wire \E_rot_step1[26]~11_combout ;
wire \E_rot_step1[30]~8_combout ;
wire \M_rot_prestep2[30]~q ;
wire \E_rot_step1[2]~9_combout ;
wire \M_rot_prestep2[6]~q ;
wire \M_rot[6]~19_combout ;
wire \A_shift_rot_result~19_combout ;
wire \A_shift_rot_result[30]~q ;
wire \M_ctrl_ld8_ld16~q ;
wire \A_ld_align_byte2_byte3_fill~q ;
wire \A_mem_baddr[1]~q ;
wire \A_mem_baddr[0]~q ;
wire \A_ctrl_ld16~q ;
wire \A_slow_ld_data_sign_bit~0_combout ;
wire \A_slow_ld_data_fill_bit~0_combout ;
wire \A_slow_inst_result_nxt[30]~19_combout ;
wire \Add14~38 ;
wire \Add14~33_sumout ;
wire \A_div_quot[8]~q ;
wire \Add14~34 ;
wire \Add14~29_sumout ;
wire \A_div_quot[9]~q ;
wire \Add14~30 ;
wire \Add14~25_sumout ;
wire \A_div_quot[10]~q ;
wire \Add14~26 ;
wire \Add14~21_sumout ;
wire \A_div_quot[11]~q ;
wire \Add14~22 ;
wire \Add14~17_sumout ;
wire \A_div_quot[12]~q ;
wire \Add14~18 ;
wire \Add14~57_sumout ;
wire \A_div_quot[13]~q ;
wire \Add14~58 ;
wire \Add14~53_sumout ;
wire \A_div_quot[14]~q ;
wire \Add14~54 ;
wire \Add14~49_sumout ;
wire \A_div_quot[15]~q ;
wire \Add14~50 ;
wire \Add14~45_sumout ;
wire \A_div_quot[16]~q ;
wire \Add14~46 ;
wire \Add14~97_sumout ;
wire \A_div_quot[17]~q ;
wire \Add14~98 ;
wire \Add14~113_sumout ;
wire \A_div_quot[18]~q ;
wire \Add14~114 ;
wire \Add14~89_sumout ;
wire \A_div_quot[19]~q ;
wire \Add14~90 ;
wire \Add14~109_sumout ;
wire \A_div_quot[20]~q ;
wire \Add14~110 ;
wire \Add14~105_sumout ;
wire \A_div_quot[21]~q ;
wire \Add14~106 ;
wire \Add14~101_sumout ;
wire \A_div_quot[22]~q ;
wire \Add14~102 ;
wire \Add14~121_sumout ;
wire \A_div_quot[23]~q ;
wire \Add14~122 ;
wire \Add14~117_sumout ;
wire \A_div_quot[24]~q ;
wire \Add14~118 ;
wire \Add14~85_sumout ;
wire \A_div_quot[25]~q ;
wire \Add14~86 ;
wire \Add14~81_sumout ;
wire \A_div_quot[26]~q ;
wire \Add14~82 ;
wire \Add14~73_sumout ;
wire \A_div_quot[27]~q ;
wire \Add14~74 ;
wire \Add14~69_sumout ;
wire \A_div_quot[28]~q ;
wire \Add14~70 ;
wire \Add14~65_sumout ;
wire \A_div_quot[29]~q ;
wire \Add14~66 ;
wire \Add14~77_sumout ;
wire \A_div_quot[30]~q ;
wire \A_slow_inst_result[30]~q ;
wire \A_wr_data_unfiltered[30]~43_combout ;
wire \A_wr_data_unfiltered[30]~44_combout ;
wire \W_wr_data[30]~q ;
wire \D_src2_reg[30]~39_combout ;
wire \D_src2[30]~8_combout ;
wire \D_src2[30]~9_combout ;
wire \E_src2[18]~1_combout ;
wire \E_src2[30]~q ;
wire \Add24~86 ;
wire \Add24~82 ;
wire \Add24~77_sumout ;
wire \E_alu_result[30]~combout ;
wire \M_alu_result[30]~q ;
wire \D_src1_reg[30]~18_combout ;
wire \E_src1[30]~q ;
wire \E_rot_step1[31]~26_combout ;
wire \M_rot_prestep2[31]~q ;
wire \E_rot_step1[19]~31_combout ;
wire \E_rot_step1[23]~28_combout ;
wire \M_rot_prestep2[23]~q ;
wire \E_rot_step1[11]~25_combout ;
wire \M_rot_prestep2[15]~q ;
wire \M_rot[7]~9_combout ;
wire \A_shift_rot_result~9_combout ;
wire \A_shift_rot_result[7]~q ;
wire \A_wr_data_unfiltered[7]~23_combout ;
wire \W_wr_data[7]~q ;
wire \D_src2_reg[7]~19_combout ;
wire \D_src2_reg[7]~20_combout ;
wire \E_src2[0]~0_combout ;
wire \E_src2[7]~q ;
wire \Add24~134_cout ;
wire \Add24~74 ;
wire \Add24~70 ;
wire \Add24~26 ;
wire \Add24~30 ;
wire \Add24~34 ;
wire \Add24~18 ;
wire \Add24~22 ;
wire \Add24~9_sumout ;
wire \E_alu_result~9_combout ;
wire \E_ctrl_jmp_indirect_nxt~0_combout ;
wire \E_valid_jmp_indirect~0_combout ;
wire \E_valid_jmp_indirect~q ;
wire \E_ctrl_jmp_indirect~q ;
wire \M_pipe_flush_waddr[0]~0_combout ;
wire \M_pipe_flush_waddr[0]~1_combout ;
wire \M_pipe_flush_waddr_nxt[5]~5_combout ;
wire \D_pc[5]~q ;
wire \E_pc[5]~q ;
wire \M_pipe_flush_waddr[0]~2_combout ;
wire \M_pipe_flush_waddr[5]~q ;
wire \D_pc[12]~q ;
wire \D_pc[11]~q ;
wire \D_pc[10]~q ;
wire \Add3~5_sumout ;
wire \Add0~5_sumout ;
wire \D_br_taken_waddr_partial[0]~q ;
wire \D_pc_plus_one[0]~q ;
wire \E_ctrl_br_cond_nxt~0_combout ;
wire \D_br_pred_not_taken~combout ;
wire \E_extra_pc[0]~q ;
wire \M_pipe_flush_waddr_nxt[0]~11_combout ;
wire \D_pc[0]~q ;
wire \E_pc[0]~q ;
wire \M_pipe_flush_waddr[0]~q ;
wire \F_ic_valid~4_combout ;
wire \F_ic_valid~0_combout ;
wire \F_ic_hit~0_combout ;
wire \D_pc[14]~q ;
wire \D_pc[13]~q ;
wire \Add3~50 ;
wire \Add3~45_sumout ;
wire \D_pc_plus_one[13]~q ;
wire \Add0~6 ;
wire \Add0~38 ;
wire \Add0~2 ;
wire \Add0~10 ;
wire \Add0~34 ;
wire \Add0~30 ;
wire \Add0~26 ;
wire \Add0~22 ;
wire \Add0~18 ;
wire \Add0~14 ;
wire \Add0~41_sumout ;
wire \D_br_taken_waddr_partial[10]~q ;
wire \Add1~22_cout ;
wire \Add1~2 ;
wire \Add1~18 ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \F_pc_nxt~8_combout ;
wire \F_pc_nxt~9_combout ;
wire \E_extra_pc[13]~q ;
wire \M_pipe_flush_waddr_nxt[13]~10_combout ;
wire \E_pc[13]~q ;
wire \M_pipe_flush_waddr[13]~q ;
wire \F_pc[13]~q ;
wire \Add3~46 ;
wire \Add3~41_sumout ;
wire \D_pc_plus_one[14]~q ;
wire \Add1~10 ;
wire \Add1~5_sumout ;
wire \F_pc_nxt~6_combout ;
wire \F_pc_nxt~7_combout ;
wire \M_pipe_flush_waddr[12]~3_combout ;
wire \E_extra_pc[14]~q ;
wire \E_pc[14]~q ;
wire \M_pipe_flush_waddr_nxt[14]~14_combout ;
wire \M_pipe_flush_waddr[14]~5_combout ;
wire \M_pipe_flush_waddr[14]~q ;
wire \M_pipe_flush_waddr[14]~_wirecell_combout ;
wire \F_pc[14]~q ;
wire \F_ic_hit~1_combout ;
wire \F_issue~combout ;
wire \D_issue~q ;
wire \F_ctrl_br~0_combout ;
wire \D_ctrl_br~q ;
wire \F_ctrl_br_uncond~0_combout ;
wire \D_ctrl_br_uncond~q ;
wire \D_br_pred_taken~0_combout ;
wire \F_kill~2_combout ;
wire \F_kill~0_combout ;
wire \F_kill~1_combout ;
wire \D_kill~q ;
wire \F_pc[14]~1_combout ;
wire \F_ic_data_rd_addr_nxt[0]~0_combout ;
wire \F_ic_data_rd_addr_nxt[0]~1_combout ;
wire \F_pc[0]~q ;
wire \Add3~6 ;
wire \Add3~57_sumout ;
wire \Add0~37_sumout ;
wire \D_br_taken_waddr_partial[1]~q ;
wire \D_pc_plus_one[1]~q ;
wire \E_extra_pc[1]~q ;
wire \M_pipe_flush_waddr_nxt[1]~12_combout ;
wire \D_pc[1]~q ;
wire \E_pc[1]~q ;
wire \M_pipe_flush_waddr[1]~q ;
wire \F_ic_data_rd_addr_nxt[1]~2_combout ;
wire \F_ic_data_rd_addr_nxt[1]~3_combout ;
wire \F_pc[1]~q ;
wire \Add3~58 ;
wire \Add3~1_sumout ;
wire \Add0~1_sumout ;
wire \D_br_taken_waddr_partial[2]~q ;
wire \D_pc_plus_one[2]~q ;
wire \E_extra_pc[2]~q ;
wire \M_pipe_flush_waddr_nxt[2]~13_combout ;
wire \D_pc[2]~q ;
wire \E_pc[2]~q ;
wire \M_pipe_flush_waddr[2]~q ;
wire \F_ic_data_rd_addr_nxt[2]~4_combout ;
wire \F_ic_data_rd_addr_nxt[2]~5_combout ;
wire \F_pc[2]~q ;
wire \Add3~2 ;
wire \Add3~9_sumout ;
wire \Add0~9_sumout ;
wire \D_br_taken_waddr_partial[3]~q ;
wire \D_pc_plus_one[3]~q ;
wire \E_extra_pc[3]~q ;
wire \M_pipe_flush_waddr_nxt[3]~7_combout ;
wire \D_pc[3]~q ;
wire \E_pc[3]~q ;
wire \M_pipe_flush_waddr[3]~q ;
wire \F_ic_tag_rd_addr_nxt[0]~12_combout ;
wire \F_ic_tag_rd_addr_nxt[0]~13_combout ;
wire \F_pc[3]~q ;
wire \Add3~10 ;
wire \Add3~37_sumout ;
wire \Add0~33_sumout ;
wire \D_br_taken_waddr_partial[4]~q ;
wire \D_pc_plus_one[4]~q ;
wire \E_extra_pc[4]~q ;
wire \M_pipe_flush_waddr_nxt[4]~4_combout ;
wire \D_pc[4]~q ;
wire \E_pc[4]~q ;
wire \M_pipe_flush_waddr[4]~q ;
wire \F_ic_tag_rd_addr_nxt[1]~8_combout ;
wire \F_ic_tag_rd_addr_nxt[1]~9_combout ;
wire \F_pc[4]~q ;
wire \Add3~38 ;
wire \Add3~34 ;
wire \Add3~29_sumout ;
wire \Add0~25_sumout ;
wire \D_br_taken_waddr_partial[6]~q ;
wire \D_pc_plus_one[6]~q ;
wire \E_extra_pc[6]~q ;
wire \M_pipe_flush_waddr_nxt[6]~3_combout ;
wire \D_pc[6]~q ;
wire \E_pc[6]~q ;
wire \M_pipe_flush_waddr[6]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~6_combout ;
wire \F_ic_tag_rd_addr_nxt[3]~7_combout ;
wire \F_pc[6]~q ;
wire \Add3~30 ;
wire \Add3~25_sumout ;
wire \Add0~21_sumout ;
wire \D_br_taken_waddr_partial[7]~q ;
wire \D_pc_plus_one[7]~q ;
wire \E_extra_pc[7]~q ;
wire \M_pipe_flush_waddr_nxt[7]~1_combout ;
wire \D_pc[7]~q ;
wire \E_pc[7]~q ;
wire \M_pipe_flush_waddr[7]~q ;
wire \F_ic_tag_rd_addr_nxt[4]~2_combout ;
wire \F_ic_tag_rd_addr_nxt[4]~3_combout ;
wire \F_pc[7]~q ;
wire \Add3~26 ;
wire \Add3~21_sumout ;
wire \Add0~17_sumout ;
wire \D_br_taken_waddr_partial[8]~q ;
wire \D_pc_plus_one[8]~q ;
wire \E_extra_pc[8]~q ;
wire \M_pipe_flush_waddr_nxt[8]~2_combout ;
wire \D_pc[8]~q ;
wire \E_pc[8]~q ;
wire \M_pipe_flush_waddr[8]~q ;
wire \F_ic_tag_rd_addr_nxt[5]~4_combout ;
wire \F_ic_tag_rd_addr_nxt[5]~5_combout ;
wire \F_pc[8]~q ;
wire \Add3~22 ;
wire \Add3~17_sumout ;
wire \Add0~13_sumout ;
wire \D_br_taken_waddr_partial[9]~q ;
wire \D_pc_plus_one[9]~q ;
wire \E_extra_pc[9]~q ;
wire \M_pipe_flush_waddr_nxt[9]~0_combout ;
wire \D_pc[9]~q ;
wire \E_pc[9]~q ;
wire \M_pipe_flush_waddr[9]~q ;
wire \F_ic_tag_rd_addr_nxt[6]~0_combout ;
wire \F_ic_tag_rd_addr_nxt[6]~1_combout ;
wire \F_pc[9]~q ;
wire \Add3~18 ;
wire \Add3~13_sumout ;
wire \D_pc_plus_one[10]~q ;
wire \Add1~1_sumout ;
wire \F_pc_nxt~2_combout ;
wire \F_pc_nxt~3_combout ;
wire \E_extra_pc[10]~q ;
wire \M_pipe_flush_waddr_nxt[10]~8_combout ;
wire \E_pc[10]~q ;
wire \M_pipe_flush_waddr[10]~q ;
wire \F_pc[10]~q ;
wire \Add3~14 ;
wire \Add3~53_sumout ;
wire \D_pc_plus_one[11]~q ;
wire \Add1~17_sumout ;
wire \F_pc_nxt~4_combout ;
wire \F_pc_nxt~5_combout ;
wire \E_extra_pc[11]~q ;
wire \M_pipe_flush_waddr_nxt[11]~9_combout ;
wire \E_pc[11]~q ;
wire \M_pipe_flush_waddr[11]~q ;
wire \F_pc[11]~q ;
wire \Add3~54 ;
wire \Add3~49_sumout ;
wire \D_pc_plus_one[12]~q ;
wire \Add1~13_sumout ;
wire \F_pc_nxt~0_combout ;
wire \F_pc_nxt~1_combout ;
wire \E_pc[12]~q ;
wire \E_extra_pc[12]~q ;
wire \M_pipe_flush_waddr_nxt[12]~6_combout ;
wire \M_pipe_flush_waddr[12]~q ;
wire \M_pipe_flush_waddr[12]~_wirecell_combout ;
wire \F_pc[12]~q ;
wire \F_ic_hit~2_combout ;
wire \D_iw_valid~q ;
wire \F_pc[14]~0_combout ;
wire \F_ic_tag_rd_addr_nxt[2]~10_combout ;
wire \F_ic_tag_rd_addr_nxt[2]~11_combout ;
wire \F_pc[5]~q ;
wire \Add3~33_sumout ;
wire \Add0~29_sumout ;
wire \D_br_taken_waddr_partial[5]~q ;
wire \D_pc_plus_one[5]~q ;
wire \E_extra_pc[5]~q ;
wire \E_alu_result[7]~combout ;
wire \M_alu_result[7]~q ;
wire \D_src1_reg[7]~8_combout ;
wire \E_src1[7]~q ;
wire \E_rot_step1[7]~24_combout ;
wire \M_rot_prestep2[11]~q ;
wire \M_rot_prestep2[3]~q ;
wire \M_rot_prestep2[27]~q ;
wire \M_rot[3]~5_combout ;
wire \A_shift_rot_result~5_combout ;
wire \A_shift_rot_result[11]~q ;
wire \A_inst_result[11]~q ;
wire \A_inst_result[27]~q ;
wire \A_ld_align_byte1_fill~q ;
wire \A_slow_inst_result[15]~0_combout ;
wire \A_slow_inst_result[15]~1_combout ;
wire \A_slow_inst_result_nxt[11]~5_combout ;
wire \A_slow_inst_result[11]~q ;
wire \A_data_ram_ld_align_fill_bit~combout ;
wire \A_wr_data_unfiltered[8]~10_combout ;
wire \A_wr_data_unfiltered[8]~11_combout ;
wire \A_wr_data_unfiltered[11]~14_combout ;
wire \A_wr_data_unfiltered[11]~15_combout ;
wire \W_wr_data[11]~q ;
wire \D_src1_reg[11]~4_combout ;
wire \E_src1[11]~q ;
wire \Add24~10 ;
wire \Add24~2 ;
wire \Add24~6 ;
wire \Add24~14 ;
wire \Add24~45_sumout ;
wire \E_logic_result[11]~1_combout ;
wire \E_alu_result[11]~5_combout ;
wire \E_alu_result[11]~combout ;
wire \M_alu_result[11]~q ;
wire \D_src2_reg[11]~15_combout ;
wire \D_src2_reg[11]~92_combout ;
wire \D_src2_reg[11]~123_combout ;
wire \E_src2[11]~q ;
wire \Add24~46 ;
wire \Add24~42 ;
wire \Add24~62 ;
wire \Add24~58 ;
wire \Add24~54 ;
wire \Add24~50 ;
wire \Add24~106 ;
wire \Add24~122 ;
wire \Add24~102 ;
wire \Add24~118 ;
wire \Add24~114 ;
wire \Add24~110 ;
wire \Add24~129_sumout ;
wire \E_alu_result[23]~combout ;
wire \M_alu_result[23]~q ;
wire \M_rot[7]~30_combout ;
wire \A_shift_rot_result~30_combout ;
wire \A_shift_rot_result[23]~q ;
wire \A_slow_inst_result_nxt[23]~30_combout ;
wire \A_slow_inst_result[23]~q ;
wire \A_wr_data_unfiltered[23]~65_combout ;
wire \A_wr_data_unfiltered[23]~66_combout ;
wire \W_wr_data[23]~q ;
wire \D_src1_reg[23]~30_combout ;
wire \E_src1[23]~q ;
wire \E_alu_result~30_combout ;
wire \D_src2_reg[23]~58_combout ;
wire \D_src2_reg[23]~59_combout ;
wire \D_src2[23]~26_combout ;
wire \D_src2[23]~27_combout ;
wire \E_src2[23]~q ;
wire \Add24~130 ;
wire \Add24~125_sumout ;
wire \E_alu_result[24]~combout ;
wire \M_alu_result[24]~q ;
wire \M_rot[0]~29_combout ;
wire \A_shift_rot_result~29_combout ;
wire \A_shift_rot_result[24]~q ;
wire \A_slow_inst_result_nxt[24]~29_combout ;
wire \A_slow_inst_result[24]~q ;
wire \A_wr_data_unfiltered[24]~63_combout ;
wire \A_wr_data_unfiltered[24]~64_combout ;
wire \W_wr_data[24]~q ;
wire \D_src1_reg[24]~29_combout ;
wire \E_src1[24]~q ;
wire \E_alu_result~29_combout ;
wire \D_src2_reg[24]~56_combout ;
wire \D_src2_reg[24]~57_combout ;
wire \D_src2[24]~24_combout ;
wire \D_src2[24]~25_combout ;
wire \E_src2[24]~q ;
wire \Add24~126 ;
wire \Add24~97_sumout ;
wire \E_alu_result[25]~combout ;
wire \M_alu_result[25]~q ;
wire \A_inst_result[25]~q ;
wire \E_rot_step1[21]~21_combout ;
wire \E_rot_step1[25]~18_combout ;
wire \M_rot_prestep2[25]~q ;
wire \E_rot_step1[29]~19_combout ;
wire \E_rot_step1[1]~16_combout ;
wire \M_rot_prestep2[1]~q ;
wire \M_rot[1]~21_combout ;
wire \A_shift_rot_result~21_combout ;
wire \A_shift_rot_result[25]~q ;
wire \A_slow_inst_result_nxt[25]~21_combout ;
wire \A_slow_inst_result[25]~q ;
wire \A_wr_data_unfiltered[25]~47_combout ;
wire \A_wr_data_unfiltered[25]~48_combout ;
wire \W_wr_data[25]~q ;
wire \D_src1_reg[25]~20_combout ;
wire \E_src1[25]~q ;
wire \E_alu_result~22_combout ;
wire \D_src2_reg[25]~42_combout ;
wire \D_src2_reg[25]~43_combout ;
wire \D_src2[25]~12_combout ;
wire \D_src2[25]~13_combout ;
wire \E_src2[25]~q ;
wire \Add24~98 ;
wire \Add24~93_sumout ;
wire \E_alu_result[26]~combout ;
wire \M_alu_result[26]~q ;
wire \A_inst_result[26]~q ;
wire \E_rot_step1[22]~10_combout ;
wire \M_rot_prestep2[26]~q ;
wire \M_rot_prestep2[2]~q ;
wire \M_rot[2]~20_combout ;
wire \A_shift_rot_result~20_combout ;
wire \A_shift_rot_result[26]~q ;
wire \A_slow_inst_result_nxt[26]~20_combout ;
wire \A_slow_inst_result[26]~q ;
wire \A_wr_data_unfiltered[26]~45_combout ;
wire \A_wr_data_unfiltered[26]~46_combout ;
wire \W_wr_data[26]~q ;
wire \D_src1_reg[26]~19_combout ;
wire \E_src1[26]~q ;
wire \E_alu_result~21_combout ;
wire \D_src2_reg[26]~40_combout ;
wire \D_src2_reg[26]~41_combout ;
wire \D_src2[26]~10_combout ;
wire \D_src2[26]~11_combout ;
wire \E_src2[26]~q ;
wire \Add24~94 ;
wire \Add24~89_sumout ;
wire \E_alu_result[27]~combout ;
wire \M_alu_result[27]~q ;
wire \M_rot[3]~18_combout ;
wire \A_shift_rot_result~18_combout ;
wire \A_shift_rot_result[27]~q ;
wire \A_slow_inst_result_nxt[27]~18_combout ;
wire \A_slow_inst_result[27]~q ;
wire \A_wr_data_unfiltered[27]~41_combout ;
wire \A_wr_data_unfiltered[27]~42_combout ;
wire \W_wr_data[27]~q ;
wire \D_src1_reg[27]~17_combout ;
wire \E_src1[27]~q ;
wire \E_logic_result[27]~11_combout ;
wire \E_alu_result~19_combout ;
wire \D_src2_reg[27]~36_combout ;
wire \D_src2_reg[27]~37_combout ;
wire \D_src2[27]~6_combout ;
wire \D_src2[27]~7_combout ;
wire \E_src2[27]~q ;
wire \Add24~90 ;
wire \Add24~85_sumout ;
wire \D_src2_reg[28]~34_combout ;
wire \A_inst_result[28]~q ;
wire \M_rot_prestep2[28]~q ;
wire \M_rot_prestep2[20]~q ;
wire \E_rot_step1[0]~0_combout ;
wire \M_rot_prestep2[4]~q ;
wire \M_rot[4]~17_combout ;
wire \A_shift_rot_result~17_combout ;
wire \A_shift_rot_result[28]~q ;
wire \A_slow_inst_result_nxt[28]~17_combout ;
wire \A_slow_inst_result[28]~q ;
wire \A_wr_data_unfiltered[28]~39_combout ;
wire \A_wr_data_unfiltered[28]~40_combout ;
wire \W_wr_data[28]~q ;
wire \D_src2_reg[28]~35_combout ;
wire \D_src2[28]~4_combout ;
wire \D_src2[28]~5_combout ;
wire \E_src2[28]~q ;
wire \E_logic_result[28]~10_combout ;
wire \E_alu_result~18_combout ;
wire \E_alu_result[28]~combout ;
wire \M_alu_result[28]~q ;
wire \D_src1_reg[28]~16_combout ;
wire \E_src1[28]~q ;
wire \E_rot_step1[28]~3_combout ;
wire \M_rot_prestep2[0]~q ;
wire \M_rot[0]~8_combout ;
wire \A_shift_rot_result~8_combout ;
wire \A_shift_rot_result[8]~q ;
wire \A_slow_inst_result_nxt[8]~8_combout ;
wire \A_slow_inst_result[8]~q ;
wire \A_wr_data_unfiltered[8]~20_combout ;
wire \A_wr_data_unfiltered[8]~21_combout ;
wire \W_wr_data[8]~q ;
wire \D_src2_reg[8]~18_combout ;
wire \D_src2_reg[8]~95_combout ;
wire \E_logic_result[8]~4_combout ;
wire \E_alu_result[8]~8_combout ;
wire \D_src2_reg[8]~111_combout ;
wire \E_src2[8]~q ;
wire \Add24~1_sumout ;
wire \E_alu_result[8]~combout ;
wire \M_alu_result[8]~q ;
wire \D_src1_reg[8]~7_combout ;
wire \E_src1[8]~q ;
wire \E_rot_step1[8]~6_combout ;
wire \M_rot_prestep2[12]~q ;
wire \M_rot[4]~4_combout ;
wire \A_shift_rot_result~4_combout ;
wire \A_shift_rot_result[12]~q ;
wire \A_inst_result[12]~q ;
wire \A_slow_inst_result_nxt[12]~4_combout ;
wire \A_slow_inst_result[12]~q ;
wire \A_wr_data_unfiltered[12]~12_combout ;
wire \A_wr_data_unfiltered[12]~13_combout ;
wire \W_wr_data[12]~q ;
wire \D_src2_reg[12]~14_combout ;
wire \D_src2_reg[12]~91_combout ;
wire \E_logic_result[12]~0_combout ;
wire \E_alu_result[12]~4_combout ;
wire \D_src2_reg[12]~127_combout ;
wire \E_src2[12]~q ;
wire \Add24~41_sumout ;
wire \E_alu_result[12]~combout ;
wire \M_alu_result[12]~q ;
wire \D_src1_reg[12]~3_combout ;
wire \E_src1[12]~q ;
wire \E_rot_step1[13]~23_combout ;
wire \M_rot_prestep2[17]~q ;
wire \M_rot[1]~24_combout ;
wire \A_shift_rot_result~24_combout ;
wire \A_shift_rot_result[17]~q ;
wire \A_slow_inst_result_nxt[17]~24_combout ;
wire \A_slow_inst_result[17]~q ;
wire \A_wr_data_unfiltered[17]~53_combout ;
wire \A_wr_data_unfiltered[17]~54_combout ;
wire \W_wr_data[17]~q ;
wire \D_src2_reg[17]~47_combout ;
wire \Add24~105_sumout ;
wire \D_src2_reg[17]~48_combout ;
wire \D_src2[17]~15_combout ;
wire \D_src2[17]~16_combout ;
wire \E_src2[17]~q ;
wire \E_alu_result~24_combout ;
wire \E_alu_result[17]~combout ;
wire \M_alu_result[17]~q ;
wire \D_src1_reg[17]~24_combout ;
wire \E_src1[17]~q ;
wire \E_rot_step1[17]~20_combout ;
wire \M_rot_prestep2[21]~q ;
wire \M_rot_prestep2[5]~q ;
wire \M_rot_prestep2[29]~q ;
wire \M_rot[5]~26_combout ;
wire \A_shift_rot_result~26_combout ;
wire \A_shift_rot_result[21]~q ;
wire \A_slow_inst_result_nxt[21]~26_combout ;
wire \A_slow_inst_result[21]~q ;
wire \A_wr_data_unfiltered[21]~57_combout ;
wire \A_wr_data_unfiltered[21]~58_combout ;
wire \W_wr_data[21]~q ;
wire \D_src1_reg[21]~26_combout ;
wire \E_src1[21]~q ;
wire \Add24~113_sumout ;
wire \D_src2_reg[21]~51_combout ;
wire \D_src2_reg[21]~52_combout ;
wire \D_src2[21]~19_combout ;
wire \D_src2[21]~20_combout ;
wire \E_src2[21]~q ;
wire \E_logic_result[21]~14_combout ;
wire \E_alu_result~26_combout ;
wire \E_alu_result[21]~combout ;
wire \M_alu_result[21]~q ;
wire \A_inst_result[21]~q ;
wire \A_inst_result[13]~q ;
wire \A_wr_data_unfiltered[5]~8_combout ;
wire \M_rot[5]~3_combout ;
wire \A_shift_rot_result~3_combout ;
wire \A_shift_rot_result[5]~q ;
wire \A_wr_data_unfiltered[5]~9_combout ;
wire \W_wr_data[5]~q ;
wire \D_src2_reg[5]~11_combout ;
wire \D_src2_reg[5]~12_combout ;
wire \E_src2[5]~q ;
wire \Add24~17_sumout ;
wire \E_alu_result~3_combout ;
wire \E_alu_result[5]~combout ;
wire \M_alu_result[5]~q ;
wire \D_src1_reg[5]~2_combout ;
wire \E_src1[5]~q ;
wire \E_rot_step1[5]~17_combout ;
wire \M_rot_prestep2[9]~q ;
wire \M_rot[1]~7_combout ;
wire \A_shift_rot_result~7_combout ;
wire \A_shift_rot_result[9]~q ;
wire \A_inst_result[9]~q ;
wire \A_slow_inst_result_nxt[9]~7_combout ;
wire \A_slow_inst_result[9]~q ;
wire \A_wr_data_unfiltered[9]~18_combout ;
wire \A_wr_data_unfiltered[9]~19_combout ;
wire \W_wr_data[9]~q ;
wire \D_src2_reg[9]~17_combout ;
wire \D_src2_reg[9]~94_combout ;
wire \E_logic_result[9]~3_combout ;
wire \E_alu_result[9]~7_combout ;
wire \D_src2_reg[9]~115_combout ;
wire \E_src2[9]~q ;
wire \Add24~5_sumout ;
wire \E_alu_result[9]~combout ;
wire \M_alu_result[9]~q ;
wire \D_src1_reg[9]~6_combout ;
wire \E_src1[9]~q ;
wire \E_rot_step1[9]~22_combout ;
wire \M_rot_prestep2[13]~q ;
wire \M_rot[5]~14_combout ;
wire \A_shift_rot_result~14_combout ;
wire \A_shift_rot_result[13]~q ;
wire \A_slow_inst_result_nxt[13]~14_combout ;
wire \A_slow_inst_result[13]~q ;
wire \A_wr_data_unfiltered[13]~33_combout ;
wire \A_wr_data_unfiltered[13]~34_combout ;
wire \W_wr_data[13]~q ;
wire \D_src2_reg[13]~27_combout ;
wire \D_src2_reg[13]~98_combout ;
wire \E_logic_result[13]~8_combout ;
wire \E_alu_result[13]~14_combout ;
wire \D_src2_reg[13]~99_combout ;
wire \E_src2[13]~q ;
wire \Add24~61_sumout ;
wire \E_alu_result[13]~combout ;
wire \M_alu_result[13]~q ;
wire \D_src1_reg[13]~13_combout ;
wire \E_src1[13]~q ;
wire \E_rot_step1[14]~12_combout ;
wire \M_rot_prestep2[18]~q ;
wire \M_rot[2]~28_combout ;
wire \A_shift_rot_result~28_combout ;
wire \A_shift_rot_result[18]~q ;
wire \A_slow_inst_result_nxt[18]~28_combout ;
wire \A_slow_inst_result[18]~q ;
wire \A_wr_data_unfiltered[18]~61_combout ;
wire \A_wr_data_unfiltered[18]~62_combout ;
wire \W_wr_data[18]~q ;
wire \D_src2_reg[18]~54_combout ;
wire \Add24~121_sumout ;
wire \D_src2_reg[18]~55_combout ;
wire \D_src2[18]~22_combout ;
wire \D_src2[18]~23_combout ;
wire \E_src2[18]~q ;
wire \E_alu_result~28_combout ;
wire \E_alu_result[18]~combout ;
wire \M_alu_result[18]~q ;
wire \D_src1_reg[18]~28_combout ;
wire \E_src1[18]~q ;
wire \E_rot_step1[18]~13_combout ;
wire \M_rot_prestep2[22]~q ;
wire \M_rot[6]~25_combout ;
wire \A_shift_rot_result~25_combout ;
wire \A_shift_rot_result[22]~q ;
wire \A_slow_inst_result_nxt[22]~25_combout ;
wire \A_slow_inst_result[22]~q ;
wire \A_wr_data_unfiltered[22]~55_combout ;
wire \A_wr_data_unfiltered[22]~56_combout ;
wire \W_wr_data[22]~q ;
wire \D_src1_reg[22]~25_combout ;
wire \E_src1[22]~q ;
wire \Add24~109_sumout ;
wire \D_src2_reg[22]~49_combout ;
wire \D_src2_reg[22]~50_combout ;
wire \D_src2[22]~17_combout ;
wire \D_src2[22]~18_combout ;
wire \E_src2[22]~q ;
wire \E_logic_result[22]~13_combout ;
wire \E_alu_result~25_combout ;
wire \E_alu_result[22]~combout ;
wire \M_alu_result[22]~q ;
wire \A_inst_result[22]~q ;
wire \A_inst_result[14]~q ;
wire \A_wr_data_unfiltered[6]~24_combout ;
wire \M_rot[6]~10_combout ;
wire \A_shift_rot_result~10_combout ;
wire \A_shift_rot_result[6]~q ;
wire \A_wr_data_unfiltered[6]~25_combout ;
wire \W_wr_data[6]~q ;
wire \D_src2_reg[6]~21_combout ;
wire \D_src2_reg[6]~22_combout ;
wire \E_src2[6]~q ;
wire \Add24~21_sumout ;
wire \E_alu_result~10_combout ;
wire \E_alu_result[6]~combout ;
wire \M_alu_result[6]~q ;
wire \D_src1_reg[6]~9_combout ;
wire \E_src1[6]~q ;
wire \E_rot_step1[6]~14_combout ;
wire \M_rot_prestep2[10]~q ;
wire \M_rot[2]~6_combout ;
wire \A_shift_rot_result~6_combout ;
wire \A_shift_rot_result[10]~q ;
wire \A_inst_result[10]~q ;
wire \A_slow_inst_result_nxt[10]~6_combout ;
wire \A_slow_inst_result[10]~q ;
wire \A_wr_data_unfiltered[10]~16_combout ;
wire \A_wr_data_unfiltered[10]~17_combout ;
wire \W_wr_data[10]~q ;
wire \D_src2_reg[10]~16_combout ;
wire \D_src2_reg[10]~93_combout ;
wire \E_logic_result[10]~2_combout ;
wire \E_alu_result[10]~6_combout ;
wire \D_src2_reg[10]~119_combout ;
wire \E_src2[10]~q ;
wire \Add24~13_sumout ;
wire \E_alu_result[10]~combout ;
wire \M_alu_result[10]~q ;
wire \D_src1_reg[10]~5_combout ;
wire \E_src1[10]~q ;
wire \E_rot_step1[10]~15_combout ;
wire \M_rot_prestep2[14]~q ;
wire \M_rot[6]~13_combout ;
wire \A_shift_rot_result~13_combout ;
wire \A_shift_rot_result[14]~q ;
wire \A_slow_inst_result_nxt[14]~13_combout ;
wire \A_slow_inst_result[14]~q ;
wire \A_wr_data_unfiltered[14]~31_combout ;
wire \A_wr_data_unfiltered[14]~32_combout ;
wire \W_wr_data[14]~q ;
wire \D_src2_reg[14]~26_combout ;
wire \D_src2_reg[14]~97_combout ;
wire \E_logic_result[14]~7_combout ;
wire \E_alu_result[14]~13_combout ;
wire \D_src2_reg[14]~103_combout ;
wire \E_src2[14]~q ;
wire \Add24~57_sumout ;
wire \E_alu_result[14]~combout ;
wire \M_alu_result[14]~q ;
wire \D_src1_reg[14]~12_combout ;
wire \E_src1[14]~q ;
wire \E_rot_step1[15]~30_combout ;
wire \M_rot_prestep2[19]~q ;
wire \M_rot[3]~22_combout ;
wire \A_shift_rot_result~22_combout ;
wire \A_shift_rot_result[19]~q ;
wire \A_slow_inst_result_nxt[19]~22_combout ;
wire \A_slow_inst_result[19]~q ;
wire \A_wr_data_unfiltered[19]~49_combout ;
wire \A_wr_data_unfiltered[19]~50_combout ;
wire \W_wr_data[19]~q ;
wire \D_src2_reg[19]~89_combout ;
wire \Add24~101_sumout ;
wire \D_src2_reg[19]~90_combout ;
wire \D_src2_reg[19]~44_combout ;
wire \D_src2[19]~14_combout ;
wire \E_src2[19]~q ;
wire \E_alu_result~23_combout ;
wire \E_alu_result[19]~combout ;
wire \M_alu_result[19]~q ;
wire \A_inst_result[19]~q ;
wire \A_wr_data_unfiltered[3]~35_combout ;
wire \M_rot[3]~15_combout ;
wire \A_shift_rot_result~15_combout ;
wire \A_shift_rot_result[3]~q ;
wire \A_wr_data_unfiltered[3]~36_combout ;
wire \W_wr_data[3]~q ;
wire \D_src1_reg[3]~14_combout ;
wire \E_src1[3]~q ;
wire \Add24~29_sumout ;
wire \E_alu_result~15_combout ;
wire \E_alu_result[3]~combout ;
wire \M_alu_result[3]~q ;
wire \D_src2_reg[3]~28_combout ;
wire \D_src2_reg[3]~29_combout ;
wire \E_src2[3]~q ;
wire \E_rot_pass2~0_combout ;
wire \M_rot_pass2~q ;
wire \M_rot[4]~27_combout ;
wire \A_shift_rot_result~27_combout ;
wire \A_shift_rot_result[20]~q ;
wire \A_slow_inst_result_nxt[20]~27_combout ;
wire \A_slow_inst_result[20]~q ;
wire \A_wr_data_unfiltered[20]~59_combout ;
wire \A_wr_data_unfiltered[20]~60_combout ;
wire \W_wr_data[20]~q ;
wire \D_src2_reg[20]~87_combout ;
wire \Add24~117_sumout ;
wire \D_src2_reg[20]~88_combout ;
wire \D_src2_reg[20]~53_combout ;
wire \D_src2[20]~21_combout ;
wire \E_src2[20]~q ;
wire \E_alu_result~27_combout ;
wire \E_alu_result[20]~combout ;
wire \M_alu_result[20]~q ;
wire \A_inst_result[20]~q ;
wire \A_wr_data_unfiltered[4]~0_combout ;
wire \M_rot[4]~0_combout ;
wire \A_shift_rot_result~0_combout ;
wire \A_shift_rot_result[4]~q ;
wire \A_wr_data_unfiltered[4]~3_combout ;
wire \W_wr_data[4]~q ;
wire \D_src2_reg[4]~5_combout ;
wire \D_src2_reg[4]~6_combout ;
wire \E_src2[4]~q ;
wire \Add24~33_sumout ;
wire \E_alu_result~1_combout ;
wire \E_alu_result[4]~combout ;
wire \M_alu_result[4]~q ;
wire \A_mem_baddr[4]~q ;
wire \M_sel_data_master~q ;
wire \M_ctrl_st_nxt~0_combout ;
wire \E_st_cache~0_combout ;
wire \M_ctrl_st_non_bypass~q ;
wire \M_dc_valid_st_cache_hit~0_combout ;
wire \M_dc_valid_st_cache_hit~1_combout ;
wire \A_dc_valid_st_cache_hit~q ;
wire \A_mem_baddr[10]~q ;
wire \A_mem_baddr[7]~q ;
wire \A_mem_baddr[5]~q ;
wire \A_mem_baddr[6]~q ;
wire \Equal261~0_combout ;
wire \A_mem_baddr[9]~q ;
wire \A_mem_baddr[8]~q ;
wire \Equal261~1_combout ;
wire \Equal261~2_combout ;
wire \M_dc_dirty~combout ;
wire \A_dc_dirty~q ;
wire \A_dc_xfer_rd_addr_has_started_nxt~0_combout ;
wire \A_dc_xfer_rd_addr_has_started~q ;
wire \Equal191~0_combout ;
wire \M_ctrl_dc_index_wb_inv~q ;
wire \A_ctrl_dc_index_wb_inv~q ;
wire \A_dc_hit~q ;
wire \E_ctrl_dc_addr_inv~0_combout ;
wire \Equal179~0_combout ;
wire \M_ctrl_dc_addr_wb_inv~q ;
wire \A_ctrl_dc_addr_wb_inv~q ;
wire \A_dc_xfer_rd_addr_starting~0_combout ;
wire \A_dc_xfer_rd_addr_starting~1_combout ;
wire \A_dc_xfer_rd_data_starting~q ;
wire \A_dc_xfer_wr_starting~q ;
wire \A_dc_wb_rd_addr_starting~q ;
wire \A_dc_wb_rd_data_starting~q ;
wire \A_dc_wb_rd_data_first_nxt~0_combout ;
wire \A_dc_wb_rd_data_first~q ;
wire \A_dc_wb_wr_starting~combout ;
wire \av_wr_data_transfer~0_combout ;
wire \A_dc_wr_data_cnt_nxt[0]~3_combout ;
wire \A_dc_wb_wr_active_nxt~0_combout ;
wire \A_dc_wb_wr_active~q ;
wire \A_dc_wr_data_cnt[0]~0_combout ;
wire \A_dc_wr_data_cnt[0]~q ;
wire \A_dc_wr_data_cnt_nxt[1]~2_combout ;
wire \A_dc_wr_data_cnt[1]~q ;
wire \A_dc_wr_data_cnt_nxt[2]~1_combout ;
wire \A_dc_wr_data_cnt[2]~q ;
wire \A_dc_wr_data_cnt_nxt[3]~0_combout ;
wire \A_dc_wr_data_cnt[3]~q ;
wire \A_dc_wb_active_nxt~0_combout ;
wire \A_dc_wb_active~q ;
wire \A_dc_fill_has_started_nxt~0_combout ;
wire \A_dc_fill_has_started~q ;
wire \A_dc_fill_starting~0_combout ;
wire \A_dc_fill_dp_offset_nxt[0]~1_combout ;
wire \A_dc_rd_data_cnt[0]~1_combout ;
wire \A_dc_fill_dp_offset[0]~q ;
wire \A_dc_fill_dp_offset_nxt[1]~2_combout ;
wire \A_dc_fill_dp_offset[1]~q ;
wire \A_dc_fill_dp_offset_nxt[2]~0_combout ;
wire \A_dc_fill_dp_offset[2]~q ;
wire \Equal263~0_combout ;
wire \A_mem_baddr[3]~q ;
wire \A_dc_rd_data_cnt_nxt[0]~3_combout ;
wire \A_dc_rd_data_cnt[0]~0_combout ;
wire \A_dc_rd_data_cnt[0]~q ;
wire \A_dc_rd_data_cnt_nxt[1]~2_combout ;
wire \A_dc_rd_data_cnt[1]~q ;
wire \A_dc_rd_data_cnt_nxt[2]~1_combout ;
wire \A_dc_rd_data_cnt[2]~q ;
wire \A_dc_rd_data_cnt_nxt[3]~0_combout ;
wire \A_dc_rd_data_cnt[3]~q ;
wire \A_ld_bypass_done~combout ;
wire \M_ctrl_ld_st_nxt~0_combout ;
wire \M_ctrl_ld_st~q ;
wire \M_valid_mem_d1~0_combout ;
wire \M_valid_mem_d1~q ;
wire \M_A_dc_line_match_d1~q ;
wire \A_dc_fill_need_extra_stall_nxt~combout ;
wire \A_dc_fill_need_extra_stall~q ;
wire \A_dc_rd_last_transfer_d1~q ;
wire \A_dc_fill_active_nxt~0_combout ;
wire \A_dc_fill_active~q ;
wire \A_mem_baddr[2]~q ;
wire \A_dc_fill_wr_data~0_combout ;
wire \A_slow_inst_result_en~0_combout ;
wire \A_slow_inst_result[2]~q ;
wire \A_inst_result[2]~q ;
wire \A_wr_data_unfiltered[2]~6_combout ;
wire \M_rot[2]~2_combout ;
wire \A_shift_rot_result~2_combout ;
wire \A_shift_rot_result[2]~q ;
wire \A_wr_data_unfiltered[2]~7_combout ;
wire \W_wr_data[2]~q ;
wire \D_src1_reg[2]~1_combout ;
wire \E_src1[2]~q ;
wire \Add24~25_sumout ;
wire \E_alu_result~2_combout ;
wire \E_alu_result[2]~combout ;
wire \M_alu_result[2]~q ;
wire \D_src2_reg[2]~9_combout ;
wire \D_src2_reg[2]~10_combout ;
wire \E_src2[2]~q ;
wire \E_rot_mask[5]~3_combout ;
wire \M_rot_mask[5]~q ;
wire \M_rot[5]~16_combout ;
wire \A_shift_rot_result~16_combout ;
wire \A_shift_rot_result[29]~q ;
wire \A_slow_inst_result_nxt[29]~16_combout ;
wire \A_slow_inst_result[29]~q ;
wire \A_wr_data_unfiltered[29]~37_combout ;
wire \A_wr_data_unfiltered[29]~38_combout ;
wire \W_wr_data[29]~q ;
wire \D_src1_reg[29]~15_combout ;
wire \E_src1[29]~q ;
wire \Add24~81_sumout ;
wire \D_src2_reg[29]~32_combout ;
wire \D_src2_reg[29]~33_combout ;
wire \D_src2[29]~2_combout ;
wire \D_src2[29]~3_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~9_combout ;
wire \Equal305~0_combout ;
wire \Equal305~1_combout ;
wire \Equal305~2_combout ;
wire \Equal305~3_combout ;
wire \Equal305~4_combout ;
wire \Equal305~5_combout ;
wire \Equal305~6_combout ;
wire \Equal305~7_combout ;
wire \Equal305~8_combout ;
wire \Equal305~9_combout ;
wire \Equal305~10_combout ;
wire \Equal305~11_combout ;
wire \Equal305~12_combout ;
wire \Equal305~13_combout ;
wire \Equal305~14_combout ;
wire \Equal305~15_combout ;
wire \E_compare_op[1]~q ;
wire \E_br_result~0_combout ;
wire \E_br_result~1_combout ;
wire \E_logic_result[0]~15_combout ;
wire \Add24~73_sumout ;
wire \E_alu_result[0]~16_combout ;
wire \E_alu_result[0]~combout ;
wire \M_alu_result[0]~q ;
wire \M_ld_align_sh8~0_combout ;
wire \A_ld_align_sh8~q ;
wire \A_slow_inst_result_nxt[1]~23_combout ;
wire \A_slow_inst_result[1]~q ;
wire \M_inst_result[1]~1_combout ;
wire \A_ienable_reg_irq1~q ;
wire \A_ipending_reg_irq1_nxt~combout ;
wire \A_ipending_reg_irq1~q ;
wire \D_control_reg_rddata_muxed[1]~2_combout ;
wire \E_control_reg_rddata[1]~q ;
wire \M_control_reg_rddata[1]~q ;
wire \A_inst_result[1]~q ;
wire \A_wr_data_unfiltered[1]~51_combout ;
wire \M_rot[1]~23_combout ;
wire \A_shift_rot_result~23_combout ;
wire \A_shift_rot_result[1]~q ;
wire \A_wr_data_unfiltered[1]~52_combout ;
wire \W_wr_data[1]~q ;
wire \D_src2_reg[1]~45_combout ;
wire \D_src2_reg[1]~46_combout ;
wire \E_src2[1]~q ;
wire \Add24~69_sumout ;
wire \E_logic_result[1]~16_combout ;
wire \E_alu_result[1]~combout ;
wire \M_alu_result[1]~q ;
wire \M_data_ram_ld_align_sign_bit_16_hi~0_combout ;
wire \M_data_ram_ld_align_sign_bit_16_hi~q ;
wire \M_data_ram_ld_align_sign_bit~0_combout ;
wire \A_data_ram_ld_align_sign_bit~q ;
wire \M_rot[0]~11_combout ;
wire \A_shift_rot_result~11_combout ;
wire \A_shift_rot_result[16]~q ;
wire \A_slow_inst_result_nxt[16]~11_combout ;
wire \A_slow_inst_result[16]~q ;
wire \A_wr_data_unfiltered[16]~27_combout ;
wire \A_wr_data_unfiltered[16]~28_combout ;
wire \W_wr_data[16]~q ;
wire \D_src2_reg[16]~23_combout ;
wire \E_logic_result[16]~5_combout ;
wire \E_alu_result[16]~11_combout ;
wire \D_src2_reg[16]~24_combout ;
wire \D_src2[16]~0_combout ;
wire \D_src2[16]~1_combout ;
wire \E_src2[16]~q ;
wire \Add24~49_sumout ;
wire \E_alu_result[16]~combout ;
wire \M_alu_result[16]~q ;
wire \M_dc_hit~0_combout ;
wire \M_dc_hit~1_combout ;
wire \M_dc_hit~combout ;
wire \M_dc_valid_st_bypass_hit~0_combout ;
wire \A_dc_valid_st_bypass_hit~q ;
wire \A_st_bypass_transfer_done~combout ;
wire \A_st_bypass_transfer_done_d1~q ;
wire \A_ctrl_st_bypass~q ;
wire \E_ctrl_dc_nowb_inv~0_combout ;
wire \M_ctrl_dc_nowb_inv~q ;
wire \A_ctrl_dc_nowb_inv~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ;
wire \A_dc_xfer_rd_addr_offset[0]~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ;
wire \A_dc_xfer_rd_addr_offset[1]~q ;
wire \A_dc_xfer_rd_addr_active_nxt~0_combout ;
wire \A_dc_xfer_rd_addr_active~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ;
wire \A_dc_xfer_rd_addr_offset[2]~q ;
wire \A_dc_xfer_rd_addr_done_nxt~combout ;
wire \A_dc_xfer_rd_addr_done~q ;
wire \A_dc_dcache_management_done_nxt~0_combout ;
wire \A_dc_dcache_management_done_nxt~combout ;
wire \A_dc_dcache_management_done~q ;
wire \M_dc_potential_hazard_after_st_unfiltered~0_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~1_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~2_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~3_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~4_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~5_combout ;
wire \A_dc_potential_hazard_after_st~q ;
wire \A_mem_stall_nxt~1_combout ;
wire \A_mem_stall_nxt~2_combout ;
wire \A_mem_stall_nxt~3_combout ;
wire \A_mem_stall_nxt~4_combout ;
wire \A_mem_stall_nxt~5_combout ;
wire \A_mem_stall~q ;
wire \always138~0_combout ;
wire \A_mul_cnt_nxt[0]~2_combout ;
wire \A_mul_cnt[0]~q ;
wire \A_mul_cnt_nxt[1]~1_combout ;
wire \A_mul_cnt[1]~q ;
wire \A_mul_cnt_nxt[2]~0_combout ;
wire \A_mul_cnt[2]~q ;
wire \A_mul_stall_nxt~0_combout ;
wire \A_mul_stall~q ;
wire \A_mul_stall_d1~q ;
wire \A_mul_stall_d2~q ;
wire \A_mul_stall_d3~q ;
wire \A_mul_result[0]~q ;
wire \Add26~6 ;
wire \Add26~93_sumout ;
wire \A_mul_result[1]~q ;
wire \Add26~94 ;
wire \Add26~9_sumout ;
wire \A_mul_result[2]~q ;
wire \Add26~10 ;
wire \Add26~61_sumout ;
wire \A_mul_result[3]~q ;
wire \Add26~62 ;
wire \Add26~1_sumout ;
wire \A_mul_result[4]~q ;
wire \Add26~2 ;
wire \Add26~13_sumout ;
wire \A_mul_result[5]~q ;
wire \Add26~14 ;
wire \Add26~41_sumout ;
wire \A_mul_result[6]~q ;
wire \Add26~42 ;
wire \Add26~37_sumout ;
wire \A_mul_result[7]~q ;
wire \Add26~38 ;
wire \Add26~33_sumout ;
wire \A_mul_result[8]~q ;
wire \Add26~34 ;
wire \Add26~29_sumout ;
wire \A_mul_result[9]~q ;
wire \Add26~30 ;
wire \Add26~25_sumout ;
wire \A_mul_result[10]~q ;
wire \Add26~26 ;
wire \Add26~21_sumout ;
wire \A_mul_result[11]~q ;
wire \Add26~22 ;
wire \Add26~17_sumout ;
wire \A_mul_result[12]~q ;
wire \Add26~18 ;
wire \Add26~57_sumout ;
wire \A_mul_result[13]~q ;
wire \Add26~58 ;
wire \Add26~53_sumout ;
wire \A_mul_result[14]~q ;
wire \Add26~54 ;
wire \Add26~49_sumout ;
wire \A_mul_result[15]~q ;
wire \M_rot[7]~12_combout ;
wire \A_shift_rot_result~12_combout ;
wire \A_shift_rot_result[15]~q ;
wire \A_slow_inst_result_nxt[15]~12_combout ;
wire \A_slow_inst_result[15]~q ;
wire \A_wr_data_unfiltered[15]~29_combout ;
wire \A_wr_data_unfiltered[15]~30_combout ;
wire \W_wr_data[15]~q ;
wire \D_src2_reg[15]~25_combout ;
wire \D_src2_reg[15]~96_combout ;
wire \E_logic_result[15]~6_combout ;
wire \E_alu_result[15]~12_combout ;
wire \D_src2_reg[15]~107_combout ;
wire \E_src2[15]~q ;
wire \Add24~53_sumout ;
wire \E_alu_result[15]~combout ;
wire \M_alu_result[15]~q ;
wire \M_dc_want_fill~0_combout ;
wire \E_ld_st_cache~0_combout ;
wire \M_ctrl_ld_st_non_bypass~q ;
wire \M_dc_want_fill~1_combout ;
wire \M_dc_want_fill~combout ;
wire \A_dc_want_fill~q ;
wire \A_slow_inst_sel_nxt~0_combout ;
wire \A_slow_inst_sel~q ;
wire \A_wr_data_unfiltered[22]~26_combout ;
wire \A_mul_partial_prod[31]~q ;
wire \Add26~78 ;
wire \Add26~125_sumout ;
wire \A_mul_result[31]~q ;
wire \M_rot[7]~31_combout ;
wire \A_shift_rot_result~31_combout ;
wire \A_shift_rot_result[31]~q ;
wire \A_slow_inst_result_nxt[31]~31_combout ;
wire \Add14~78 ;
wire \Add14~125_sumout ;
wire \A_div_quot[31]~q ;
wire \A_slow_inst_result[31]~q ;
wire \A_wr_data_unfiltered[31]~67_combout ;
wire \A_wr_data_unfiltered[31]~68_combout ;
wire \W_wr_data[31]~q ;
wire \D_src1_reg[31]~31_combout ;
wire \E_src1[31]~q ;
wire \Add24~78 ;
wire \Add24~37_sumout ;
wire \D_src2_reg[31]~60_combout ;
wire \D_src2_reg[31]~61_combout ;
wire \D_src2[31]~28_combout ;
wire \D_src2[31]~29_combout ;
wire \E_src2[31]~q ;
wire \Add24~38 ;
wire \Add24~65_sumout ;
wire \E_br_result~2_combout ;
wire \E_ctrl_br_cond~q ;
wire \D_ctrl_flush_pipe_always~0_combout ;
wire \D_ctrl_flush_pipe_always~1_combout ;
wire \E_ctrl_flush_pipe_always~q ;
wire \M_pipe_flush_nxt~0_combout ;
wire \M_pipe_flush~q ;
wire \E_wr_dst_reg_from_D~q ;
wire \E_wr_dst_reg~0_combout ;
wire \E_regnum_b_cmp_F~0_combout ;
wire \E_regnum_b_cmp_F~1_combout ;
wire \E_regnum_b_cmp_F~combout ;
wire \M_regnum_b_cmp_D~q ;
wire \D_src2_reg[29]~0_combout ;
wire \D_src2_reg[29]~1_combout ;
wire \D_src2_reg[0]~7_combout ;
wire \D_src2_reg[0]~8_combout ;
wire \E_src2[0]~q ;
wire \Add9~17_sumout ;
wire \M_div_src2[0]~q ;
wire \A_div_den[0]~0_combout ;
wire \A_div_den[0]~q ;
wire \Add9~18 ;
wire \Add9~21_sumout ;
wire \M_div_src2[1]~q ;
wire \A_div_den_en~combout ;
wire \A_div_den[1]~q ;
wire \Add9~22 ;
wire \Add9~25_sumout ;
wire \M_div_src2[2]~q ;
wire \A_div_den[2]~q ;
wire \Add9~26 ;
wire \Add9~29_sumout ;
wire \M_div_src2[3]~q ;
wire \A_div_den[3]~q ;
wire \Add9~30 ;
wire \Add9~33_sumout ;
wire \M_div_src2[4]~q ;
wire \A_div_den[4]~q ;
wire \Add9~34 ;
wire \Add9~37_sumout ;
wire \M_div_src2[5]~q ;
wire \A_div_den[5]~q ;
wire \Add9~38 ;
wire \Add9~41_sumout ;
wire \M_div_src2[6]~q ;
wire \A_div_den[6]~q ;
wire \Add9~42 ;
wire \Add9~45_sumout ;
wire \M_div_src2[7]~q ;
wire \A_div_den[7]~q ;
wire \Add9~46 ;
wire \Add9~49_sumout ;
wire \M_div_src2[8]~q ;
wire \A_div_den[8]~q ;
wire \Add9~50 ;
wire \Add9~53_sumout ;
wire \M_div_src2[9]~q ;
wire \A_div_den[9]~q ;
wire \Add9~54 ;
wire \Add9~57_sumout ;
wire \M_div_src2[10]~q ;
wire \A_div_den[10]~q ;
wire \Add9~58 ;
wire \Add9~61_sumout ;
wire \M_div_src2[11]~q ;
wire \A_div_den[11]~q ;
wire \Add9~62 ;
wire \Add9~65_sumout ;
wire \M_div_src2[12]~q ;
wire \A_div_den[12]~q ;
wire \Add9~66 ;
wire \Add9~69_sumout ;
wire \M_div_src2[13]~q ;
wire \A_div_den[13]~q ;
wire \Add9~70 ;
wire \Add9~73_sumout ;
wire \M_div_src2[14]~q ;
wire \A_div_den[14]~q ;
wire \Add9~74 ;
wire \Add9~77_sumout ;
wire \M_div_src2[15]~q ;
wire \A_div_den[15]~q ;
wire \Add9~78 ;
wire \Add9~85_sumout ;
wire \M_div_src2[16]~q ;
wire \A_div_den[16]~q ;
wire \Add9~86 ;
wire \Add9~89_sumout ;
wire \M_div_src2[17]~q ;
wire \A_div_den[17]~q ;
wire \Add9~90 ;
wire \Add9~93_sumout ;
wire \M_div_src2[18]~q ;
wire \A_div_den[18]~q ;
wire \Add9~94 ;
wire \Add9~97_sumout ;
wire \M_div_src2[19]~q ;
wire \A_div_den[19]~q ;
wire \Add9~98 ;
wire \Add9~101_sumout ;
wire \M_div_src2[20]~q ;
wire \A_div_den[20]~q ;
wire \Add9~102 ;
wire \Add9~105_sumout ;
wire \M_div_src2[21]~q ;
wire \A_div_den[21]~q ;
wire \Add9~106 ;
wire \Add9~109_sumout ;
wire \M_div_src2[22]~q ;
wire \A_div_den[22]~q ;
wire \Add9~110 ;
wire \Add9~113_sumout ;
wire \M_div_src2[23]~q ;
wire \A_div_den[23]~q ;
wire \Add9~114 ;
wire \Add9~117_sumout ;
wire \M_div_src2[24]~q ;
wire \A_div_den[24]~q ;
wire \Add9~118 ;
wire \Add9~121_sumout ;
wire \M_div_src2[25]~q ;
wire \A_div_den[25]~q ;
wire \Add9~122 ;
wire \Add9~125_sumout ;
wire \M_div_src2[26]~q ;
wire \A_div_den[26]~q ;
wire \Add9~126 ;
wire \Add9~81_sumout ;
wire \M_div_src2[27]~q ;
wire \A_div_den[27]~q ;
wire \Add9~82 ;
wire \Add9~13_sumout ;
wire \M_div_src2[28]~q ;
wire \A_div_den[28]~q ;
wire \Add9~14 ;
wire \Add9~9_sumout ;
wire \M_div_src2[29]~q ;
wire \A_div_den[29]~q ;
wire \Add9~10 ;
wire \Add9~5_sumout ;
wire \M_div_src2[30]~q ;
wire \A_div_den[30]~q ;
wire \Add9~6 ;
wire \Add9~1_sumout ;
wire \M_div_src2[31]~q ;
wire \A_div_den[31]~q ;
wire \Add8~9_sumout ;
wire \M_div_src1[0]~q ;
wire \A_div_rem[0]~0_combout ;
wire \A_div_rem[0]~q ;
wire \Add11~134_cout ;
wire \Add11~129_sumout ;
wire \Add8~10 ;
wire \Add8~13_sumout ;
wire \M_div_src1[1]~q ;
wire \A_div_rem_en~combout ;
wire \A_div_rem[1]~q ;
wire \Add11~130 ;
wire \Add11~125_sumout ;
wire \Add8~14 ;
wire \Add8~17_sumout ;
wire \M_div_src1[2]~q ;
wire \A_div_rem[2]~q ;
wire \Add11~126 ;
wire \Add11~121_sumout ;
wire \Add8~18 ;
wire \Add8~21_sumout ;
wire \M_div_src1[3]~q ;
wire \A_div_rem[3]~q ;
wire \Add11~122 ;
wire \Add11~117_sumout ;
wire \Add8~22 ;
wire \Add8~25_sumout ;
wire \M_div_src1[4]~q ;
wire \A_div_rem[4]~q ;
wire \Add11~118 ;
wire \Add11~113_sumout ;
wire \Add8~26 ;
wire \Add8~29_sumout ;
wire \M_div_src1[5]~q ;
wire \A_div_rem[5]~q ;
wire \Add11~114 ;
wire \Add11~109_sumout ;
wire \Add8~30 ;
wire \Add8~33_sumout ;
wire \M_div_src1[6]~q ;
wire \A_div_rem[6]~q ;
wire \Add11~110 ;
wire \Add11~105_sumout ;
wire \Add8~34 ;
wire \Add8~37_sumout ;
wire \M_div_src1[7]~q ;
wire \A_div_rem[7]~q ;
wire \Add11~106 ;
wire \Add11~101_sumout ;
wire \Add8~38 ;
wire \Add8~41_sumout ;
wire \M_div_src1[8]~q ;
wire \A_div_rem[8]~q ;
wire \Add11~102 ;
wire \Add11~97_sumout ;
wire \Add8~42 ;
wire \Add8~45_sumout ;
wire \M_div_src1[9]~q ;
wire \A_div_rem[9]~q ;
wire \Add11~98 ;
wire \Add11~93_sumout ;
wire \Add8~46 ;
wire \Add8~49_sumout ;
wire \M_div_src1[10]~q ;
wire \A_div_rem[10]~q ;
wire \Add11~94 ;
wire \Add11~89_sumout ;
wire \Add8~50 ;
wire \Add8~53_sumout ;
wire \M_div_src1[11]~q ;
wire \A_div_rem[11]~q ;
wire \Add11~90 ;
wire \Add11~85_sumout ;
wire \Add8~54 ;
wire \Add8~57_sumout ;
wire \M_div_src1[12]~q ;
wire \A_div_rem[12]~q ;
wire \Add11~86 ;
wire \Add11~81_sumout ;
wire \Add8~58 ;
wire \Add8~61_sumout ;
wire \M_div_src1[13]~q ;
wire \A_div_rem[13]~q ;
wire \Add11~82 ;
wire \Add11~77_sumout ;
wire \Add8~62 ;
wire \Add8~65_sumout ;
wire \M_div_src1[14]~q ;
wire \A_div_rem[14]~q ;
wire \Add11~78 ;
wire \Add11~73_sumout ;
wire \Add8~66 ;
wire \Add8~69_sumout ;
wire \M_div_src1[15]~q ;
wire \A_div_rem[15]~q ;
wire \Add11~74 ;
wire \Add11~69_sumout ;
wire \Add8~70 ;
wire \Add8~77_sumout ;
wire \M_div_src1[16]~q ;
wire \A_div_rem[16]~q ;
wire \Add11~70 ;
wire \Add11~65_sumout ;
wire \Add8~78 ;
wire \Add8~81_sumout ;
wire \M_div_src1[17]~q ;
wire \A_div_rem[17]~q ;
wire \Add11~66 ;
wire \Add11~61_sumout ;
wire \Add8~82 ;
wire \Add8~85_sumout ;
wire \M_div_src1[18]~q ;
wire \A_div_rem[18]~q ;
wire \Add11~62 ;
wire \Add11~57_sumout ;
wire \Add8~86 ;
wire \Add8~89_sumout ;
wire \M_div_src1[19]~q ;
wire \A_div_rem[19]~q ;
wire \Add11~58 ;
wire \Add11~53_sumout ;
wire \Add8~90 ;
wire \Add8~93_sumout ;
wire \M_div_src1[20]~q ;
wire \A_div_rem[20]~q ;
wire \Add11~54 ;
wire \Add11~49_sumout ;
wire \Add8~94 ;
wire \Add8~97_sumout ;
wire \M_div_src1[21]~q ;
wire \A_div_rem[21]~q ;
wire \Add11~50 ;
wire \Add11~45_sumout ;
wire \Add8~98 ;
wire \Add8~101_sumout ;
wire \M_div_src1[22]~q ;
wire \A_div_rem[22]~q ;
wire \Add11~46 ;
wire \Add11~41_sumout ;
wire \Add8~102 ;
wire \Add8~105_sumout ;
wire \M_div_src1[23]~q ;
wire \A_div_rem[23]~q ;
wire \Add11~42 ;
wire \Add11~37_sumout ;
wire \Add8~106 ;
wire \Add8~109_sumout ;
wire \M_div_src1[24]~q ;
wire \A_div_rem[24]~q ;
wire \Add11~38 ;
wire \Add11~33_sumout ;
wire \Add8~110 ;
wire \Add8~113_sumout ;
wire \M_div_src1[25]~q ;
wire \A_div_rem[25]~q ;
wire \Add11~34 ;
wire \Add11~29_sumout ;
wire \Add8~114 ;
wire \Add8~117_sumout ;
wire \M_div_src1[26]~q ;
wire \A_div_rem[26]~q ;
wire \Add11~30 ;
wire \Add11~25_sumout ;
wire \Add8~118 ;
wire \Add8~121_sumout ;
wire \M_div_src1[27]~q ;
wire \A_div_rem[27]~q ;
wire \Add11~26 ;
wire \Add11~21_sumout ;
wire \Add8~122 ;
wire \Add8~125_sumout ;
wire \M_div_src1[28]~q ;
wire \A_div_rem[28]~q ;
wire \Add11~22 ;
wire \Add11~17_sumout ;
wire \Add8~126 ;
wire \Add8~73_sumout ;
wire \M_div_src1[29]~q ;
wire \A_div_rem[29]~q ;
wire \Add11~18 ;
wire \Add11~13_sumout ;
wire \Add8~74 ;
wire \Add8~5_sumout ;
wire \M_div_src1[30]~q ;
wire \A_div_rem[30]~q ;
wire \Add11~14 ;
wire \Add11~9_sumout ;
wire \Add8~6 ;
wire \Add8~1_sumout ;
wire \M_div_src1[31]~q ;
wire \A_div_rem[31]~q ;
wire \Add11~10 ;
wire \Add11~5_sumout ;
wire \A_div_rem[32]~q ;
wire \Add11~6 ;
wire \Add11~1_sumout ;
wire \A_div_discover_quotient_bits~combout ;
wire \Add13~9_sumout ;
wire \A_div_norm_cnt_nxt[0]~0_combout ;
wire \A_div_norm_cnt[0]~q ;
wire \Add13~10 ;
wire \Add13~17_sumout ;
wire \A_div_norm_cnt[1]~q ;
wire \Add13~18 ;
wire \Add13~21_sumout ;
wire \A_div_norm_cnt[2]~q ;
wire \Add13~22 ;
wire \Add13~5_sumout ;
wire \A_div_norm_cnt[3]~q ;
wire \Add13~6 ;
wire \Add13~13_sumout ;
wire \A_div_norm_cnt[4]~q ;
wire \Add13~14 ;
wire \Add13~1_sumout ;
wire \A_div_norm_cnt[5]~q ;
wire \A_div_last_quotient_bit_nxt~0_combout ;
wire \A_div_last_quotient_bit_nxt~combout ;
wire \A_div_last_quotient_bit~q ;
wire \A_div_quot_ready~q ;
wire \A_div_done~q ;
wire \A_stall~combout ;
wire \M_ctrl_late_result~q ;
wire \D_data_depend~1_combout ;
wire \D_dep_stall~0_combout ;
wire \F_stall~combout ;
wire \D_iw[14]~q ;
wire \D_ctrl_break~0_combout ;
wire \E_ctrl_break~q ;
wire \M_ctrl_break~q ;
wire \M_iw[14]~q ;
wire \M_iw[11]~q ;
wire \M_iw[5]~q ;
wire \M_iw[0]~q ;
wire \M_iw[16]~q ;
wire \M_iw[15]~q ;
wire \M_iw[13]~q ;
wire \M_iw[12]~q ;
wire \M_op_eret~0_combout ;
wire \M_iw[4]~q ;
wire \M_iw[3]~q ;
wire \M_iw[2]~q ;
wire \M_iw[1]~q ;
wire \M_op_eret~1_combout ;
wire \M_op_eret~2_combout ;
wire \A_status_reg_pie_inst_nxt~0_combout ;
wire \A_status_reg_pie_inst_nxt~1_combout ;
wire \A_status_reg_pie_inst_nxt~2_combout ;
wire \A_status_reg_pie~q ;
wire \A_valid_wrctl_ienable~q ;
wire \norm_intr_req~0_combout ;
wire \F_iw[5]~1_combout ;
wire \D_iw[5]~q ;
wire \Equal169~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_late_result~2_combout ;
wire \D_ctrl_late_result~0_combout ;
wire \D_ctrl_late_result~1_combout ;
wire \E_ctrl_late_result~q ;
wire \D_data_depend~0_combout ;
wire \D_valid~combout ;
wire \E_valid_from_D~q ;
wire \E_valid~0_combout ;
wire \latched_oci_tb_hbreak_req_next~0_combout ;
wire \latched_oci_tb_hbreak_req~q ;
wire \F_iw~0_combout ;
wire \F_iw[0]~9_combout ;
wire \D_iw[0]~q ;
wire \E_iw[0]~q ;
wire \E_ld_st_bus~0_combout ;
wire \M_ctrl_ld_st_bypass~q ;
wire \A_ctrl_ld_st_bypass~q ;
wire \A_mem_bypass_pending~combout ;
wire \d_address_offset_field[0]~0_combout ;
wire \Add21~0_combout ;
wire \d_address_offset_field_nxt[2]~0_combout ;
wire \d_address_offset_field[0]~1_combout ;
wire \d_address_offset_field[0]~2_combout ;
wire \A_dc_wb_update_av_writedata~combout ;
wire \E_src2_reg[0]~q ;
wire \M_st_data[0]~q ;
wire \A_st_data[0]~q ;
wire \d_writedata_nxt[0]~0_combout ;
wire \d_writedata[14]~0_combout ;
wire \d_address_offset_field_nxt[0]~1_combout ;
wire \A_st_bypass_delayed~0_combout ;
wire \A_st_bypass_delayed~q ;
wire \A_st_bypass_delayed_started~0_combout ;
wire \A_st_bypass_delayed_started~q ;
wire \d_write_nxt~0_combout ;
wire \d_write_nxt~1_combout ;
wire \A_dc_wb_wr_want_dmaster~combout ;
wire \A_dc_wb_line[0]~q ;
wire \d_address_tag_field_nxt~0_combout ;
wire \d_address_line_field_nxt[0]~0_combout ;
wire \A_dc_actual_tag[1]~q ;
wire \A_dc_wb_tag[1]~q ;
wire \A_mem_baddr[12]~q ;
wire \d_address_tag_field_nxt[1]~1_combout ;
wire \A_dc_actual_tag[0]~q ;
wire \A_dc_wb_tag[0]~q ;
wire \A_mem_baddr[11]~q ;
wire \d_address_tag_field_nxt[0]~2_combout ;
wire \A_dc_wb_line[5]~q ;
wire \d_address_line_field_nxt[5]~1_combout ;
wire \A_dc_wb_line[4]~q ;
wire \d_address_line_field_nxt[4]~2_combout ;
wire \A_dc_wb_line[3]~q ;
wire \d_address_line_field_nxt[3]~3_combout ;
wire \A_dc_wb_line[2]~q ;
wire \d_address_line_field_nxt[2]~4_combout ;
wire \A_dc_wb_line[1]~q ;
wire \d_address_line_field_nxt[1]~5_combout ;
wire \A_dc_actual_tag[5]~q ;
wire \A_dc_wb_tag[5]~q ;
wire \A_mem_baddr[16]~q ;
wire \d_address_tag_field_nxt[5]~3_combout ;
wire \A_dc_actual_tag[4]~q ;
wire \A_dc_wb_tag[4]~q ;
wire \A_mem_baddr[15]~q ;
wire \d_address_tag_field_nxt[4]~4_combout ;
wire \A_dc_actual_tag[3]~q ;
wire \A_dc_wb_tag[3]~q ;
wire \A_mem_baddr[14]~q ;
wire \d_address_tag_field_nxt[3]~5_combout ;
wire \A_dc_actual_tag[2]~q ;
wire \A_dc_wb_tag[2]~q ;
wire \A_mem_baddr[13]~q ;
wire \d_address_tag_field_nxt[2]~6_combout ;
wire \d_address_offset_field_nxt[1]~2_combout ;
wire \A_ld_bypass_delayed~0_combout ;
wire \A_ld_bypass_delayed~q ;
wire \A_ld_bypass_delayed_started~0_combout ;
wire \A_ld_bypass_delayed_started~q ;
wire \d_read_nxt~0_combout ;
wire \d_read_nxt~1_combout ;
wire \A_dc_rd_addr_cnt_nxt[0]~3_combout ;
wire \A_dc_rd_addr_cnt[0]~0_combout ;
wire \A_dc_rd_addr_cnt[0]~q ;
wire \A_dc_rd_addr_cnt_nxt[1]~2_combout ;
wire \A_dc_rd_addr_cnt[1]~q ;
wire \A_dc_rd_addr_cnt_nxt[2]~1_combout ;
wire \A_dc_rd_addr_cnt[2]~q ;
wire \Add22~0_combout ;
wire \A_dc_rd_addr_cnt_nxt[3]~0_combout ;
wire \A_dc_rd_addr_cnt[3]~q ;
wire \d_read_nxt~2_combout ;
wire \F_ic_fill_same_tag_line~0_combout ;
wire \F_ic_fill_same_tag_line~1_combout ;
wire \F_ic_fill_same_tag_line~2_combout ;
wire \F_ic_fill_same_tag_line~3_combout ;
wire \F_ic_fill_same_tag_line~4_combout ;
wire \F_ic_fill_same_tag_line~5_combout ;
wire \F_ic_fill_same_tag_line~combout ;
wire \D_ic_fill_same_tag_line~q ;
wire \E_ctrl_invalidate_i~0_combout ;
wire \E_ctrl_invalidate_i~1_combout ;
wire \M_ctrl_invalidate_i~q ;
wire \ic_tag_clr_valid_bits_nxt~0_combout ;
wire \ic_fill_prevent_refill_nxt~combout ;
wire \ic_fill_prevent_refill~q ;
wire \ic_fill_initial_offset[2]~q ;
wire \D_ic_fill_starting_d1~q ;
wire \ic_fill_initial_offset[0]~q ;
wire \ic_fill_dp_offset_nxt[0]~1_combout ;
wire \i_readdatavalid_d1~q ;
wire \ic_fill_dp_offset_en~0_combout ;
wire \ic_fill_dp_offset[0]~q ;
wire \ic_fill_initial_offset[1]~q ;
wire \ic_fill_dp_offset_nxt[1]~2_combout ;
wire \ic_fill_dp_offset[1]~q ;
wire \ic_fill_dp_offset[2]~q ;
wire \ic_fill_dp_offset_nxt[2]~0_combout ;
wire \ic_fill_active_nxt~0_combout ;
wire \ic_fill_active_nxt~1_combout ;
wire \ic_fill_active~q ;
wire \D_ic_fill_starting~0_combout ;
wire \ic_fill_ap_cnt_nxt[0]~3_combout ;
wire \ic_fill_ap_cnt[3]~0_combout ;
wire \ic_fill_ap_cnt[0]~q ;
wire \ic_fill_ap_cnt_nxt[1]~2_combout ;
wire \ic_fill_ap_cnt[1]~q ;
wire \ic_fill_ap_cnt_nxt[2]~1_combout ;
wire \ic_fill_ap_cnt[2]~q ;
wire \ic_fill_ap_cnt_nxt[3]~0_combout ;
wire \ic_fill_ap_cnt[3]~q ;
wire \i_read_nxt~0_combout ;
wire \i_read_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~0_combout ;
wire \hbreak_enabled~0_combout ;
wire \ic_tag_wraddress_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~2_combout ;
wire \ic_tag_wraddress_nxt~3_combout ;
wire \ic_tag_wraddress_nxt~4_combout ;
wire \ic_tag_wraddress_nxt~5_combout ;
wire \ic_tag_wraddress_nxt~6_combout ;
wire \E_src2_reg[7]~q ;
wire \M_st_data[7]~q ;
wire \A_st_data[7]~q ;
wire \d_writedata_nxt[7]~1_combout ;
wire \ic_fill_ap_offset_nxt[0]~0_combout ;
wire \ic_fill_ap_offset_nxt[2]~1_combout ;
wire \ic_fill_ap_offset_nxt[1]~2_combout ;
wire \E_mem_byte_en~0_combout ;
wire \M_mem_byte_en[0]~q ;
wire \A_mem_byte_en[0]~q ;
wire \d_byteenable_nxt[0]~0_combout ;
wire \d_byteenable_nxt[0]~1_combout ;
wire \E_src2_reg[3]~q ;
wire \M_st_data[3]~q ;
wire \A_st_data[3]~q ;
wire \d_writedata_nxt[3]~2_combout ;
wire \E_src2_reg[1]~q ;
wire \M_st_data[1]~q ;
wire \A_st_data[1]~q ;
wire \d_writedata_nxt[1]~3_combout ;
wire \E_src2_reg[4]~q ;
wire \M_st_data[4]~q ;
wire \A_st_data[4]~q ;
wire \d_writedata_nxt[4]~4_combout ;
wire \E_src2_reg[20]~q ;
wire \M_st_data[20]~q ;
wire \A_st_data[20]~q ;
wire \d_writedata_nxt[20]~5_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \M_mem_byte_en[2]~q ;
wire \A_mem_byte_en[2]~q ;
wire \d_byteenable_nxt[2]~2_combout ;
wire \E_src2_reg[12]~q ;
wire \Equal0~0_combout ;
wire \M_st_data[12]~q ;
wire \A_st_data[12]~q ;
wire \d_writedata_nxt[12]~6_combout ;
wire \E_mem_byte_en[1]~2_combout ;
wire \M_mem_byte_en[1]~q ;
wire \A_mem_byte_en[1]~q ;
wire \d_byteenable_nxt[1]~3_combout ;
wire \D_src2_reg[28]~62_combout ;
wire \D_src2_reg[28]~63_combout ;
wire \E_src2_reg[28]~q ;
wire \E_st_data[28]~0_combout ;
wire \M_st_data[28]~q ;
wire \A_st_data[28]~q ;
wire \d_writedata_nxt[28]~7_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \M_mem_byte_en[3]~q ;
wire \A_mem_byte_en[3]~q ;
wire \d_byteenable_nxt[3]~4_combout ;
wire \D_src2_reg[16]~64_combout ;
wire \E_src2_reg[16]~q ;
wire \M_st_data[16]~q ;
wire \A_st_data[16]~q ;
wire \d_writedata_nxt[16]~8_combout ;
wire \E_src2_reg[8]~q ;
wire \M_st_data[8]~q ;
wire \A_st_data[8]~q ;
wire \d_writedata_nxt[8]~9_combout ;
wire \D_src2_reg[24]~65_combout ;
wire \D_src2_reg[24]~66_combout ;
wire \E_src2_reg[24]~q ;
wire \E_st_data[24]~1_combout ;
wire \M_st_data[24]~q ;
wire \A_st_data[24]~q ;
wire \d_writedata_nxt[24]~10_combout ;
wire \E_src2_reg[2]~q ;
wire \M_st_data[2]~q ;
wire \A_st_data[2]~q ;
wire \d_writedata_nxt[2]~11_combout ;
wire \D_src2_reg[18]~67_combout ;
wire \E_src2_reg[18]~q ;
wire \M_st_data[18]~q ;
wire \A_st_data[18]~q ;
wire \d_writedata_nxt[18]~12_combout ;
wire \E_src2_reg[10]~q ;
wire \M_st_data[10]~q ;
wire \A_st_data[10]~q ;
wire \d_writedata_nxt[10]~13_combout ;
wire \D_src2_reg[26]~68_combout ;
wire \D_src2_reg[26]~69_combout ;
wire \E_src2_reg[26]~q ;
wire \E_st_data[26]~2_combout ;
wire \M_st_data[26]~q ;
wire \A_st_data[26]~q ;
wire \d_writedata_nxt[26]~14_combout ;
wire \E_src2_reg[5]~q ;
wire \M_st_data[5]~q ;
wire \A_st_data[5]~q ;
wire \d_writedata_nxt[5]~15_combout ;
wire \D_src2_reg[21]~70_combout ;
wire \D_src2_reg[21]~71_combout ;
wire \E_src2_reg[21]~q ;
wire \M_st_data[21]~q ;
wire \A_st_data[21]~q ;
wire \d_writedata_nxt[21]~16_combout ;
wire \E_src2_reg[13]~q ;
wire \M_st_data[13]~q ;
wire \A_st_data[13]~q ;
wire \d_writedata_nxt[13]~17_combout ;
wire \D_src2_reg[29]~72_combout ;
wire \D_src2_reg[29]~73_combout ;
wire \E_src2_reg[29]~q ;
wire \E_st_data[29]~3_combout ;
wire \M_st_data[29]~q ;
wire \A_st_data[29]~q ;
wire \d_writedata_nxt[29]~18_combout ;
wire \D_src2_reg[23]~74_combout ;
wire \D_src2_reg[23]~75_combout ;
wire \E_src2_reg[23]~q ;
wire \M_st_data[23]~q ;
wire \A_st_data[23]~q ;
wire \d_writedata_nxt[23]~19_combout ;
wire \E_src2_reg[15]~q ;
wire \M_st_data[15]~q ;
wire \A_st_data[15]~q ;
wire \d_writedata_nxt[15]~20_combout ;
wire \D_src2_reg[31]~76_combout ;
wire \D_src2_reg[31]~77_combout ;
wire \E_src2_reg[31]~q ;
wire \E_st_data[31]~4_combout ;
wire \M_st_data[31]~q ;
wire \A_st_data[31]~q ;
wire \d_writedata_nxt[31]~21_combout ;
wire \E_src2_reg[11]~q ;
wire \M_st_data[11]~q ;
wire \A_st_data[11]~q ;
wire \d_writedata_nxt[11]~22_combout ;
wire \D_src2_reg[27]~78_combout ;
wire \D_src2_reg[27]~79_combout ;
wire \E_src2_reg[27]~q ;
wire \E_st_data[27]~5_combout ;
wire \M_st_data[27]~q ;
wire \A_st_data[27]~q ;
wire \d_writedata_nxt[27]~23_combout ;
wire \E_src2_reg[9]~q ;
wire \M_st_data[9]~q ;
wire \A_st_data[9]~q ;
wire \d_writedata_nxt[9]~24_combout ;
wire \D_src2_reg[25]~80_combout ;
wire \D_src2_reg[25]~81_combout ;
wire \E_src2_reg[25]~q ;
wire \E_st_data[25]~6_combout ;
wire \M_st_data[25]~q ;
wire \A_st_data[25]~q ;
wire \d_writedata_nxt[25]~25_combout ;
wire \E_src2_reg[6]~q ;
wire \M_st_data[6]~q ;
wire \A_st_data[6]~q ;
wire \d_writedata_nxt[6]~26_combout ;
wire \D_src2_reg[22]~82_combout ;
wire \D_src2_reg[22]~83_combout ;
wire \E_src2_reg[22]~q ;
wire \M_st_data[22]~q ;
wire \A_st_data[22]~q ;
wire \d_writedata_nxt[22]~27_combout ;
wire \E_src2_reg[14]~q ;
wire \M_st_data[14]~q ;
wire \A_st_data[14]~q ;
wire \d_writedata_nxt[14]~28_combout ;
wire \D_src2_reg[30]~84_combout ;
wire \D_src2_reg[30]~85_combout ;
wire \E_src2_reg[30]~q ;
wire \E_st_data[30]~7_combout ;
wire \M_st_data[30]~q ;
wire \A_st_data[30]~q ;
wire \d_writedata_nxt[30]~29_combout ;
wire \E_src2_reg[19]~q ;
wire \M_st_data[19]~q ;
wire \A_st_data[19]~q ;
wire \d_writedata_nxt[19]~30_combout ;
wire \D_src2_reg[17]~86_combout ;
wire \E_src2_reg[17]~q ;
wire \M_st_data[17]~q ;
wire \A_st_data[17]~q ;
wire \d_writedata_nxt[17]~31_combout ;


Qsys_system_Qsys_system_nios2_qsys_0_bht_module Qsys_system_nios2_qsys_0_bht(
	.q_b_1(\Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ),
	.F_stall(\F_stall~combout ),
	.M_bht_wr_en_unfiltered(\M_bht_wr_en_unfiltered~combout ),
	.M_bht_wr_data_unfiltered_1(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.M_bht_ptr_unfiltered_0(\M_bht_ptr_unfiltered[0]~q ),
	.M_bht_ptr_unfiltered_1(\M_bht_ptr_unfiltered[1]~q ),
	.M_bht_ptr_unfiltered_2(\M_bht_ptr_unfiltered[2]~q ),
	.M_bht_ptr_unfiltered_3(\M_bht_ptr_unfiltered[3]~q ),
	.M_bht_ptr_unfiltered_4(\M_bht_ptr_unfiltered[4]~q ),
	.M_bht_ptr_unfiltered_5(\M_bht_ptr_unfiltered[5]~q ),
	.M_bht_ptr_unfiltered_6(\M_bht_ptr_unfiltered[6]~q ),
	.M_bht_ptr_unfiltered_7(\M_bht_ptr_unfiltered[7]~q ),
	.F_bht_ptr_nxt_0(\F_bht_ptr_nxt[0]~combout ),
	.F_bht_ptr_nxt_1(\F_bht_ptr_nxt[1]~combout ),
	.F_bht_ptr_nxt_2(\F_bht_ptr_nxt[2]~combout ),
	.F_bht_ptr_nxt_3(\F_bht_ptr_nxt[3]~combout ),
	.F_bht_ptr_nxt_4(\F_bht_ptr_nxt[4]~combout ),
	.F_bht_ptr_nxt_5(\F_bht_ptr_nxt[5]~combout ),
	.F_bht_ptr_nxt_6(\F_bht_ptr_nxt[6]~combout ),
	.F_bht_ptr_nxt_7(\F_bht_ptr_nxt[7]~combout ),
	.M_br_mispredict(\M_br_mispredict~_wirecell_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_ic_tag_module Qsys_system_nios2_qsys_0_ic_tag(
	.q_b_2(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.ic_fill_valid_bits_5(\ic_fill_valid_bits[5]~q ),
	.ic_fill_valid_bits_7(\ic_fill_valid_bits[7]~q ),
	.ic_fill_valid_bits_4(\ic_fill_valid_bits[4]~q ),
	.q_b_6(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.ic_fill_valid_bits_6(\ic_fill_valid_bits[6]~q ),
	.ic_fill_valid_bits_1(\ic_fill_valid_bits[1]~q ),
	.ic_fill_valid_bits_3(\ic_fill_valid_bits[3]~q ),
	.ic_fill_valid_bits_0(\ic_fill_valid_bits[0]~q ),
	.ic_fill_valid_bits_2(\ic_fill_valid_bits[2]~q ),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.F_stall(\F_stall~combout ),
	.F_ic_tag_rd_addr_nxt_6(\F_ic_tag_rd_addr_nxt[6]~1_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~3_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~9_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~11_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~13_combout ),
	.ic_tag_wren(\ic_tag_wren~combout ),
	.ic_tag_wraddress_0(\ic_tag_wraddress[0]~q ),
	.ic_tag_wraddress_1(\ic_tag_wraddress[1]~q ),
	.ic_tag_wraddress_2(\ic_tag_wraddress[2]~q ),
	.ic_tag_wraddress_3(\ic_tag_wraddress[3]~q ),
	.ic_tag_wraddress_4(\ic_tag_wraddress[4]~q ),
	.ic_tag_wraddress_5(\ic_tag_wraddress[5]~q ),
	.ic_tag_wraddress_6(\ic_tag_wraddress[6]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_dc_tag_module Qsys_system_nios2_qsys_0_dc_tag(
	.q_b_4(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[7] ),
	.dc_tag_wr_port_en(\dc_tag_wr_port_en~combout ),
	.dc_tag_wr_port_data_4(\dc_tag_wr_port_data[4]~1_combout ),
	.dc_tag_wr_port_addr_0(\dc_tag_wr_port_addr[0]~0_combout ),
	.dc_tag_wr_port_addr_1(\dc_tag_wr_port_addr[1]~1_combout ),
	.dc_tag_wr_port_addr_2(\dc_tag_wr_port_addr[2]~2_combout ),
	.dc_tag_wr_port_addr_3(\dc_tag_wr_port_addr[3]~3_combout ),
	.dc_tag_wr_port_addr_4(\dc_tag_wr_port_addr[4]~4_combout ),
	.dc_tag_wr_port_addr_5(\dc_tag_wr_port_addr[5]~5_combout ),
	.dc_tag_rd_port_addr_0(\dc_tag_rd_port_addr[0]~0_combout ),
	.dc_tag_rd_port_addr_1(\dc_tag_rd_port_addr[1]~1_combout ),
	.dc_tag_rd_port_addr_2(\dc_tag_rd_port_addr[2]~2_combout ),
	.dc_tag_rd_port_addr_3(\dc_tag_rd_port_addr[3]~3_combout ),
	.dc_tag_rd_port_addr_4(\dc_tag_rd_port_addr[4]~4_combout ),
	.dc_tag_rd_port_addr_5(\dc_tag_rd_port_addr[5]~5_combout ),
	.dc_tag_wr_port_data_5(\dc_tag_wr_port_data[5]~2_combout ),
	.dc_tag_wr_port_data_6(\dc_tag_wr_port_data[6]~3_combout ),
	.dc_tag_wr_port_data_0(\dc_tag_wr_port_data[0]~4_combout ),
	.dc_tag_wr_port_data_1(\dc_tag_wr_port_data[1]~5_combout ),
	.dc_tag_wr_port_data_2(\dc_tag_wr_port_data[2]~6_combout ),
	.dc_tag_wr_port_data_3(\dc_tag_wr_port_data[3]~7_combout ),
	.dc_tag_wr_port_data_7(\dc_tag_wr_port_data[7]~8_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_register_bank_b_module Qsys_system_nios2_qsys_0_register_bank_b(
	.q_b_4(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_16(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_29(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_30(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_26(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_19(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_17(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_22(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_18(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_24(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_31(\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~3_combout ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~5_combout ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~7_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~9_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~13_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~15_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~17_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~19_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~21_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~23_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~25_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~28_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~30_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~32_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~34_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~36_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~38_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~40_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~42_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~44_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~46_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~48_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~50_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~52_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~54_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~56_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~58_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~60_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~62_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~64_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~66_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~68_combout ),
	.A_dst_regnum_from_M_4(\A_dst_regnum_from_M[4]~q ),
	.A_wr_dst_reg_from_M(\A_wr_dst_reg_from_M~q ),
	.A_dst_regnum_from_M_0(\A_dst_regnum_from_M[0]~q ),
	.A_dst_regnum_from_M_1(\A_dst_regnum_from_M[1]~q ),
	.A_dst_regnum_from_M_2(\A_dst_regnum_from_M[2]~q ),
	.A_dst_regnum_from_M_3(\A_dst_regnum_from_M[3]~q ),
	.rf_b_rd_port_addr_0(\rf_b_rd_port_addr[0]~0_combout ),
	.rf_b_rd_port_addr_1(\rf_b_rd_port_addr[1]~1_combout ),
	.rf_b_rd_port_addr_2(\rf_b_rd_port_addr[2]~2_combout ),
	.rf_b_rd_port_addr_3(\rf_b_rd_port_addr[3]~3_combout ),
	.rf_b_rd_port_addr_4(\rf_b_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_register_bank_a_module Qsys_system_nios2_qsys_0_register_bank_a(
	.q_b_4(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_16(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_29(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_30(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_26(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_19(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_17(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_22(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_18(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_24(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_31(\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~3_combout ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~5_combout ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~7_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~9_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~13_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~15_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~17_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~19_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~21_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~23_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~25_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~28_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~30_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~32_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~34_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~36_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~38_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~40_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~42_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~44_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~46_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~48_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~50_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~52_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~54_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~56_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~58_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~60_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~62_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~64_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~66_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~68_combout ),
	.A_dst_regnum_from_M_4(\A_dst_regnum_from_M[4]~q ),
	.A_wr_dst_reg_from_M(\A_wr_dst_reg_from_M~q ),
	.A_dst_regnum_from_M_0(\A_dst_regnum_from_M[0]~q ),
	.A_dst_regnum_from_M_1(\A_dst_regnum_from_M[1]~q ),
	.A_dst_regnum_from_M_2(\A_dst_regnum_from_M[2]~q ),
	.A_dst_regnum_from_M_3(\A_dst_regnum_from_M[3]~q ),
	.rf_a_rd_port_addr_0(\rf_a_rd_port_addr[0]~0_combout ),
	.rf_a_rd_port_addr_1(\rf_a_rd_port_addr[1]~1_combout ),
	.rf_a_rd_port_addr_2(\rf_a_rd_port_addr[2]~2_combout ),
	.rf_a_rd_port_addr_3(\rf_a_rd_port_addr[3]~3_combout ),
	.rf_a_rd_port_addr_4(\rf_a_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_dc_victim_module Qsys_system_nios2_qsys_0_dc_victim(
	.q_b_0(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ),
	.A_dc_xfer_wr_data_0(\A_dc_xfer_wr_data[0]~q ),
	.q_b_7(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ),
	.A_dc_xfer_wr_data_7(\A_dc_xfer_wr_data[7]~q ),
	.q_b_1(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ),
	.A_dc_xfer_wr_data_3(\A_dc_xfer_wr_data[3]~q ),
	.q_b_4(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_20(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_28(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_16(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_24(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_18(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_26(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_21(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_13(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_29(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_23(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_15(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_31(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_27(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_25(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_22(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_30(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_19(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ),
	.A_dc_xfer_wr_data_1(\A_dc_xfer_wr_data[1]~q ),
	.q_b_17(\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ),
	.A_dc_xfer_wr_data_4(\A_dc_xfer_wr_data[4]~q ),
	.A_dc_xfer_wr_data_20(\A_dc_xfer_wr_data[20]~q ),
	.A_dc_xfer_wr_data_12(\A_dc_xfer_wr_data[12]~q ),
	.A_dc_xfer_wr_data_28(\A_dc_xfer_wr_data[28]~q ),
	.A_dc_xfer_wr_data_16(\A_dc_xfer_wr_data[16]~q ),
	.A_dc_xfer_wr_data_8(\A_dc_xfer_wr_data[8]~q ),
	.A_dc_xfer_wr_data_24(\A_dc_xfer_wr_data[24]~q ),
	.A_dc_xfer_wr_data_2(\A_dc_xfer_wr_data[2]~q ),
	.A_dc_xfer_wr_data_18(\A_dc_xfer_wr_data[18]~q ),
	.A_dc_xfer_wr_data_10(\A_dc_xfer_wr_data[10]~q ),
	.A_dc_xfer_wr_data_26(\A_dc_xfer_wr_data[26]~q ),
	.A_dc_xfer_wr_data_5(\A_dc_xfer_wr_data[5]~q ),
	.A_dc_xfer_wr_data_21(\A_dc_xfer_wr_data[21]~q ),
	.A_dc_xfer_wr_data_13(\A_dc_xfer_wr_data[13]~q ),
	.A_dc_xfer_wr_data_29(\A_dc_xfer_wr_data[29]~q ),
	.A_dc_xfer_wr_data_23(\A_dc_xfer_wr_data[23]~q ),
	.A_dc_xfer_wr_data_15(\A_dc_xfer_wr_data[15]~q ),
	.A_dc_xfer_wr_data_31(\A_dc_xfer_wr_data[31]~q ),
	.A_dc_xfer_wr_data_11(\A_dc_xfer_wr_data[11]~q ),
	.A_dc_xfer_wr_data_27(\A_dc_xfer_wr_data[27]~q ),
	.A_dc_xfer_wr_data_9(\A_dc_xfer_wr_data[9]~q ),
	.A_dc_xfer_wr_data_25(\A_dc_xfer_wr_data[25]~q ),
	.A_dc_xfer_wr_data_6(\A_dc_xfer_wr_data[6]~q ),
	.A_dc_xfer_wr_data_22(\A_dc_xfer_wr_data[22]~q ),
	.A_dc_xfer_wr_data_14(\A_dc_xfer_wr_data[14]~q ),
	.A_dc_xfer_wr_data_30(\A_dc_xfer_wr_data[30]~q ),
	.A_dc_xfer_wr_data_19(\A_dc_xfer_wr_data[19]~q ),
	.A_dc_xfer_wr_data_17(\A_dc_xfer_wr_data[17]~q ),
	.A_dc_xfer_wr_active(\A_dc_xfer_wr_active~q ),
	.A_dc_wb_rd_en(\A_dc_wb_rd_en~combout ),
	.A_dc_xfer_wr_offset_0(\A_dc_xfer_wr_offset[0]~q ),
	.A_dc_xfer_wr_offset_1(\A_dc_xfer_wr_offset[1]~q ),
	.A_dc_xfer_wr_offset_2(\A_dc_xfer_wr_offset[2]~q ),
	.A_dc_wb_rd_addr_offset_0(\A_dc_wb_rd_addr_offset[0]~q ),
	.A_dc_wb_rd_addr_offset_1(\A_dc_wb_rd_addr_offset[1]~q ),
	.A_dc_wb_rd_addr_offset_2(\A_dc_wb_rd_addr_offset[2]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_dc_data_module Qsys_system_nios2_qsys_0_dc_data(
	.q_b_0(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_4(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_20(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_28(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_16(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_24(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_18(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_26(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_5(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_21(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_13(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_29(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_23(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_15(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_31(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_27(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_25(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_22(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_30(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_19(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_17(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.dc_data_wr_port_en(\dc_data_wr_port_en~combout ),
	.dc_data_wr_port_data_0(\dc_data_wr_port_data[0]~1_combout ),
	.dc_data_wr_port_addr_0(\dc_data_wr_port_addr[0]~0_combout ),
	.dc_data_wr_port_addr_1(\dc_data_wr_port_addr[1]~1_combout ),
	.dc_data_wr_port_addr_2(\dc_data_wr_port_addr[2]~2_combout ),
	.dc_data_wr_port_addr_3(\dc_data_wr_port_addr[3]~3_combout ),
	.dc_data_wr_port_addr_4(\dc_data_wr_port_addr[4]~4_combout ),
	.dc_data_wr_port_addr_5(\dc_data_wr_port_addr[5]~5_combout ),
	.dc_data_wr_port_addr_6(\dc_data_wr_port_addr[6]~6_combout ),
	.dc_data_wr_port_addr_7(\dc_data_wr_port_addr[7]~7_combout ),
	.dc_data_wr_port_addr_8(\dc_data_wr_port_addr[8]~8_combout ),
	.dc_data_rd_port_addr_0(\dc_data_rd_port_addr[0]~0_combout ),
	.dc_data_rd_port_addr_1(\dc_data_rd_port_addr[1]~1_combout ),
	.dc_data_rd_port_addr_2(\dc_data_rd_port_addr[2]~2_combout ),
	.dc_data_rd_port_addr_3(\dc_data_rd_port_addr[3]~3_combout ),
	.dc_data_rd_port_addr_4(\dc_data_rd_port_addr[4]~4_combout ),
	.dc_data_rd_port_addr_5(\dc_data_rd_port_addr[5]~5_combout ),
	.dc_data_rd_port_addr_6(\dc_data_rd_port_addr[6]~6_combout ),
	.dc_data_rd_port_addr_7(\dc_data_rd_port_addr[7]~7_combout ),
	.dc_data_rd_port_addr_8(\dc_data_rd_port_addr[8]~8_combout ),
	.dc_data_wr_port_data_4(\dc_data_wr_port_data[4]~2_combout ),
	.dc_data_wr_port_data_20(\dc_data_wr_port_data[20]~4_combout ),
	.dc_data_wr_port_data_12(\dc_data_wr_port_data[12]~6_combout ),
	.dc_data_wr_port_data_28(\dc_data_wr_port_data[28]~8_combout ),
	.dc_data_wr_port_data_16(\dc_data_wr_port_data[16]~9_combout ),
	.dc_data_wr_port_data_8(\dc_data_wr_port_data[8]~10_combout ),
	.dc_data_wr_port_data_24(\dc_data_wr_port_data[24]~11_combout ),
	.dc_data_wr_port_data_2(\dc_data_wr_port_data[2]~12_combout ),
	.dc_data_wr_port_data_18(\dc_data_wr_port_data[18]~13_combout ),
	.dc_data_wr_port_data_10(\dc_data_wr_port_data[10]~14_combout ),
	.dc_data_wr_port_data_26(\dc_data_wr_port_data[26]~15_combout ),
	.dc_data_wr_port_data_5(\dc_data_wr_port_data[5]~16_combout ),
	.dc_data_wr_port_data_21(\dc_data_wr_port_data[21]~17_combout ),
	.dc_data_wr_port_data_13(\dc_data_wr_port_data[13]~18_combout ),
	.dc_data_wr_port_data_29(\dc_data_wr_port_data[29]~19_combout ),
	.dc_data_wr_port_data_7(\dc_data_wr_port_data[7]~20_combout ),
	.dc_data_wr_port_data_23(\dc_data_wr_port_data[23]~21_combout ),
	.dc_data_wr_port_data_15(\dc_data_wr_port_data[15]~22_combout ),
	.dc_data_wr_port_data_31(\dc_data_wr_port_data[31]~23_combout ),
	.dc_data_wr_port_data_11(\dc_data_wr_port_data[11]~24_combout ),
	.dc_data_wr_port_data_27(\dc_data_wr_port_data[27]~25_combout ),
	.dc_data_wr_port_data_9(\dc_data_wr_port_data[9]~26_combout ),
	.dc_data_wr_port_data_25(\dc_data_wr_port_data[25]~27_combout ),
	.dc_data_wr_port_data_6(\dc_data_wr_port_data[6]~28_combout ),
	.dc_data_wr_port_data_22(\dc_data_wr_port_data[22]~29_combout ),
	.dc_data_wr_port_data_14(\dc_data_wr_port_data[14]~30_combout ),
	.dc_data_wr_port_data_30(\dc_data_wr_port_data[30]~31_combout ),
	.dc_data_wr_port_data_3(\dc_data_wr_port_data[3]~32_combout ),
	.dc_data_wr_port_data_19(\dc_data_wr_port_data[19]~33_combout ),
	.dc_data_wr_port_data_1(\dc_data_wr_port_data[1]~34_combout ),
	.dc_data_wr_port_data_17(\dc_data_wr_port_data[17]~35_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_ic_data_module Qsys_system_nios2_qsys_0_ic_data(
	.q_b_5(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_3(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_1(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_4(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_2(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_28(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_30(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_27(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_29(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_0(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_23(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_25(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_26(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_22(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_24(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_16(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_13(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_12(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_8(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_18(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_21(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_6(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_20(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_9(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_7(\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.ic_fill_line_6(ic_fill_line_6),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_0(ic_fill_line_0),
	.F_stall(\F_stall~combout ),
	.ic_fill_dp_offset_0(\ic_fill_dp_offset[0]~q ),
	.ic_fill_dp_offset_1(\ic_fill_dp_offset[1]~q ),
	.ic_fill_dp_offset_2(\ic_fill_dp_offset[2]~q ),
	.i_readdatavalid_d1(\i_readdatavalid_d1~q ),
	.F_ic_tag_rd_addr_nxt_6(\F_ic_tag_rd_addr_nxt[6]~1_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~3_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~9_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~11_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~13_combout ),
	.i_readdata_d1_5(\i_readdata_d1[5]~q ),
	.F_ic_data_rd_addr_nxt_0(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.F_ic_data_rd_addr_nxt_1(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.F_ic_data_rd_addr_nxt_2(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.i_readdata_d1_3(\i_readdata_d1[3]~q ),
	.i_readdata_d1_1(\i_readdata_d1[1]~q ),
	.i_readdata_d1_4(\i_readdata_d1[4]~q ),
	.i_readdata_d1_2(\i_readdata_d1[2]~q ),
	.i_readdata_d1_28(\i_readdata_d1[28]~q ),
	.i_readdata_d1_30(\i_readdata_d1[30]~q ),
	.i_readdata_d1_31(\i_readdata_d1[31]~q ),
	.i_readdata_d1_27(\i_readdata_d1[27]~q ),
	.i_readdata_d1_29(\i_readdata_d1[29]~q ),
	.i_readdata_d1_0(\i_readdata_d1[0]~q ),
	.i_readdata_d1_23(\i_readdata_d1[23]~q ),
	.i_readdata_d1_25(\i_readdata_d1[25]~q ),
	.i_readdata_d1_26(\i_readdata_d1[26]~q ),
	.i_readdata_d1_22(\i_readdata_d1[22]~q ),
	.i_readdata_d1_24(\i_readdata_d1[24]~q ),
	.i_readdata_d1_16(\i_readdata_d1[16]~q ),
	.i_readdata_d1_15(\i_readdata_d1[15]~q ),
	.i_readdata_d1_13(\i_readdata_d1[13]~q ),
	.i_readdata_d1_14(\i_readdata_d1[14]~q ),
	.i_readdata_d1_12(\i_readdata_d1[12]~q ),
	.i_readdata_d1_11(\i_readdata_d1[11]~q ),
	.i_readdata_d1_10(\i_readdata_d1[10]~q ),
	.i_readdata_d1_8(\i_readdata_d1[8]~q ),
	.i_readdata_d1_18(\i_readdata_d1[18]~q ),
	.i_readdata_d1_17(\i_readdata_d1[17]~q ),
	.i_readdata_d1_21(\i_readdata_d1[21]~q ),
	.i_readdata_d1_6(\i_readdata_d1[6]~q ),
	.i_readdata_d1_20(\i_readdata_d1[20]~q ),
	.i_readdata_d1_19(\i_readdata_d1[19]~q ),
	.i_readdata_d1_9(\i_readdata_d1[9]~q ),
	.i_readdata_d1_7(\i_readdata_d1[7]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_mult_cell the_Qsys_system_nios2_qsys_0_mult_cell(
	.Add0(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~1_sumout ),
	.Add01(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~5_sumout ),
	.Add02(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~9_sumout ),
	.Add03(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~13_sumout ),
	.Add04(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~17_sumout ),
	.Add05(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~21_sumout ),
	.Add06(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~25_sumout ),
	.Add07(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~29_sumout ),
	.Add08(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~33_sumout ),
	.Add09(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~37_sumout ),
	.Add010(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~41_sumout ),
	.Add011(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~45_sumout ),
	.Add012(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~49_sumout ),
	.Add013(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~53_sumout ),
	.Add014(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~57_sumout ),
	.Add015(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~61_sumout ),
	.A_mul_src2_0(\A_mul_src2[0]~q ),
	.A_mul_src2_1(\A_mul_src2[1]~q ),
	.A_mul_src2_2(\A_mul_src2[2]~q ),
	.A_mul_src2_3(\A_mul_src2[3]~q ),
	.A_mul_src2_4(\A_mul_src2[4]~q ),
	.A_mul_src2_5(\A_mul_src2[5]~q ),
	.A_mul_src2_6(\A_mul_src2[6]~q ),
	.A_mul_src2_7(\A_mul_src2[7]~q ),
	.A_mul_src2_8(\A_mul_src2[8]~q ),
	.A_mul_src2_9(\A_mul_src2[9]~q ),
	.A_mul_src2_10(\A_mul_src2[10]~q ),
	.A_mul_src2_11(\A_mul_src2[11]~q ),
	.A_mul_src2_12(\A_mul_src2[12]~q ),
	.A_mul_src2_13(\A_mul_src2[13]~q ),
	.A_mul_src2_14(\A_mul_src2[14]~q ),
	.A_mul_src2_15(\A_mul_src2[15]~q ),
	.A_mul_src1_0(\A_mul_src1[0]~q ),
	.A_mul_src1_1(\A_mul_src1[1]~q ),
	.A_mul_src1_2(\A_mul_src1[2]~q ),
	.A_mul_src1_3(\A_mul_src1[3]~q ),
	.A_mul_src1_4(\A_mul_src1[4]~q ),
	.A_mul_src1_5(\A_mul_src1[5]~q ),
	.A_mul_src1_6(\A_mul_src1[6]~q ),
	.A_mul_src1_7(\A_mul_src1[7]~q ),
	.A_mul_src1_8(\A_mul_src1[8]~q ),
	.A_mul_src1_9(\A_mul_src1[9]~q ),
	.A_mul_src1_10(\A_mul_src1[10]~q ),
	.A_mul_src1_11(\A_mul_src1[11]~q ),
	.A_mul_src1_12(\A_mul_src1[12]~q ),
	.A_mul_src1_13(\A_mul_src1[13]~q ),
	.A_mul_src1_14(\A_mul_src1[14]~q ),
	.A_mul_src1_15(\A_mul_src1[15]~q ),
	.A_mul_src1_16(\A_mul_src1[16]~q ),
	.A_mul_src1_17(\A_mul_src1[17]~q ),
	.A_mul_src1_18(\A_mul_src1[18]~q ),
	.A_mul_src1_19(\A_mul_src1[19]~q ),
	.A_mul_src1_20(\A_mul_src1[20]~q ),
	.A_mul_src1_21(\A_mul_src1[21]~q ),
	.A_mul_src1_22(\A_mul_src1[22]~q ),
	.A_mul_src1_23(\A_mul_src1[23]~q ),
	.A_mul_src1_24(\A_mul_src1[24]~q ),
	.A_mul_src1_25(\A_mul_src1[25]~q ),
	.A_mul_src1_26(\A_mul_src1[26]~q ),
	.A_mul_src1_27(\A_mul_src1[27]~q ),
	.A_mul_src1_28(\A_mul_src1[28]~q ),
	.A_mul_src1_29(\A_mul_src1[29]~q ),
	.A_mul_src1_30(\A_mul_src1[30]~q ),
	.A_mul_src1_31(\A_mul_src1[31]~q ),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_4(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_0(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_2(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_5(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_12(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_11(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_10(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_9(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_8(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_7(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_6(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_15(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_14(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_13(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_3(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_1(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci the_Qsys_system_nios2_qsys_0_nios2_oci(
	.readdata_4(readdata_4),
	.readdata_20(readdata_20),
	.readdata_12(readdata_12),
	.readdata_28(readdata_28),
	.readdata_16(readdata_16),
	.readdata_8(readdata_8),
	.readdata_24(readdata_24),
	.readdata_2(readdata_2),
	.readdata_18(readdata_18),
	.readdata_10(readdata_10),
	.readdata_26(readdata_26),
	.readdata_5(readdata_5),
	.readdata_21(readdata_21),
	.readdata_13(readdata_13),
	.readdata_29(readdata_29),
	.readdata_7(readdata_7),
	.readdata_23(readdata_23),
	.readdata_15(readdata_15),
	.readdata_31(readdata_31),
	.readdata_11(readdata_11),
	.readdata_27(readdata_27),
	.readdata_9(readdata_9),
	.readdata_25(readdata_25),
	.readdata_6(readdata_6),
	.readdata_22(readdata_22),
	.readdata_14(readdata_14),
	.readdata_30(readdata_30),
	.readdata_3(readdata_3),
	.readdata_19(readdata_19),
	.readdata_17(readdata_17),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_write(d_write1),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.waitrequest(jtag_debug_module_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr1),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled(hbreak_enabled1),
	.jtag_break(\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.oci_single_step_mode(\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ),
	.r_early_rst(r_early_rst),
	.writedata_nxt({src_payload26,src_payload32,src_payload22,src_payload17,src_payload11,src_payload10,src_payload12,src_payload8,src_payload24,src_payload30,src_payload14,src_payload6,src_payload7,src_payload15,src_payload13,src_payload5,src_payload25,src_payload31,src_payload21,src_payload16,
src_payload27,src_payload19,src_payload28,src_payload18,src_payload23,src_payload29,src_payload20,src_payload9,src_payload2,src_payload4,src_payload3,src_payload}),
	.debugaccess_nxt(src_payload1),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.oci_ienable_0(\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_ienable_1(\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[1]~q ),
	.readdata_0(readdata_0),
	.resetrequest(jtag_debug_module_resetrequest),
	.readdata_1(readdata_1),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

dffeas \A_dc_xfer_wr_data[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[0]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[0] .power_up = "low";

dffeas \ic_fill_valid_bits[5] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[5]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[5] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[5] .power_up = "low";

dffeas \ic_fill_valid_bits[7] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[7]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[7] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[7] .power_up = "low";

dffeas \ic_fill_valid_bits[4] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[4]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[4] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[4] .power_up = "low";

dffeas \ic_fill_valid_bits[6] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[6]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[6] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[6] .power_up = "low";

dffeas \A_dc_xfer_wr_data[7] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[7]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[7]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[7] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[7] .power_up = "low";

dffeas \ic_fill_valid_bits[1] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[1]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[1] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[1] .power_up = "low";

dffeas \ic_fill_valid_bits[3] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[3]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[3] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[3] .power_up = "low";

dffeas \ic_fill_valid_bits[0] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[0]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[0] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[0] .power_up = "low";

dffeas \ic_fill_valid_bits[2] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[2]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[2] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[2] .power_up = "low";

dffeas \A_dc_xfer_wr_data[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[3]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[3]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[3] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[3] .power_up = "low";

dffeas \A_mul_src2[0] (
	.clk(clk_clk),
	.d(\M_div_src2[0]~q ),
	.asdata(\A_mul_src2[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[0]~q ),
	.prn(vcc));
defparam \A_mul_src2[0] .is_wysiwyg = "true";
defparam \A_mul_src2[0] .power_up = "low";

dffeas \A_mul_src2[1] (
	.clk(clk_clk),
	.d(\M_div_src2[1]~q ),
	.asdata(\A_mul_src2[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[1]~q ),
	.prn(vcc));
defparam \A_mul_src2[1] .is_wysiwyg = "true";
defparam \A_mul_src2[1] .power_up = "low";

dffeas \A_mul_src2[2] (
	.clk(clk_clk),
	.d(\M_div_src2[2]~q ),
	.asdata(\A_mul_src2[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[2]~q ),
	.prn(vcc));
defparam \A_mul_src2[2] .is_wysiwyg = "true";
defparam \A_mul_src2[2] .power_up = "low";

dffeas \A_mul_src2[3] (
	.clk(clk_clk),
	.d(\M_div_src2[3]~q ),
	.asdata(\A_mul_src2[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[3]~q ),
	.prn(vcc));
defparam \A_mul_src2[3] .is_wysiwyg = "true";
defparam \A_mul_src2[3] .power_up = "low";

dffeas \A_mul_src2[4] (
	.clk(clk_clk),
	.d(\M_div_src2[4]~q ),
	.asdata(\A_mul_src2[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[4]~q ),
	.prn(vcc));
defparam \A_mul_src2[4] .is_wysiwyg = "true";
defparam \A_mul_src2[4] .power_up = "low";

dffeas \A_mul_src2[5] (
	.clk(clk_clk),
	.d(\M_div_src2[5]~q ),
	.asdata(\A_mul_src2[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[5]~q ),
	.prn(vcc));
defparam \A_mul_src2[5] .is_wysiwyg = "true";
defparam \A_mul_src2[5] .power_up = "low";

dffeas \A_mul_src2[6] (
	.clk(clk_clk),
	.d(\M_div_src2[6]~q ),
	.asdata(\A_mul_src2[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[6]~q ),
	.prn(vcc));
defparam \A_mul_src2[6] .is_wysiwyg = "true";
defparam \A_mul_src2[6] .power_up = "low";

dffeas \A_mul_src2[7] (
	.clk(clk_clk),
	.d(\M_div_src2[7]~q ),
	.asdata(\A_mul_src2[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[7]~q ),
	.prn(vcc));
defparam \A_mul_src2[7] .is_wysiwyg = "true";
defparam \A_mul_src2[7] .power_up = "low";

dffeas \A_mul_src2[8] (
	.clk(clk_clk),
	.d(\M_div_src2[8]~q ),
	.asdata(\A_mul_src2[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[8]~q ),
	.prn(vcc));
defparam \A_mul_src2[8] .is_wysiwyg = "true";
defparam \A_mul_src2[8] .power_up = "low";

dffeas \A_mul_src2[9] (
	.clk(clk_clk),
	.d(\M_div_src2[9]~q ),
	.asdata(\A_mul_src2[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[9]~q ),
	.prn(vcc));
defparam \A_mul_src2[9] .is_wysiwyg = "true";
defparam \A_mul_src2[9] .power_up = "low";

dffeas \A_mul_src2[10] (
	.clk(clk_clk),
	.d(\M_div_src2[10]~q ),
	.asdata(\A_mul_src2[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[10]~q ),
	.prn(vcc));
defparam \A_mul_src2[10] .is_wysiwyg = "true";
defparam \A_mul_src2[10] .power_up = "low";

dffeas \A_mul_src2[11] (
	.clk(clk_clk),
	.d(\M_div_src2[11]~q ),
	.asdata(\A_mul_src2[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[11]~q ),
	.prn(vcc));
defparam \A_mul_src2[11] .is_wysiwyg = "true";
defparam \A_mul_src2[11] .power_up = "low";

dffeas \A_mul_src2[12] (
	.clk(clk_clk),
	.d(\M_div_src2[12]~q ),
	.asdata(\A_mul_src2[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[12]~q ),
	.prn(vcc));
defparam \A_mul_src2[12] .is_wysiwyg = "true";
defparam \A_mul_src2[12] .power_up = "low";

dffeas \A_mul_src2[13] (
	.clk(clk_clk),
	.d(\M_div_src2[13]~q ),
	.asdata(\A_mul_src2[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[13]~q ),
	.prn(vcc));
defparam \A_mul_src2[13] .is_wysiwyg = "true";
defparam \A_mul_src2[13] .power_up = "low";

dffeas \A_mul_src2[14] (
	.clk(clk_clk),
	.d(\M_div_src2[14]~q ),
	.asdata(\A_mul_src2[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[14]~q ),
	.prn(vcc));
defparam \A_mul_src2[14] .is_wysiwyg = "true";
defparam \A_mul_src2[14] .power_up = "low";

dffeas \A_mul_src2[15] (
	.clk(clk_clk),
	.d(\M_div_src2[15]~q ),
	.asdata(\A_mul_src2[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[15]~q ),
	.prn(vcc));
defparam \A_mul_src2[15] .is_wysiwyg = "true";
defparam \A_mul_src2[15] .power_up = "low";

dffeas \A_mul_src1[0] (
	.clk(clk_clk),
	.d(\M_div_src1[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[0]~q ),
	.prn(vcc));
defparam \A_mul_src1[0] .is_wysiwyg = "true";
defparam \A_mul_src1[0] .power_up = "low";

dffeas \A_mul_src1[1] (
	.clk(clk_clk),
	.d(\M_div_src1[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[1]~q ),
	.prn(vcc));
defparam \A_mul_src1[1] .is_wysiwyg = "true";
defparam \A_mul_src1[1] .power_up = "low";

dffeas \A_mul_src1[2] (
	.clk(clk_clk),
	.d(\M_div_src1[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[2]~q ),
	.prn(vcc));
defparam \A_mul_src1[2] .is_wysiwyg = "true";
defparam \A_mul_src1[2] .power_up = "low";

dffeas \A_mul_src1[3] (
	.clk(clk_clk),
	.d(\M_div_src1[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[3]~q ),
	.prn(vcc));
defparam \A_mul_src1[3] .is_wysiwyg = "true";
defparam \A_mul_src1[3] .power_up = "low";

dffeas \A_mul_src1[4] (
	.clk(clk_clk),
	.d(\M_div_src1[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[4]~q ),
	.prn(vcc));
defparam \A_mul_src1[4] .is_wysiwyg = "true";
defparam \A_mul_src1[4] .power_up = "low";

dffeas \A_mul_src1[5] (
	.clk(clk_clk),
	.d(\M_div_src1[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[5]~q ),
	.prn(vcc));
defparam \A_mul_src1[5] .is_wysiwyg = "true";
defparam \A_mul_src1[5] .power_up = "low";

dffeas \A_mul_src1[6] (
	.clk(clk_clk),
	.d(\M_div_src1[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[6]~q ),
	.prn(vcc));
defparam \A_mul_src1[6] .is_wysiwyg = "true";
defparam \A_mul_src1[6] .power_up = "low";

dffeas \A_mul_src1[7] (
	.clk(clk_clk),
	.d(\M_div_src1[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[7]~q ),
	.prn(vcc));
defparam \A_mul_src1[7] .is_wysiwyg = "true";
defparam \A_mul_src1[7] .power_up = "low";

dffeas \A_mul_src1[8] (
	.clk(clk_clk),
	.d(\M_div_src1[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[8]~q ),
	.prn(vcc));
defparam \A_mul_src1[8] .is_wysiwyg = "true";
defparam \A_mul_src1[8] .power_up = "low";

dffeas \A_mul_src1[9] (
	.clk(clk_clk),
	.d(\M_div_src1[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[9]~q ),
	.prn(vcc));
defparam \A_mul_src1[9] .is_wysiwyg = "true";
defparam \A_mul_src1[9] .power_up = "low";

dffeas \A_mul_src1[10] (
	.clk(clk_clk),
	.d(\M_div_src1[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[10]~q ),
	.prn(vcc));
defparam \A_mul_src1[10] .is_wysiwyg = "true";
defparam \A_mul_src1[10] .power_up = "low";

dffeas \A_mul_src1[11] (
	.clk(clk_clk),
	.d(\M_div_src1[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[11]~q ),
	.prn(vcc));
defparam \A_mul_src1[11] .is_wysiwyg = "true";
defparam \A_mul_src1[11] .power_up = "low";

dffeas \A_mul_src1[12] (
	.clk(clk_clk),
	.d(\M_div_src1[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[12]~q ),
	.prn(vcc));
defparam \A_mul_src1[12] .is_wysiwyg = "true";
defparam \A_mul_src1[12] .power_up = "low";

dffeas \A_mul_src1[13] (
	.clk(clk_clk),
	.d(\M_div_src1[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[13]~q ),
	.prn(vcc));
defparam \A_mul_src1[13] .is_wysiwyg = "true";
defparam \A_mul_src1[13] .power_up = "low";

dffeas \A_mul_src1[14] (
	.clk(clk_clk),
	.d(\M_div_src1[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[14]~q ),
	.prn(vcc));
defparam \A_mul_src1[14] .is_wysiwyg = "true";
defparam \A_mul_src1[14] .power_up = "low";

dffeas \A_mul_src1[15] (
	.clk(clk_clk),
	.d(\M_div_src1[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[15]~q ),
	.prn(vcc));
defparam \A_mul_src1[15] .is_wysiwyg = "true";
defparam \A_mul_src1[15] .power_up = "low";

dffeas \A_dc_xfer_wr_data[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[1]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[1] .power_up = "low";

dffeas \A_dc_xfer_wr_data[4] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[4]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[4]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[4] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[4] .power_up = "low";

dffeas \A_dc_xfer_wr_data[20] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[20]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[20]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[20] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[20] .power_up = "low";

dffeas \A_dc_xfer_wr_data[12] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[12]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[12]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[12] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[12] .power_up = "low";

dffeas \A_dc_xfer_wr_data[28] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[28]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[28]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[28] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[28] .power_up = "low";

dffeas \A_mul_src2[16] (
	.clk(clk_clk),
	.d(\M_div_src2[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[16]~q ),
	.prn(vcc));
defparam \A_mul_src2[16] .is_wysiwyg = "true";
defparam \A_mul_src2[16] .power_up = "low";

dffeas \A_mul_src2[17] (
	.clk(clk_clk),
	.d(\M_div_src2[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[17]~q ),
	.prn(vcc));
defparam \A_mul_src2[17] .is_wysiwyg = "true";
defparam \A_mul_src2[17] .power_up = "low";

dffeas \A_mul_src2[18] (
	.clk(clk_clk),
	.d(\M_div_src2[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[18]~q ),
	.prn(vcc));
defparam \A_mul_src2[18] .is_wysiwyg = "true";
defparam \A_mul_src2[18] .power_up = "low";

dffeas \A_mul_src2[19] (
	.clk(clk_clk),
	.d(\M_div_src2[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[19]~q ),
	.prn(vcc));
defparam \A_mul_src2[19] .is_wysiwyg = "true";
defparam \A_mul_src2[19] .power_up = "low";

dffeas \A_mul_src2[20] (
	.clk(clk_clk),
	.d(\M_div_src2[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[20]~q ),
	.prn(vcc));
defparam \A_mul_src2[20] .is_wysiwyg = "true";
defparam \A_mul_src2[20] .power_up = "low";

dffeas \A_mul_src2[21] (
	.clk(clk_clk),
	.d(\M_div_src2[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[21]~q ),
	.prn(vcc));
defparam \A_mul_src2[21] .is_wysiwyg = "true";
defparam \A_mul_src2[21] .power_up = "low";

dffeas \A_mul_src2[22] (
	.clk(clk_clk),
	.d(\M_div_src2[22]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[22]~q ),
	.prn(vcc));
defparam \A_mul_src2[22] .is_wysiwyg = "true";
defparam \A_mul_src2[22] .power_up = "low";

dffeas \A_mul_src2[23] (
	.clk(clk_clk),
	.d(\M_div_src2[23]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[23]~q ),
	.prn(vcc));
defparam \A_mul_src2[23] .is_wysiwyg = "true";
defparam \A_mul_src2[23] .power_up = "low";

dffeas \A_mul_src2[24] (
	.clk(clk_clk),
	.d(\M_div_src2[24]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[24]~q ),
	.prn(vcc));
defparam \A_mul_src2[24] .is_wysiwyg = "true";
defparam \A_mul_src2[24] .power_up = "low";

dffeas \A_mul_src2[25] (
	.clk(clk_clk),
	.d(\M_div_src2[25]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[25]~q ),
	.prn(vcc));
defparam \A_mul_src2[25] .is_wysiwyg = "true";
defparam \A_mul_src2[25] .power_up = "low";

dffeas \A_mul_src2[26] (
	.clk(clk_clk),
	.d(\M_div_src2[26]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[26]~q ),
	.prn(vcc));
defparam \A_mul_src2[26] .is_wysiwyg = "true";
defparam \A_mul_src2[26] .power_up = "low";

dffeas \A_mul_src2[27] (
	.clk(clk_clk),
	.d(\M_div_src2[27]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[27]~q ),
	.prn(vcc));
defparam \A_mul_src2[27] .is_wysiwyg = "true";
defparam \A_mul_src2[27] .power_up = "low";

dffeas \A_mul_src2[28] (
	.clk(clk_clk),
	.d(\M_div_src2[28]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[28]~q ),
	.prn(vcc));
defparam \A_mul_src2[28] .is_wysiwyg = "true";
defparam \A_mul_src2[28] .power_up = "low";

dffeas \A_mul_src2[29] (
	.clk(clk_clk),
	.d(\M_div_src2[29]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[29]~q ),
	.prn(vcc));
defparam \A_mul_src2[29] .is_wysiwyg = "true";
defparam \A_mul_src2[29] .power_up = "low";

dffeas \A_mul_src2[30] (
	.clk(clk_clk),
	.d(\M_div_src2[30]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[30]~q ),
	.prn(vcc));
defparam \A_mul_src2[30] .is_wysiwyg = "true";
defparam \A_mul_src2[30] .power_up = "low";

dffeas \A_mul_src2[31] (
	.clk(clk_clk),
	.d(\M_div_src2[31]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[31]~q ),
	.prn(vcc));
defparam \A_mul_src2[31] .is_wysiwyg = "true";
defparam \A_mul_src2[31] .power_up = "low";

dffeas \A_dc_xfer_wr_data[16] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[16]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[16]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[16] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[16] .power_up = "low";

dffeas \A_dc_xfer_wr_data[8] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[8]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[8]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[8] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[8] .power_up = "low";

dffeas \A_dc_xfer_wr_data[24] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[24]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[24]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[24] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[24] .power_up = "low";

dffeas \A_dc_xfer_wr_data[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[2]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[2] .power_up = "low";

dffeas \A_dc_xfer_wr_data[18] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[18]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[18]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[18] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[18] .power_up = "low";

dffeas \A_dc_xfer_wr_data[10] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[10]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[10]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[10] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[10] .power_up = "low";

dffeas \A_dc_xfer_wr_data[26] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[26]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[26]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[26] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[26] .power_up = "low";

dffeas \A_dc_xfer_wr_data[5] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[5]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[5]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[5] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[5] .power_up = "low";

dffeas \A_dc_xfer_wr_data[21] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[21]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[21]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[21] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[21] .power_up = "low";

dffeas \A_dc_xfer_wr_data[13] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[13]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[13]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[13] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[13] .power_up = "low";

dffeas \A_dc_xfer_wr_data[29] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[29]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[29]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[29] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[29] .power_up = "low";

dffeas \A_dc_xfer_wr_data[23] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[23]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[23]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[23] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[23] .power_up = "low";

dffeas \A_dc_xfer_wr_data[15] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[15]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[15]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[15] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[15] .power_up = "low";

dffeas \A_dc_xfer_wr_data[31] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[31]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[31]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[31] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[31] .power_up = "low";

dffeas \A_dc_xfer_wr_data[11] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[11]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[11]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[11] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[11] .power_up = "low";

dffeas \A_dc_xfer_wr_data[27] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[27]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[27]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[27] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[27] .power_up = "low";

dffeas \A_dc_xfer_wr_data[9] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[9]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[9]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[9] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[9] .power_up = "low";

dffeas \A_dc_xfer_wr_data[25] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[25]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[25]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[25] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[25] .power_up = "low";

dffeas \A_dc_xfer_wr_data[6] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[6]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[6]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[6] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[6] .power_up = "low";

dffeas \A_dc_xfer_wr_data[22] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[22]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[22]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[22] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[22] .power_up = "low";

dffeas \A_dc_xfer_wr_data[14] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[14]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[14]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[14] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[14] .power_up = "low";

dffeas \A_dc_xfer_wr_data[30] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[30]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[30]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[30] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[30] .power_up = "low";

dffeas \A_mul_src1[16] (
	.clk(clk_clk),
	.d(\M_div_src1[16]~q ),
	.asdata(\A_mul_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[16]~q ),
	.prn(vcc));
defparam \A_mul_src1[16] .is_wysiwyg = "true";
defparam \A_mul_src1[16] .power_up = "low";

dffeas \A_mul_src1[17] (
	.clk(clk_clk),
	.d(\M_div_src1[17]~q ),
	.asdata(\A_mul_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[17]~q ),
	.prn(vcc));
defparam \A_mul_src1[17] .is_wysiwyg = "true";
defparam \A_mul_src1[17] .power_up = "low";

dffeas \A_mul_src1[18] (
	.clk(clk_clk),
	.d(\M_div_src1[18]~q ),
	.asdata(\A_mul_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[18]~q ),
	.prn(vcc));
defparam \A_mul_src1[18] .is_wysiwyg = "true";
defparam \A_mul_src1[18] .power_up = "low";

dffeas \A_mul_src1[19] (
	.clk(clk_clk),
	.d(\M_div_src1[19]~q ),
	.asdata(\A_mul_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[19]~q ),
	.prn(vcc));
defparam \A_mul_src1[19] .is_wysiwyg = "true";
defparam \A_mul_src1[19] .power_up = "low";

dffeas \A_mul_src1[20] (
	.clk(clk_clk),
	.d(\M_div_src1[20]~q ),
	.asdata(\A_mul_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[20]~q ),
	.prn(vcc));
defparam \A_mul_src1[20] .is_wysiwyg = "true";
defparam \A_mul_src1[20] .power_up = "low";

dffeas \A_mul_src1[21] (
	.clk(clk_clk),
	.d(\M_div_src1[21]~q ),
	.asdata(\A_mul_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[21]~q ),
	.prn(vcc));
defparam \A_mul_src1[21] .is_wysiwyg = "true";
defparam \A_mul_src1[21] .power_up = "low";

dffeas \A_mul_src1[22] (
	.clk(clk_clk),
	.d(\M_div_src1[22]~q ),
	.asdata(\A_mul_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[22]~q ),
	.prn(vcc));
defparam \A_mul_src1[22] .is_wysiwyg = "true";
defparam \A_mul_src1[22] .power_up = "low";

dffeas \A_mul_src1[23] (
	.clk(clk_clk),
	.d(\M_div_src1[23]~q ),
	.asdata(\A_mul_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[23]~q ),
	.prn(vcc));
defparam \A_mul_src1[23] .is_wysiwyg = "true";
defparam \A_mul_src1[23] .power_up = "low";

dffeas \A_mul_src1[24] (
	.clk(clk_clk),
	.d(\M_div_src1[24]~q ),
	.asdata(\A_mul_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[24]~q ),
	.prn(vcc));
defparam \A_mul_src1[24] .is_wysiwyg = "true";
defparam \A_mul_src1[24] .power_up = "low";

dffeas \A_mul_src1[25] (
	.clk(clk_clk),
	.d(\M_div_src1[25]~q ),
	.asdata(\A_mul_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[25]~q ),
	.prn(vcc));
defparam \A_mul_src1[25] .is_wysiwyg = "true";
defparam \A_mul_src1[25] .power_up = "low";

dffeas \A_mul_src1[26] (
	.clk(clk_clk),
	.d(\M_div_src1[26]~q ),
	.asdata(\A_mul_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[26]~q ),
	.prn(vcc));
defparam \A_mul_src1[26] .is_wysiwyg = "true";
defparam \A_mul_src1[26] .power_up = "low";

dffeas \A_mul_src1[27] (
	.clk(clk_clk),
	.d(\M_div_src1[27]~q ),
	.asdata(\A_mul_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[27]~q ),
	.prn(vcc));
defparam \A_mul_src1[27] .is_wysiwyg = "true";
defparam \A_mul_src1[27] .power_up = "low";

dffeas \A_mul_src1[28] (
	.clk(clk_clk),
	.d(\M_div_src1[28]~q ),
	.asdata(\A_mul_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[28]~q ),
	.prn(vcc));
defparam \A_mul_src1[28] .is_wysiwyg = "true";
defparam \A_mul_src1[28] .power_up = "low";

dffeas \A_mul_src1[29] (
	.clk(clk_clk),
	.d(\M_div_src1[29]~q ),
	.asdata(\A_mul_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[29]~q ),
	.prn(vcc));
defparam \A_mul_src1[29] .is_wysiwyg = "true";
defparam \A_mul_src1[29] .power_up = "low";

dffeas \A_mul_src1[30] (
	.clk(clk_clk),
	.d(\M_div_src1[30]~q ),
	.asdata(\A_mul_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[30]~q ),
	.prn(vcc));
defparam \A_mul_src1[30] .is_wysiwyg = "true";
defparam \A_mul_src1[30] .power_up = "low";

dffeas \A_mul_src1[31] (
	.clk(clk_clk),
	.d(\M_div_src1[31]~q ),
	.asdata(\A_mul_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[31]~q ),
	.prn(vcc));
defparam \A_mul_src1[31] .is_wysiwyg = "true";
defparam \A_mul_src1[31] .power_up = "low";

dffeas \A_dc_xfer_wr_data[19] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[19]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[19]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[19] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[19] .power_up = "low";

dffeas \A_dc_xfer_wr_data[17] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[17]~q ),
	.asdata(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[17]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[17] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[17] .power_up = "low";

dffeas A_dc_xfer_wr_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_data_active~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_active~q ),
	.prn(vcc));
defparam A_dc_xfer_wr_active.is_wysiwyg = "true";
defparam A_dc_xfer_wr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_wb_rd_en~0 (
	.dataa(!\A_dc_wb_rd_data_starting~q ),
	.datab(!\A_dc_wb_rd_addr_starting~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_en~0 .extended_lut = "off";
defparam \A_dc_wb_rd_en~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_wb_rd_en~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_wb_rd_en(
	.dataa(!rst1),
	.datab(!d_write1),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(!\A_dc_wb_wr_starting~combout ),
	.dataf(!\A_dc_wb_rd_en~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_rd_en.extended_lut = "off";
defparam A_dc_wb_rd_en.lut_mask = 64'hFFFFFFFFFFF7FFFF;
defparam A_dc_wb_rd_en.shared_arith = "off";

dffeas \A_dc_xfer_wr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[0] .power_up = "low";

dffeas \A_dc_xfer_wr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[1] .power_up = "low";

dffeas \A_dc_xfer_wr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[2] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[0] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[1] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[2] .power_up = "low";

dffeas A_dc_fill_starting_d1(
	.clk(clk_clk),
	.d(\A_dc_fill_starting~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_starting_d1~q ),
	.prn(vcc));
defparam A_dc_fill_starting_d1.is_wysiwyg = "true";
defparam A_dc_fill_starting_d1.power_up = "low";

dffeas A_en_d1(
	.clk(clk_clk),
	.d(\A_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_en_d1~q ),
	.prn(vcc));
defparam A_en_d1.is_wysiwyg = "true";
defparam A_en_d1.power_up = "low";

dffeas A_ctrl_dc_index_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_index_inv~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_index_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_index_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_index_inv.power_up = "low";

dffeas A_ctrl_dc_addr_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_addr_inv~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_addr_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_addr_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_addr_inv.power_up = "low";

cyclonev_lcell_comb \A_dc_tag_dcache_management_wr_en~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_dc_hit~q ),
	.datac(!\A_en_d1~q ),
	.datad(!\A_ctrl_dc_index_inv~q ),
	.datae(!\A_ctrl_dc_addr_inv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_tag_dcache_management_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_tag_dcache_management_wr_en~0 .extended_lut = "off";
defparam \A_dc_tag_dcache_management_wr_en~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \A_dc_tag_dcache_management_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[5]~0 (
	.dataa(!\A_dc_fill_starting_d1~q ),
	.datab(!\A_dc_tag_dcache_management_wr_en~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[5]~0 .extended_lut = "off";
defparam \dc_tag_wr_port_data[5]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \dc_tag_wr_port_data[5]~0 .shared_arith = "off";

cyclonev_lcell_comb dc_tag_wr_port_en(
	.dataa(!\A_div_done~q ),
	.datab(!\A_mem_stall~q ),
	.datac(!\A_mul_stall~q ),
	.datad(!\A_div_stall~0_combout ),
	.datae(!\M_dc_valid_st_cache_hit~0_combout ),
	.dataf(!\dc_tag_wr_port_data[5]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam dc_tag_wr_port_en.extended_lut = "off";
defparam dc_tag_wr_port_en.lut_mask = 64'hFFFFFFFFFFFDFFFF;
defparam dc_tag_wr_port_en.shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[4]~1 (
	.dataa(!\A_mem_baddr[15]~q ),
	.datab(!\M_alu_result[15]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[4]~1 .extended_lut = "off";
defparam \dc_tag_wr_port_data[4]~1 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[0]~0 (
	.dataa(!\A_mem_baddr[5]~q ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[0]~0 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[0]~0 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[1]~1 (
	.dataa(!\A_mem_baddr[6]~q ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[1]~1 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[1]~1 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[2]~2 (
	.dataa(!\A_mem_baddr[7]~q ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[2]~2 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[2]~2 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[3]~3 (
	.dataa(!\A_mem_baddr[8]~q ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[3]~3 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[3]~3 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[4]~4 (
	.dataa(!\A_mem_baddr[9]~q ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[4]~4 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[4]~4 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[5]~5 (
	.dataa(!\A_mem_baddr[10]~q ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[5]~5 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[5]~5 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\Add24~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[0]~0 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\Add24~21_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[1]~1 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\Add24~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[2]~2 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\Add24~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[3]~3 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\Add24~5_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[4]~4 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[5]~5 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\Add24~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[5]~5 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[5]~2 (
	.dataa(!\A_mem_baddr[16]~q ),
	.datab(!\M_alu_result[16]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[5]~2 .extended_lut = "off";
defparam \dc_tag_wr_port_data[5]~2 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[6]~3 (
	.dataa(!\A_dc_fill_starting_d1~q ),
	.datab(!\A_dc_tag_dcache_management_wr_en~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[6]~3 .extended_lut = "off";
defparam \dc_tag_wr_port_data[6]~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \dc_tag_wr_port_data[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[0]~4 (
	.dataa(!\A_mem_baddr[11]~q ),
	.datab(!\M_alu_result[11]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[0]~4 .extended_lut = "off";
defparam \dc_tag_wr_port_data[0]~4 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[1]~5 (
	.dataa(!\A_mem_baddr[12]~q ),
	.datab(!\M_alu_result[12]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[1]~5 .extended_lut = "off";
defparam \dc_tag_wr_port_data[1]~5 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[2]~6 (
	.dataa(!\A_mem_baddr[13]~q ),
	.datab(!\M_alu_result[13]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[2]~6 .extended_lut = "off";
defparam \dc_tag_wr_port_data[2]~6 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[3]~7 (
	.dataa(!\A_mem_baddr[14]~q ),
	.datab(!\M_alu_result[14]~q ),
	.datac(!\dc_tag_wr_port_data[5]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[3]~7 .extended_lut = "off";
defparam \dc_tag_wr_port_data[3]~7 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[3]~7 .shared_arith = "off";

dffeas A_dc_xfer_rd_data_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_active~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_active~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_active.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_active.power_up = "low";

dffeas \A_dc_rd_data[0] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[0] .is_wysiwyg = "true";
defparam \A_dc_rd_data[0] .power_up = "low";

dffeas A_dc_xfer_rd_data_offset_match(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_match~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_offset_match~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_offset_match.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_offset_match.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[0]~0 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_starting~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[1]~1 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_offset[1]~q ),
	.datac(!\A_dc_xfer_wr_starting~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .lut_mask = 64'hF6F6F6F6F6F6F6F6;
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[2]~2 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_offset[1]~q ),
	.datac(!\A_dc_xfer_wr_offset[2]~q ),
	.datad(!\A_dc_xfer_wr_starting~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .lut_mask = 64'hFF96FF96FF96FF96;
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[0]~0 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[1]~1 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(!\A_dc_wb_rd_addr_offset[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[2]~2 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(!\A_dc_wb_rd_addr_offset[1]~q ),
	.datad(!\A_dc_wb_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .shared_arith = "off";

dffeas M_ctrl_dc_index_inv(
	.clk(clk_clk),
	.d(\E_ctrl_dc_index_inv~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_index_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_index_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_index_inv.power_up = "low";

dffeas M_ctrl_dc_addr_inv(
	.clk(clk_clk),
	.d(\E_ctrl_dc_addr_inv~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_addr_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_addr_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_addr_inv.power_up = "low";

dffeas A_valid_st_writes_mem(
	.clk(clk_clk),
	.d(\M_valid_st_writes_mem~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_valid_st_writes_mem~q ),
	.prn(vcc));
defparam A_valid_st_writes_mem.is_wysiwyg = "true";
defparam A_valid_st_writes_mem.power_up = "low";

cyclonev_lcell_comb \dc_tag_wr_port_data[7]~8 (
	.dataa(!\A_dc_fill_starting_d1~q ),
	.datab(!\A_dc_tag_dcache_management_wr_en~0_combout ),
	.datac(!\A_valid_st_writes_mem~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[7]~8 .extended_lut = "off";
defparam \dc_tag_wr_port_data[7]~8 .lut_mask = 64'h8D8D8D8D8D8D8D8D;
defparam \dc_tag_wr_port_data[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[22]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_b_rd_port_addr[0]~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[23]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_b_rd_port_addr[1]~1 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[24]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_b_rd_port_addr[2]~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[25]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_b_rd_port_addr[3]~3 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[26]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_b_rd_port_addr[4]~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[27]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_a_rd_port_addr[0]~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[28]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_a_rd_port_addr[1]~1 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[29]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_a_rd_port_addr[2]~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[30]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_a_rd_port_addr[3]~3 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[31]~q ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_a_rd_port_addr[4]~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb A_dc_valid_st_bypass_hit_wr_en(
	.dataa(!\A_dc_valid_st_bypass_hit~q ),
	.datab(!\A_en_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_valid_st_bypass_hit_wr_en.extended_lut = "off";
defparam A_dc_valid_st_bypass_hit_wr_en.lut_mask = 64'h7777777777777777;
defparam A_dc_valid_st_bypass_hit_wr_en.shared_arith = "off";

cyclonev_lcell_comb dc_data_wr_port_en(
	.dataa(!\A_stall~combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\d_readdatavalid_d1~q ),
	.datad(!\M_dc_valid_st_cache_hit~0_combout ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam dc_data_wr_port_en.extended_lut = "off";
defparam dc_data_wr_port_en.lut_mask = 64'h47FFFFFF47FFFFFF;
defparam dc_data_wr_port_en.shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[0]~0 (
	.dataa(!\M_st_data[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\M_mem_byte_en[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[0]~0 .extended_lut = "off";
defparam \M_dc_st_data[0]~0 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[0]~0 .shared_arith = "off";

dffeas \A_dc_st_data[0] (
	.clk(clk_clk),
	.d(\M_dc_st_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[0]~q ),
	.prn(vcc));
defparam \A_dc_st_data[0] .is_wysiwyg = "true";
defparam \A_dc_st_data[0] .power_up = "low";

dffeas A_ctrl_st(
	.clk(clk_clk),
	.d(\M_ctrl_st~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_st~q ),
	.prn(vcc));
defparam A_ctrl_st.is_wysiwyg = "true";
defparam A_ctrl_st.power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[6]~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal263~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_mem_byte_en[0]~q ),
	.dataf(!\A_ctrl_st~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[6]~0 .extended_lut = "off";
defparam \dc_data_wr_port_data[6]~0 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[0]~1 (
	.dataa(!\M_dc_st_data[0]~0_combout ),
	.datab(!\A_dc_st_data[0]~q ),
	.datac(!\d_readdata_d1[0]~q ),
	.datad(!\A_st_data[0]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[0]~1 .extended_lut = "off";
defparam \dc_data_wr_port_data[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[0]~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[2]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\A_dc_fill_dp_offset[0]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[0]~0 .extended_lut = "off";
defparam \dc_data_wr_port_addr[0]~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_wr_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[1]~1 (
	.dataa(!\A_mem_baddr[3]~q ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\A_dc_fill_active~q ),
	.datad(!\A_dc_fill_dp_offset[1]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[1]~1 .extended_lut = "off";
defparam \dc_data_wr_port_addr[1]~1 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \dc_data_wr_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[2]~2 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[4]~q ),
	.datac(!\M_alu_result[4]~q ),
	.datad(!\A_dc_fill_dp_offset[2]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[2]~2 .extended_lut = "off";
defparam \dc_data_wr_port_addr[2]~2 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_wr_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[3]~3 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[5]~q ),
	.datac(!\M_alu_result[5]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[3]~3 .extended_lut = "off";
defparam \dc_data_wr_port_addr[3]~3 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[4]~4 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[6]~q ),
	.datac(!\M_alu_result[6]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[4]~4 .extended_lut = "off";
defparam \dc_data_wr_port_addr[4]~4 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[5]~5 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[7]~q ),
	.datac(!\M_alu_result[7]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[5]~5 .extended_lut = "off";
defparam \dc_data_wr_port_addr[5]~5 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[6]~6 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[8]~q ),
	.datac(!\M_alu_result[8]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[6]~6 .extended_lut = "off";
defparam \dc_data_wr_port_addr[6]~6 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[7]~7 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[9]~q ),
	.datac(!\M_alu_result[9]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[7]~7 .extended_lut = "off";
defparam \dc_data_wr_port_addr[7]~7 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[8]~8 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[10]~q ),
	.datac(!\M_alu_result[10]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[8]~8 .extended_lut = "off";
defparam \dc_data_wr_port_addr[8]~8 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[2]~q ),
	.datac(!\Add24~25_sumout ),
	.datad(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[0]~0 .extended_lut = "off";
defparam \dc_data_rd_port_addr[0]~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\Add24~29_sumout ),
	.datad(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[1]~1 .extended_lut = "off";
defparam \dc_data_rd_port_addr[1]~1 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[4]~q ),
	.datac(!\Add24~33_sumout ),
	.datad(!\A_dc_xfer_rd_addr_active~q ),
	.datae(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[2]~2 .extended_lut = "off";
defparam \dc_data_rd_port_addr[2]~2 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \dc_data_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[5]~q ),
	.datac(!\M_alu_result[5]~q ),
	.datad(!\Add24~17_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[3]~3 .extended_lut = "off";
defparam \dc_data_rd_port_addr[3]~3 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[6]~q ),
	.datac(!\M_alu_result[6]~q ),
	.datad(!\Add24~21_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[4]~4 .extended_lut = "off";
defparam \dc_data_rd_port_addr[4]~4 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[5]~5 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[7]~q ),
	.datac(!\M_alu_result[7]~q ),
	.datad(!\Add24~9_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[5]~5 .extended_lut = "off";
defparam \dc_data_rd_port_addr[5]~5 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[6]~6 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[8]~q ),
	.datac(!\M_alu_result[8]~q ),
	.datad(!\Add24~1_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[6]~6 .extended_lut = "off";
defparam \dc_data_rd_port_addr[6]~6 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[7]~7 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[9]~q ),
	.datac(!\M_alu_result[9]~q ),
	.datad(!\Add24~5_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[7]~7 .extended_lut = "off";
defparam \dc_data_rd_port_addr[7]~7 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[8]~8 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[10]~q ),
	.datac(!\M_alu_result[10]~q ),
	.datad(!\Add24~13_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[8]~8 .extended_lut = "off";
defparam \dc_data_rd_port_addr[8]~8 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_match~0 (
	.dataa(!\A_mem_baddr[2]~q ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(!\A_valid_st_writes_mem~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_match~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_match~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_match~0 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \A_dc_xfer_rd_addr_offset_match~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_xfer_rd_addr_offset_match(
	.dataa(!\A_mem_baddr[3]~q ),
	.datab(!\A_mem_baddr[4]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(!\A_dc_xfer_rd_addr_offset_match~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_match~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_xfer_rd_addr_offset_match.extended_lut = "off";
defparam A_dc_xfer_rd_addr_offset_match.lut_mask = 64'h6996FFFF6996FFFF;
defparam A_dc_xfer_rd_addr_offset_match.shared_arith = "off";

dffeas ic_tag_clr_valid_bits(
	.clk(clk_clk),
	.d(\ic_tag_clr_valid_bits~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_clr_valid_bits~q ),
	.prn(vcc));
defparam ic_tag_clr_valid_bits.is_wysiwyg = "true";
defparam ic_tag_clr_valid_bits.power_up = "low";

cyclonev_lcell_comb ic_tag_wren(
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_tag_clr_valid_bits~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_wren.extended_lut = "off";
defparam ic_tag_wren.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ic_tag_wren.shared_arith = "off";

dffeas \ic_tag_wraddress[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[0]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[0] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[0] .power_up = "low";

dffeas \ic_tag_wraddress[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[1]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[1]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[1] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[1] .power_up = "low";

dffeas \ic_tag_wraddress[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[2]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[2] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[2] .power_up = "low";

dffeas \ic_tag_wraddress[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[3]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[3]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[3] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[3] .power_up = "low";

dffeas \ic_tag_wraddress[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[4]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[4]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[4] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[4] .power_up = "low";

dffeas \ic_tag_wraddress[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[5]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[5]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[5] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[5] .power_up = "low";

dffeas \ic_tag_wraddress[6] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[6]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[6]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[6] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[6] .power_up = "low";

dffeas \i_readdata_d1[5] (
	.clk(clk_clk),
	.d(i_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[5]~q ),
	.prn(vcc));
defparam \i_readdata_d1[5] .is_wysiwyg = "true";
defparam \i_readdata_d1[5] .power_up = "low";

dffeas \i_readdata_d1[3] (
	.clk(clk_clk),
	.d(i_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[3]~q ),
	.prn(vcc));
defparam \i_readdata_d1[3] .is_wysiwyg = "true";
defparam \i_readdata_d1[3] .power_up = "low";

dffeas \i_readdata_d1[1] (
	.clk(clk_clk),
	.d(i_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[1]~q ),
	.prn(vcc));
defparam \i_readdata_d1[1] .is_wysiwyg = "true";
defparam \i_readdata_d1[1] .power_up = "low";

dffeas \i_readdata_d1[4] (
	.clk(clk_clk),
	.d(i_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[4]~q ),
	.prn(vcc));
defparam \i_readdata_d1[4] .is_wysiwyg = "true";
defparam \i_readdata_d1[4] .power_up = "low";

dffeas \i_readdata_d1[2] (
	.clk(clk_clk),
	.d(i_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[2]~q ),
	.prn(vcc));
defparam \i_readdata_d1[2] .is_wysiwyg = "true";
defparam \i_readdata_d1[2] .power_up = "low";

dffeas \i_readdata_d1[28] (
	.clk(clk_clk),
	.d(i_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[28]~q ),
	.prn(vcc));
defparam \i_readdata_d1[28] .is_wysiwyg = "true";
defparam \i_readdata_d1[28] .power_up = "low";

dffeas \i_readdata_d1[30] (
	.clk(clk_clk),
	.d(i_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[30]~q ),
	.prn(vcc));
defparam \i_readdata_d1[30] .is_wysiwyg = "true";
defparam \i_readdata_d1[30] .power_up = "low";

dffeas \i_readdata_d1[31] (
	.clk(clk_clk),
	.d(i_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[31]~q ),
	.prn(vcc));
defparam \i_readdata_d1[31] .is_wysiwyg = "true";
defparam \i_readdata_d1[31] .power_up = "low";

dffeas \i_readdata_d1[27] (
	.clk(clk_clk),
	.d(i_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[27]~q ),
	.prn(vcc));
defparam \i_readdata_d1[27] .is_wysiwyg = "true";
defparam \i_readdata_d1[27] .power_up = "low";

dffeas \i_readdata_d1[29] (
	.clk(clk_clk),
	.d(i_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[29]~q ),
	.prn(vcc));
defparam \i_readdata_d1[29] .is_wysiwyg = "true";
defparam \i_readdata_d1[29] .power_up = "low";

dffeas \i_readdata_d1[0] (
	.clk(clk_clk),
	.d(i_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[0]~q ),
	.prn(vcc));
defparam \i_readdata_d1[0] .is_wysiwyg = "true";
defparam \i_readdata_d1[0] .power_up = "low";

dffeas \i_readdata_d1[23] (
	.clk(clk_clk),
	.d(i_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[23]~q ),
	.prn(vcc));
defparam \i_readdata_d1[23] .is_wysiwyg = "true";
defparam \i_readdata_d1[23] .power_up = "low";

dffeas \i_readdata_d1[25] (
	.clk(clk_clk),
	.d(i_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[25]~q ),
	.prn(vcc));
defparam \i_readdata_d1[25] .is_wysiwyg = "true";
defparam \i_readdata_d1[25] .power_up = "low";

dffeas \i_readdata_d1[26] (
	.clk(clk_clk),
	.d(i_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[26]~q ),
	.prn(vcc));
defparam \i_readdata_d1[26] .is_wysiwyg = "true";
defparam \i_readdata_d1[26] .power_up = "low";

dffeas \i_readdata_d1[22] (
	.clk(clk_clk),
	.d(i_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[22]~q ),
	.prn(vcc));
defparam \i_readdata_d1[22] .is_wysiwyg = "true";
defparam \i_readdata_d1[22] .power_up = "low";

dffeas \i_readdata_d1[24] (
	.clk(clk_clk),
	.d(i_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[24]~q ),
	.prn(vcc));
defparam \i_readdata_d1[24] .is_wysiwyg = "true";
defparam \i_readdata_d1[24] .power_up = "low";

dffeas \i_readdata_d1[16] (
	.clk(clk_clk),
	.d(i_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[16]~q ),
	.prn(vcc));
defparam \i_readdata_d1[16] .is_wysiwyg = "true";
defparam \i_readdata_d1[16] .power_up = "low";

dffeas \i_readdata_d1[15] (
	.clk(clk_clk),
	.d(i_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[15]~q ),
	.prn(vcc));
defparam \i_readdata_d1[15] .is_wysiwyg = "true";
defparam \i_readdata_d1[15] .power_up = "low";

dffeas \i_readdata_d1[13] (
	.clk(clk_clk),
	.d(i_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[13]~q ),
	.prn(vcc));
defparam \i_readdata_d1[13] .is_wysiwyg = "true";
defparam \i_readdata_d1[13] .power_up = "low";

dffeas \i_readdata_d1[14] (
	.clk(clk_clk),
	.d(i_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[14]~q ),
	.prn(vcc));
defparam \i_readdata_d1[14] .is_wysiwyg = "true";
defparam \i_readdata_d1[14] .power_up = "low";

dffeas \i_readdata_d1[12] (
	.clk(clk_clk),
	.d(i_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[12]~q ),
	.prn(vcc));
defparam \i_readdata_d1[12] .is_wysiwyg = "true";
defparam \i_readdata_d1[12] .power_up = "low";

dffeas \i_readdata_d1[11] (
	.clk(clk_clk),
	.d(i_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[11]~q ),
	.prn(vcc));
defparam \i_readdata_d1[11] .is_wysiwyg = "true";
defparam \i_readdata_d1[11] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_dc_index_inv~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_dc_index_inv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_dc_index_inv~0 .extended_lut = "off";
defparam \E_ctrl_dc_index_inv~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_ctrl_dc_index_inv~0 .shared_arith = "off";

dffeas M_ctrl_st(
	.clk(clk_clk),
	.d(\M_ctrl_st_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st~q ),
	.prn(vcc));
defparam M_ctrl_st.is_wysiwyg = "true";
defparam M_ctrl_st.power_up = "low";

cyclonev_lcell_comb M_valid_st_writes_mem(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_valid_st_writes_mem~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_valid_st_writes_mem.extended_lut = "off";
defparam M_valid_st_writes_mem.lut_mask = 64'h7777777777777777;
defparam M_valid_st_writes_mem.shared_arith = "off";

dffeas \i_readdata_d1[10] (
	.clk(clk_clk),
	.d(i_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[10]~q ),
	.prn(vcc));
defparam \i_readdata_d1[10] .is_wysiwyg = "true";
defparam \i_readdata_d1[10] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[4]~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\M_mem_byte_en[0]~q ),
	.datac(!\M_st_data[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[4]~1 .extended_lut = "off";
defparam \M_dc_st_data[4]~1 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[4]~1 .shared_arith = "off";

dffeas \A_dc_st_data[4] (
	.clk(clk_clk),
	.d(\M_dc_st_data[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[4]~q ),
	.prn(vcc));
defparam \A_dc_st_data[4] .is_wysiwyg = "true";
defparam \A_dc_st_data[4] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[4]~2 (
	.dataa(!\M_dc_st_data[4]~1_combout ),
	.datab(!\A_dc_st_data[4]~q ),
	.datac(!\d_readdata_d1[4]~q ),
	.datad(!\A_st_data[4]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[4]~2 .extended_lut = "off";
defparam \dc_data_wr_port_data[4]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[20]~2 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[20]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[20]~2 .extended_lut = "off";
defparam \M_dc_st_data[20]~2 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[20]~2 .shared_arith = "off";

dffeas \A_dc_st_data[20] (
	.clk(clk_clk),
	.d(\M_dc_st_data[20]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[20]~q ),
	.prn(vcc));
defparam \A_dc_st_data[20] .is_wysiwyg = "true";
defparam \A_dc_st_data[20] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[18]~3 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal263~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_byte_en[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[18]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[18]~3 .extended_lut = "off";
defparam \dc_data_wr_port_data[18]~3 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[18]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[20]~4 (
	.dataa(!\M_dc_st_data[20]~2_combout ),
	.datab(!\A_dc_st_data[20]~q ),
	.datac(!\d_readdata_d1[20]~q ),
	.datad(!\A_st_data[20]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[20]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[20]~4 .extended_lut = "off";
defparam \dc_data_wr_port_data[20]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[20]~4 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[12]~3 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[12]~3 .extended_lut = "off";
defparam \M_dc_st_data[12]~3 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[12]~3 .shared_arith = "off";

dffeas \A_dc_st_data[12] (
	.clk(clk_clk),
	.d(\M_dc_st_data[12]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[12]~q ),
	.prn(vcc));
defparam \A_dc_st_data[12] .is_wysiwyg = "true";
defparam \A_dc_st_data[12] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[12]~5 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal263~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_byte_en[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[12]~5 .extended_lut = "off";
defparam \dc_data_wr_port_data[12]~5 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[12]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[12]~6 (
	.dataa(!\M_dc_st_data[12]~3_combout ),
	.datab(!\A_dc_st_data[12]~q ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\A_st_data[12]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[12]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[12]~6 .extended_lut = "off";
defparam \dc_data_wr_port_data[12]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[12]~6 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[28]~4 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[28]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[28]~4 .extended_lut = "off";
defparam \M_dc_st_data[28]~4 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[28]~4 .shared_arith = "off";

dffeas \A_dc_st_data[28] (
	.clk(clk_clk),
	.d(\M_dc_st_data[28]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[28]~q ),
	.prn(vcc));
defparam \A_dc_st_data[28] .is_wysiwyg = "true";
defparam \A_dc_st_data[28] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[31]~7 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal263~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_byte_en[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[31]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[31]~7 .extended_lut = "off";
defparam \dc_data_wr_port_data[31]~7 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[31]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[28]~8 (
	.dataa(!\M_dc_st_data[28]~4_combout ),
	.datab(!\A_dc_st_data[28]~q ),
	.datac(!\d_readdata_d1[28]~q ),
	.datad(!\A_st_data[28]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[28]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[28]~8 .extended_lut = "off";
defparam \dc_data_wr_port_data[28]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[28]~8 .shared_arith = "off";

dffeas M_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_br_cond~q ),
	.prn(vcc));
defparam M_ctrl_br_cond.is_wysiwyg = "true";
defparam M_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb M_bht_wr_en_unfiltered(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_br_cond~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_en_unfiltered~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_bht_wr_en_unfiltered.extended_lut = "off";
defparam M_bht_wr_en_unfiltered.lut_mask = 64'h7777777777777777;
defparam M_bht_wr_en_unfiltered.shared_arith = "off";

dffeas \M_bht_data[1] (
	.clk(clk_clk),
	.d(\E_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_data[1]~q ),
	.prn(vcc));
defparam \M_bht_data[1] .is_wysiwyg = "true";
defparam \M_bht_data[1] .power_up = "low";

dffeas \M_bht_data[0] (
	.clk(clk_clk),
	.d(\E_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_data[0]~q ),
	.prn(vcc));
defparam \M_bht_data[0] .is_wysiwyg = "true";
defparam \M_bht_data[0] .power_up = "low";

dffeas M_br_mispredict(
	.clk(clk_clk),
	.d(\E_br_mispredict~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_br_mispredict~q ),
	.prn(vcc));
defparam M_br_mispredict.is_wysiwyg = "true";
defparam M_br_mispredict.power_up = "low";

cyclonev_lcell_comb \M_bht_wr_data_unfiltered[1]~0 (
	.dataa(!\M_bht_data[1]~q ),
	.datab(!\M_bht_data[0]~q ),
	.datac(!\M_br_mispredict~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_bht_wr_data_unfiltered[1]~0 .extended_lut = "off";
defparam \M_bht_wr_data_unfiltered[1]~0 .lut_mask = 64'h9696969696969696;
defparam \M_bht_wr_data_unfiltered[1]~0 .shared_arith = "off";

dffeas \M_bht_ptr_unfiltered[0] (
	.clk(clk_clk),
	.d(\E_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[0]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[0] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[0] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[1] (
	.clk(clk_clk),
	.d(\E_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[1]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[1] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[1] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[2] (
	.clk(clk_clk),
	.d(\E_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[2]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[2] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[2] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[3] (
	.clk(clk_clk),
	.d(\E_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[3]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[3] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[3] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[4] (
	.clk(clk_clk),
	.d(\E_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[4]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[4] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[4] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[5] (
	.clk(clk_clk),
	.d(\E_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[5]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[5] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[5] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[6] (
	.clk(clk_clk),
	.d(\E_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[6]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[6] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[6] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[7] (
	.clk(clk_clk),
	.d(\E_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[7]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[7] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[7] .power_up = "low";

dffeas \M_br_cond_taken_history[0] (
	.clk(clk_clk),
	.d(\E_br_result~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[0]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[0] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[0] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[0] (
	.dataa(!\E_src1[2]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\M_br_cond_taken_history[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[0] .extended_lut = "off";
defparam \F_bht_ptr_nxt[0] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[0] .shared_arith = "off";

dffeas \M_br_cond_taken_history[1] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[1]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[1] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[1] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[1] (
	.dataa(!\E_src1[3]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[1]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.dataf(!\M_br_cond_taken_history[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[1] .extended_lut = "off";
defparam \F_bht_ptr_nxt[1] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[1] .shared_arith = "off";

dffeas \M_br_cond_taken_history[2] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[2]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[2] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[2] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[2] (
	.dataa(!\E_src1[4]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[2]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~4_combout ),
	.dataf(!\M_br_cond_taken_history[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[2] .extended_lut = "off";
defparam \F_bht_ptr_nxt[2] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[2] .shared_arith = "off";

dffeas \M_br_cond_taken_history[3] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[3]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[3] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[3] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[3] (
	.dataa(!\E_src1[5]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[3]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[0]~12_combout ),
	.dataf(!\M_br_cond_taken_history[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[3] .extended_lut = "off";
defparam \F_bht_ptr_nxt[3] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[3] .shared_arith = "off";

dffeas \M_br_cond_taken_history[4] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[4]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[4] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[4] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[4] (
	.dataa(!\E_src1[6]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[4]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[1]~8_combout ),
	.dataf(!\M_br_cond_taken_history[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[4] .extended_lut = "off";
defparam \F_bht_ptr_nxt[4] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[4] .shared_arith = "off";

dffeas \M_br_cond_taken_history[5] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[5]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[5] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[5] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[5] (
	.dataa(!\E_src1[7]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[5]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[2]~10_combout ),
	.dataf(!\M_br_cond_taken_history[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[5] .extended_lut = "off";
defparam \F_bht_ptr_nxt[5] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[5] .shared_arith = "off";

dffeas \M_br_cond_taken_history[6] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[6]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[6] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[6] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[6] (
	.dataa(!\E_src1[8]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.dataf(!\M_br_cond_taken_history[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[6] .extended_lut = "off";
defparam \F_bht_ptr_nxt[6] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[6] .shared_arith = "off";

dffeas \M_br_cond_taken_history[7] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[7]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[7] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[7] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[7] (
	.dataa(!\E_src1[9]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[4]~2_combout ),
	.dataf(!\M_br_cond_taken_history[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[7] .extended_lut = "off";
defparam \F_bht_ptr_nxt[7] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[7] .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[16]~5 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[16]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[16]~5 .extended_lut = "off";
defparam \M_dc_st_data[16]~5 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[16]~5 .shared_arith = "off";

dffeas \A_dc_st_data[16] (
	.clk(clk_clk),
	.d(\M_dc_st_data[16]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[16]~q ),
	.prn(vcc));
defparam \A_dc_st_data[16] .is_wysiwyg = "true";
defparam \A_dc_st_data[16] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[16]~9 (
	.dataa(!\M_dc_st_data[16]~5_combout ),
	.datab(!\A_dc_st_data[16]~q ),
	.datac(!\d_readdata_d1[16]~q ),
	.datad(!\A_st_data[16]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[16]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[16]~9 .extended_lut = "off";
defparam \dc_data_wr_port_data[16]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[16]~9 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[8]~6 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[8]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[8]~6 .extended_lut = "off";
defparam \M_dc_st_data[8]~6 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[8]~6 .shared_arith = "off";

dffeas \A_dc_st_data[8] (
	.clk(clk_clk),
	.d(\M_dc_st_data[8]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[8]~q ),
	.prn(vcc));
defparam \A_dc_st_data[8] .is_wysiwyg = "true";
defparam \A_dc_st_data[8] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[8]~10 (
	.dataa(!\M_dc_st_data[8]~6_combout ),
	.datab(!\A_dc_st_data[8]~q ),
	.datac(!\d_readdata_d1[8]~q ),
	.datad(!\A_st_data[8]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[8]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[8]~10 .extended_lut = "off";
defparam \dc_data_wr_port_data[8]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[8]~10 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[24]~7 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[24]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[24]~7 .extended_lut = "off";
defparam \M_dc_st_data[24]~7 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[24]~7 .shared_arith = "off";

dffeas \A_dc_st_data[24] (
	.clk(clk_clk),
	.d(\M_dc_st_data[24]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[24]~q ),
	.prn(vcc));
defparam \A_dc_st_data[24] .is_wysiwyg = "true";
defparam \A_dc_st_data[24] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[24]~11 (
	.dataa(!\M_dc_st_data[24]~7_combout ),
	.datab(!\A_dc_st_data[24]~q ),
	.datac(!\d_readdata_d1[24]~q ),
	.datad(!\A_st_data[24]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[24]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[24]~11 .extended_lut = "off";
defparam \dc_data_wr_port_data[24]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[24]~11 .shared_arith = "off";

dffeas \i_readdata_d1[8] (
	.clk(clk_clk),
	.d(i_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[8]~q ),
	.prn(vcc));
defparam \i_readdata_d1[8] .is_wysiwyg = "true";
defparam \i_readdata_d1[8] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[2]~8 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.datac(!\M_st_data[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[2]~8 .extended_lut = "off";
defparam \M_dc_st_data[2]~8 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[2]~8 .shared_arith = "off";

dffeas \A_dc_st_data[2] (
	.clk(clk_clk),
	.d(\M_dc_st_data[2]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[2]~q ),
	.prn(vcc));
defparam \A_dc_st_data[2] .is_wysiwyg = "true";
defparam \A_dc_st_data[2] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[2]~12 (
	.dataa(!\M_dc_st_data[2]~8_combout ),
	.datab(!\A_dc_st_data[2]~q ),
	.datac(!\d_readdata_d1[2]~q ),
	.datad(!\A_st_data[2]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[2]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[2]~12 .extended_lut = "off";
defparam \dc_data_wr_port_data[2]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[2]~12 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[18]~9 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[18]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[18]~9 .extended_lut = "off";
defparam \M_dc_st_data[18]~9 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[18]~9 .shared_arith = "off";

dffeas \A_dc_st_data[18] (
	.clk(clk_clk),
	.d(\M_dc_st_data[18]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[18]~q ),
	.prn(vcc));
defparam \A_dc_st_data[18] .is_wysiwyg = "true";
defparam \A_dc_st_data[18] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[18]~13 (
	.dataa(!\M_dc_st_data[18]~9_combout ),
	.datab(!\A_dc_st_data[18]~q ),
	.datac(!\d_readdata_d1[18]~q ),
	.datad(!\A_st_data[18]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[18]~13 .extended_lut = "off";
defparam \dc_data_wr_port_data[18]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[18]~13 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[10]~10 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[10]~10 .extended_lut = "off";
defparam \M_dc_st_data[10]~10 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[10]~10 .shared_arith = "off";

dffeas \A_dc_st_data[10] (
	.clk(clk_clk),
	.d(\M_dc_st_data[10]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[10]~q ),
	.prn(vcc));
defparam \A_dc_st_data[10] .is_wysiwyg = "true";
defparam \A_dc_st_data[10] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[10]~14 (
	.dataa(!\M_dc_st_data[10]~10_combout ),
	.datab(!\A_dc_st_data[10]~q ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\A_st_data[10]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[10]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[10]~14 .extended_lut = "off";
defparam \dc_data_wr_port_data[10]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[10]~14 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[26]~11 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[26]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[26]~11 .extended_lut = "off";
defparam \M_dc_st_data[26]~11 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[26]~11 .shared_arith = "off";

dffeas \A_dc_st_data[26] (
	.clk(clk_clk),
	.d(\M_dc_st_data[26]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[26]~q ),
	.prn(vcc));
defparam \A_dc_st_data[26] .is_wysiwyg = "true";
defparam \A_dc_st_data[26] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[26]~15 (
	.dataa(!\M_dc_st_data[26]~11_combout ),
	.datab(!\A_dc_st_data[26]~q ),
	.datac(!\d_readdata_d1[26]~q ),
	.datad(!\A_st_data[26]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[26]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[26]~15 .extended_lut = "off";
defparam \dc_data_wr_port_data[26]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[26]~15 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[5]~12 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.datac(!\M_st_data[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[5]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[5]~12 .extended_lut = "off";
defparam \M_dc_st_data[5]~12 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[5]~12 .shared_arith = "off";

dffeas \A_dc_st_data[5] (
	.clk(clk_clk),
	.d(\M_dc_st_data[5]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[5]~q ),
	.prn(vcc));
defparam \A_dc_st_data[5] .is_wysiwyg = "true";
defparam \A_dc_st_data[5] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[5]~16 (
	.dataa(!\M_dc_st_data[5]~12_combout ),
	.datab(!\A_dc_st_data[5]~q ),
	.datac(!\d_readdata_d1[5]~q ),
	.datad(!\A_st_data[5]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[5]~16 .extended_lut = "off";
defparam \dc_data_wr_port_data[5]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[5]~16 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[21]~13 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[21]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[21]~13 .extended_lut = "off";
defparam \M_dc_st_data[21]~13 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[21]~13 .shared_arith = "off";

dffeas \A_dc_st_data[21] (
	.clk(clk_clk),
	.d(\M_dc_st_data[21]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[21]~q ),
	.prn(vcc));
defparam \A_dc_st_data[21] .is_wysiwyg = "true";
defparam \A_dc_st_data[21] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[21]~17 (
	.dataa(!\M_dc_st_data[21]~13_combout ),
	.datab(!\A_dc_st_data[21]~q ),
	.datac(!\d_readdata_d1[21]~q ),
	.datad(!\A_st_data[21]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[21]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[21]~17 .extended_lut = "off";
defparam \dc_data_wr_port_data[21]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[21]~17 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[13]~14 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[13]~14 .extended_lut = "off";
defparam \M_dc_st_data[13]~14 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[13]~14 .shared_arith = "off";

dffeas \A_dc_st_data[13] (
	.clk(clk_clk),
	.d(\M_dc_st_data[13]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[13]~q ),
	.prn(vcc));
defparam \A_dc_st_data[13] .is_wysiwyg = "true";
defparam \A_dc_st_data[13] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[13]~18 (
	.dataa(!\M_dc_st_data[13]~14_combout ),
	.datab(!\A_dc_st_data[13]~q ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\A_st_data[13]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[13]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[13]~18 .extended_lut = "off";
defparam \dc_data_wr_port_data[13]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[13]~18 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[29]~15 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[29]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[29]~15 .extended_lut = "off";
defparam \M_dc_st_data[29]~15 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[29]~15 .shared_arith = "off";

dffeas \A_dc_st_data[29] (
	.clk(clk_clk),
	.d(\M_dc_st_data[29]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[29]~q ),
	.prn(vcc));
defparam \A_dc_st_data[29] .is_wysiwyg = "true";
defparam \A_dc_st_data[29] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[29]~19 (
	.dataa(!\M_dc_st_data[29]~15_combout ),
	.datab(!\A_dc_st_data[29]~q ),
	.datac(!\d_readdata_d1[29]~q ),
	.datad(!\A_st_data[29]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[29]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[29]~19 .extended_lut = "off";
defparam \dc_data_wr_port_data[29]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[29]~19 .shared_arith = "off";

dffeas \i_readdata_d1[18] (
	.clk(clk_clk),
	.d(i_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[18]~q ),
	.prn(vcc));
defparam \i_readdata_d1[18] .is_wysiwyg = "true";
defparam \i_readdata_d1[18] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[7]~16 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.datac(!\M_st_data[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[7]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[7]~16 .extended_lut = "off";
defparam \M_dc_st_data[7]~16 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[7]~16 .shared_arith = "off";

dffeas \A_dc_st_data[7] (
	.clk(clk_clk),
	.d(\M_dc_st_data[7]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[7]~q ),
	.prn(vcc));
defparam \A_dc_st_data[7] .is_wysiwyg = "true";
defparam \A_dc_st_data[7] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[7]~20 (
	.dataa(!\M_dc_st_data[7]~16_combout ),
	.datab(!\A_dc_st_data[7]~q ),
	.datac(!\d_readdata_d1[7]~q ),
	.datad(!\A_st_data[7]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[7]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[7]~20 .extended_lut = "off";
defparam \dc_data_wr_port_data[7]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[23]~17 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[23]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[23]~17 .extended_lut = "off";
defparam \M_dc_st_data[23]~17 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[23]~17 .shared_arith = "off";

dffeas \A_dc_st_data[23] (
	.clk(clk_clk),
	.d(\M_dc_st_data[23]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[23]~q ),
	.prn(vcc));
defparam \A_dc_st_data[23] .is_wysiwyg = "true";
defparam \A_dc_st_data[23] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[23]~21 (
	.dataa(!\M_dc_st_data[23]~17_combout ),
	.datab(!\A_dc_st_data[23]~q ),
	.datac(!\d_readdata_d1[23]~q ),
	.datad(!\A_st_data[23]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[23]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[23]~21 .extended_lut = "off";
defparam \dc_data_wr_port_data[23]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[23]~21 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[15]~18 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[15]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[15]~18 .extended_lut = "off";
defparam \M_dc_st_data[15]~18 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[15]~18 .shared_arith = "off";

dffeas \A_dc_st_data[15] (
	.clk(clk_clk),
	.d(\M_dc_st_data[15]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[15]~q ),
	.prn(vcc));
defparam \A_dc_st_data[15] .is_wysiwyg = "true";
defparam \A_dc_st_data[15] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[15]~22 (
	.dataa(!\M_dc_st_data[15]~18_combout ),
	.datab(!\A_dc_st_data[15]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\A_st_data[15]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[15]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[15]~22 .extended_lut = "off";
defparam \dc_data_wr_port_data[15]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[15]~22 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[31]~19 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[31]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[31]~19 .extended_lut = "off";
defparam \M_dc_st_data[31]~19 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[31]~19 .shared_arith = "off";

dffeas \A_dc_st_data[31] (
	.clk(clk_clk),
	.d(\M_dc_st_data[31]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[31]~q ),
	.prn(vcc));
defparam \A_dc_st_data[31] .is_wysiwyg = "true";
defparam \A_dc_st_data[31] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[31]~23 (
	.dataa(!\M_dc_st_data[31]~19_combout ),
	.datab(!\A_dc_st_data[31]~q ),
	.datac(!\d_readdata_d1[31]~q ),
	.datad(!\A_st_data[31]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[31]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[31]~23 .extended_lut = "off";
defparam \dc_data_wr_port_data[31]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[31]~23 .shared_arith = "off";

dffeas \i_readdata_d1[17] (
	.clk(clk_clk),
	.d(i_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[17]~q ),
	.prn(vcc));
defparam \i_readdata_d1[17] .is_wysiwyg = "true";
defparam \i_readdata_d1[17] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[11]~20 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[11]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[11]~20 .extended_lut = "off";
defparam \M_dc_st_data[11]~20 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[11]~20 .shared_arith = "off";

dffeas \A_dc_st_data[11] (
	.clk(clk_clk),
	.d(\M_dc_st_data[11]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[11]~q ),
	.prn(vcc));
defparam \A_dc_st_data[11] .is_wysiwyg = "true";
defparam \A_dc_st_data[11] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[11]~24 (
	.dataa(!\M_dc_st_data[11]~20_combout ),
	.datab(!\A_dc_st_data[11]~q ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\A_st_data[11]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[11]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[11]~24 .extended_lut = "off";
defparam \dc_data_wr_port_data[11]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[11]~24 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[27]~21 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[27]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[27]~21 .extended_lut = "off";
defparam \M_dc_st_data[27]~21 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[27]~21 .shared_arith = "off";

dffeas \A_dc_st_data[27] (
	.clk(clk_clk),
	.d(\M_dc_st_data[27]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[27]~q ),
	.prn(vcc));
defparam \A_dc_st_data[27] .is_wysiwyg = "true";
defparam \A_dc_st_data[27] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[27]~25 (
	.dataa(!\M_dc_st_data[27]~21_combout ),
	.datab(!\A_dc_st_data[27]~q ),
	.datac(!\d_readdata_d1[27]~q ),
	.datad(!\A_st_data[27]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[27]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[27]~25 .extended_lut = "off";
defparam \dc_data_wr_port_data[27]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[27]~25 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[9]~22 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[9]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[9]~22 .extended_lut = "off";
defparam \M_dc_st_data[9]~22 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[9]~22 .shared_arith = "off";

dffeas \A_dc_st_data[9] (
	.clk(clk_clk),
	.d(\M_dc_st_data[9]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[9]~q ),
	.prn(vcc));
defparam \A_dc_st_data[9] .is_wysiwyg = "true";
defparam \A_dc_st_data[9] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[9]~26 (
	.dataa(!\M_dc_st_data[9]~22_combout ),
	.datab(!\A_dc_st_data[9]~q ),
	.datac(!\d_readdata_d1[9]~q ),
	.datad(!\A_st_data[9]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[9]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[9]~26 .extended_lut = "off";
defparam \dc_data_wr_port_data[9]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[9]~26 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[25]~23 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[25]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[25]~23 .extended_lut = "off";
defparam \M_dc_st_data[25]~23 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[25]~23 .shared_arith = "off";

dffeas \A_dc_st_data[25] (
	.clk(clk_clk),
	.d(\M_dc_st_data[25]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[25]~q ),
	.prn(vcc));
defparam \A_dc_st_data[25] .is_wysiwyg = "true";
defparam \A_dc_st_data[25] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[25]~27 (
	.dataa(!\M_dc_st_data[25]~23_combout ),
	.datab(!\A_dc_st_data[25]~q ),
	.datac(!\d_readdata_d1[25]~q ),
	.datad(!\A_st_data[25]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[25]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[25]~27 .extended_lut = "off";
defparam \dc_data_wr_port_data[25]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[25]~27 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[6]~24 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.datac(!\M_st_data[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[6]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[6]~24 .extended_lut = "off";
defparam \M_dc_st_data[6]~24 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[6]~24 .shared_arith = "off";

dffeas \A_dc_st_data[6] (
	.clk(clk_clk),
	.d(\M_dc_st_data[6]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[6]~q ),
	.prn(vcc));
defparam \A_dc_st_data[6] .is_wysiwyg = "true";
defparam \A_dc_st_data[6] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[6]~28 (
	.dataa(!\M_dc_st_data[6]~24_combout ),
	.datab(!\A_dc_st_data[6]~q ),
	.datac(!\d_readdata_d1[6]~q ),
	.datad(!\A_st_data[6]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[6]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[6]~28 .extended_lut = "off";
defparam \dc_data_wr_port_data[6]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[6]~28 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[22]~25 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[22]~25 .extended_lut = "off";
defparam \M_dc_st_data[22]~25 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[22]~25 .shared_arith = "off";

dffeas \A_dc_st_data[22] (
	.clk(clk_clk),
	.d(\M_dc_st_data[22]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[22]~q ),
	.prn(vcc));
defparam \A_dc_st_data[22] .is_wysiwyg = "true";
defparam \A_dc_st_data[22] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[22]~29 (
	.dataa(!\M_dc_st_data[22]~25_combout ),
	.datab(!\A_dc_st_data[22]~q ),
	.datac(!\d_readdata_d1[22]~q ),
	.datad(!\A_st_data[22]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[22]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[22]~29 .extended_lut = "off";
defparam \dc_data_wr_port_data[22]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[22]~29 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[14]~26 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\M_st_data[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[14]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[14]~26 .extended_lut = "off";
defparam \M_dc_st_data[14]~26 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[14]~26 .shared_arith = "off";

dffeas \A_dc_st_data[14] (
	.clk(clk_clk),
	.d(\M_dc_st_data[14]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[14]~q ),
	.prn(vcc));
defparam \A_dc_st_data[14] .is_wysiwyg = "true";
defparam \A_dc_st_data[14] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[14]~30 (
	.dataa(!\M_dc_st_data[14]~26_combout ),
	.datab(!\A_dc_st_data[14]~q ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\A_st_data[14]~q ),
	.datae(!\dc_data_wr_port_data[12]~5_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[14]~30 .extended_lut = "off";
defparam \dc_data_wr_port_data[14]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[14]~30 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[30]~27 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[30]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[30]~27 .extended_lut = "off";
defparam \M_dc_st_data[30]~27 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[30]~27 .shared_arith = "off";

dffeas \A_dc_st_data[30] (
	.clk(clk_clk),
	.d(\M_dc_st_data[30]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[30]~q ),
	.prn(vcc));
defparam \A_dc_st_data[30] .is_wysiwyg = "true";
defparam \A_dc_st_data[30] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[30]~31 (
	.dataa(!\M_dc_st_data[30]~27_combout ),
	.datab(!\A_dc_st_data[30]~q ),
	.datac(!\d_readdata_d1[30]~q ),
	.datad(!\A_st_data[30]~q ),
	.datae(!\dc_data_wr_port_data[31]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[30]~31 .extended_lut = "off";
defparam \dc_data_wr_port_data[30]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[30]~31 .shared_arith = "off";

dffeas \i_readdata_d1[21] (
	.clk(clk_clk),
	.d(i_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[21]~q ),
	.prn(vcc));
defparam \i_readdata_d1[21] .is_wysiwyg = "true";
defparam \i_readdata_d1[21] .power_up = "low";

dffeas \i_readdata_d1[6] (
	.clk(clk_clk),
	.d(i_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[6]~q ),
	.prn(vcc));
defparam \i_readdata_d1[6] .is_wysiwyg = "true";
defparam \i_readdata_d1[6] .power_up = "low";

dffeas \i_readdata_d1[20] (
	.clk(clk_clk),
	.d(i_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[20]~q ),
	.prn(vcc));
defparam \i_readdata_d1[20] .is_wysiwyg = "true";
defparam \i_readdata_d1[20] .power_up = "low";

dffeas \i_readdata_d1[19] (
	.clk(clk_clk),
	.d(i_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[19]~q ),
	.prn(vcc));
defparam \i_readdata_d1[19] .is_wysiwyg = "true";
defparam \i_readdata_d1[19] .power_up = "low";

dffeas \i_readdata_d1[9] (
	.clk(clk_clk),
	.d(i_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[9]~q ),
	.prn(vcc));
defparam \i_readdata_d1[9] .is_wysiwyg = "true";
defparam \i_readdata_d1[9] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[3]~28 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\M_mem_byte_en[0]~q ),
	.datac(!\M_st_data[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[3]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[3]~28 .extended_lut = "off";
defparam \M_dc_st_data[3]~28 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[3]~28 .shared_arith = "off";

dffeas \A_dc_st_data[3] (
	.clk(clk_clk),
	.d(\M_dc_st_data[3]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[3]~q ),
	.prn(vcc));
defparam \A_dc_st_data[3] .is_wysiwyg = "true";
defparam \A_dc_st_data[3] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[3]~32 (
	.dataa(!\M_dc_st_data[3]~28_combout ),
	.datab(!\A_dc_st_data[3]~q ),
	.datac(!\d_readdata_d1[3]~q ),
	.datad(!\A_st_data[3]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[3]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[3]~32 .extended_lut = "off";
defparam \dc_data_wr_port_data[3]~32 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[3]~32 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[19]~29 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[19]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[19]~29 .extended_lut = "off";
defparam \M_dc_st_data[19]~29 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[19]~29 .shared_arith = "off";

dffeas \A_dc_st_data[19] (
	.clk(clk_clk),
	.d(\M_dc_st_data[19]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[19]~q ),
	.prn(vcc));
defparam \A_dc_st_data[19] .is_wysiwyg = "true";
defparam \A_dc_st_data[19] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[19]~33 (
	.dataa(!\M_dc_st_data[19]~29_combout ),
	.datab(!\A_dc_st_data[19]~q ),
	.datac(!\d_readdata_d1[19]~q ),
	.datad(!\A_st_data[19]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[19]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[19]~33 .extended_lut = "off";
defparam \dc_data_wr_port_data[19]~33 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[19]~33 .shared_arith = "off";

cyclonev_lcell_comb ic_tag_clr_valid_bits_nxt(
	.dataa(!rst1),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_clr_valid_bits_nxt.extended_lut = "off";
defparam ic_tag_clr_valid_bits_nxt.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam ic_tag_clr_valid_bits_nxt.shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~7 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_crst~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~7 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~7 .lut_mask = 64'h7777777777777777;
defparam \ic_tag_wraddress_nxt~7 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[0]~8 (
	.dataa(!rst1),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datad(!\ic_tag_wraddress_nxt~6_combout ),
	.datae(!\ic_tag_wraddress_nxt~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[0]~8 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[0]~8 .lut_mask = 64'hBFFFB3FFBFFFB3FF;
defparam \ic_tag_wraddress_nxt[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~9 (
	.dataa(!rst1),
	.datab(!\ic_tag_wraddress_nxt~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~9 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~9 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \ic_tag_wraddress_nxt[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~10 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~4_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~10 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~10 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[1]~10 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[2]~11 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~5_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[2]~11 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[2]~11 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[3]~12 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~3_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[3]~12 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[3]~12 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[3]~12 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[4]~13 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~2_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[4]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[4]~13 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[4]~13 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[4]~13 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[5]~14 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~1_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[5]~14 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[5]~14 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[5]~14 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[6]~15 (
	.dataa(!rst1),
	.datab(!\M_alu_result[11]~q ),
	.datac(!\ic_tag_wraddress_nxt~0_combout ),
	.datad(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datae(!\ic_tag_wraddress_nxt~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[6]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[6]~15 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[6]~15 .lut_mask = 64'hBFFFBF3FBFFFBF3F;
defparam \ic_tag_wraddress_nxt[6]~15 .shared_arith = "off";

dffeas \i_readdata_d1[7] (
	.clk(clk_clk),
	.d(i_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[7]~q ),
	.prn(vcc));
defparam \i_readdata_d1[7] .is_wysiwyg = "true";
defparam \i_readdata_d1[7] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[1]~30 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.datac(!\M_st_data[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[1]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[1]~30 .extended_lut = "off";
defparam \M_dc_st_data[1]~30 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[1]~30 .shared_arith = "off";

dffeas \A_dc_st_data[1] (
	.clk(clk_clk),
	.d(\M_dc_st_data[1]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[1]~q ),
	.prn(vcc));
defparam \A_dc_st_data[1] .is_wysiwyg = "true";
defparam \A_dc_st_data[1] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[1]~34 (
	.dataa(!\M_dc_st_data[1]~30_combout ),
	.datab(!\A_dc_st_data[1]~q ),
	.datac(!\d_readdata_d1[1]~q ),
	.datad(!\A_st_data[1]~q ),
	.datae(!\dc_data_wr_port_data[6]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[1]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[1]~34 .extended_lut = "off";
defparam \dc_data_wr_port_data[1]~34 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[1]~34 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[17]~31 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\M_st_data[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[17]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[17]~31 .extended_lut = "off";
defparam \M_dc_st_data[17]~31 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[17]~31 .shared_arith = "off";

dffeas \A_dc_st_data[17] (
	.clk(clk_clk),
	.d(\M_dc_st_data[17]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[17]~q ),
	.prn(vcc));
defparam \A_dc_st_data[17] .is_wysiwyg = "true";
defparam \A_dc_st_data[17] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[17]~35 (
	.dataa(!\M_dc_st_data[17]~31_combout ),
	.datab(!\A_dc_st_data[17]~q ),
	.datac(!\d_readdata_d1[17]~q ),
	.datad(!\A_st_data[17]~q ),
	.datae(!\dc_data_wr_port_data[18]~3_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[17]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[17]~35 .extended_lut = "off";
defparam \dc_data_wr_port_data[17]~35 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[17]~35 .shared_arith = "off";

dffeas \E_bht_data[0] (
	.clk(clk_clk),
	.d(\D_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_data[0]~q ),
	.prn(vcc));
defparam \E_bht_data[0] .is_wysiwyg = "true";
defparam \E_bht_data[0] .power_up = "low";

cyclonev_lcell_comb E_br_mispredict(
	.dataa(!\E_valid~1_combout ),
	.datab(!\E_bht_data[1]~q ),
	.datac(!\Add24~65_sumout ),
	.datad(!\E_br_result~0_combout ),
	.datae(!\E_br_result~1_combout ),
	.dataf(!\E_ctrl_br_cond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_mispredict~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_br_mispredict.extended_lut = "off";
defparam E_br_mispredict.lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam E_br_mispredict.shared_arith = "off";

dffeas \E_bht_ptr[0] (
	.clk(clk_clk),
	.d(\D_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[0]~q ),
	.prn(vcc));
defparam \E_bht_ptr[0] .is_wysiwyg = "true";
defparam \E_bht_ptr[0] .power_up = "low";

dffeas \E_bht_ptr[1] (
	.clk(clk_clk),
	.d(\D_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[1]~q ),
	.prn(vcc));
defparam \E_bht_ptr[1] .is_wysiwyg = "true";
defparam \E_bht_ptr[1] .power_up = "low";

dffeas \E_bht_ptr[2] (
	.clk(clk_clk),
	.d(\D_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[2]~q ),
	.prn(vcc));
defparam \E_bht_ptr[2] .is_wysiwyg = "true";
defparam \E_bht_ptr[2] .power_up = "low";

dffeas \E_bht_ptr[3] (
	.clk(clk_clk),
	.d(\D_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[3]~q ),
	.prn(vcc));
defparam \E_bht_ptr[3] .is_wysiwyg = "true";
defparam \E_bht_ptr[3] .power_up = "low";

dffeas \E_bht_ptr[4] (
	.clk(clk_clk),
	.d(\D_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[4]~q ),
	.prn(vcc));
defparam \E_bht_ptr[4] .is_wysiwyg = "true";
defparam \E_bht_ptr[4] .power_up = "low";

dffeas \E_bht_ptr[5] (
	.clk(clk_clk),
	.d(\D_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[5]~q ),
	.prn(vcc));
defparam \E_bht_ptr[5] .is_wysiwyg = "true";
defparam \E_bht_ptr[5] .power_up = "low";

dffeas \E_bht_ptr[6] (
	.clk(clk_clk),
	.d(\D_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[6]~q ),
	.prn(vcc));
defparam \E_bht_ptr[6] .is_wysiwyg = "true";
defparam \E_bht_ptr[6] .power_up = "low";

dffeas \E_bht_ptr[7] (
	.clk(clk_clk),
	.d(\D_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[7]~q ),
	.prn(vcc));
defparam \E_bht_ptr[7] .is_wysiwyg = "true";
defparam \E_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \M_br_cond_taken_history[0]~0 (
	.dataa(!\A_div_done~q ),
	.datab(!\A_mem_stall~q ),
	.datac(!\A_mul_stall~q ),
	.datad(!\A_div_stall~0_combout ),
	.datae(!\E_valid~1_combout ),
	.dataf(!\E_ctrl_br_cond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_cond_taken_history[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_cond_taken_history[0]~0 .extended_lut = "off";
defparam \M_br_cond_taken_history[0]~0 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \M_br_cond_taken_history[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ic_fill_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_valid_bits_en(
	.dataa(!\ic_fill_dp_offset_en~0_combout ),
	.datab(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_valid_bits_en.extended_lut = "off";
defparam ic_fill_valid_bits_en.lut_mask = 64'h7777777777777777;
defparam ic_fill_valid_bits_en.shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~1 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~1 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \ic_fill_valid_bits_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~2 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~2 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \ic_fill_valid_bits_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~3 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~3 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~3 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \ic_fill_valid_bits_nxt~3 .shared_arith = "off";

dffeas \D_bht_data[0] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_data[0]~q ),
	.prn(vcc));
defparam \D_bht_data[0] .is_wysiwyg = "true";
defparam \D_bht_data[0] .power_up = "low";

dffeas \D_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[0]~q ),
	.prn(vcc));
defparam \D_bht_ptr[0] .is_wysiwyg = "true";
defparam \D_bht_ptr[0] .power_up = "low";

dffeas \D_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[1]~q ),
	.prn(vcc));
defparam \D_bht_ptr[1] .is_wysiwyg = "true";
defparam \D_bht_ptr[1] .power_up = "low";

dffeas \D_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[2]~q ),
	.prn(vcc));
defparam \D_bht_ptr[2] .is_wysiwyg = "true";
defparam \D_bht_ptr[2] .power_up = "low";

dffeas \D_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[3]~q ),
	.prn(vcc));
defparam \D_bht_ptr[3] .is_wysiwyg = "true";
defparam \D_bht_ptr[3] .power_up = "low";

dffeas \D_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[4]~q ),
	.prn(vcc));
defparam \D_bht_ptr[4] .is_wysiwyg = "true";
defparam \D_bht_ptr[4] .power_up = "low";

dffeas \D_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[5]~q ),
	.prn(vcc));
defparam \D_bht_ptr[5] .is_wysiwyg = "true";
defparam \D_bht_ptr[5] .power_up = "low";

dffeas \D_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[6]~q ),
	.prn(vcc));
defparam \D_bht_ptr[6] .is_wysiwyg = "true";
defparam \D_bht_ptr[6] .power_up = "low";

dffeas \D_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[7]~q ),
	.prn(vcc));
defparam \D_bht_ptr[7] .is_wysiwyg = "true";
defparam \D_bht_ptr[7] .power_up = "low";

dffeas \A_dc_rd_data[7] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[7]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[7] .is_wysiwyg = "true";
defparam \A_dc_rd_data[7] .power_up = "low";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~4 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~4 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~4 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \ic_fill_valid_bits_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~5 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~5 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~5 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \ic_fill_valid_bits_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~6 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~6 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~6 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \ic_fill_valid_bits_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~7 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~7 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~7 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \ic_fill_valid_bits_nxt~7 .shared_arith = "off";

dffeas \A_dc_rd_data[3] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[3] .is_wysiwyg = "true";
defparam \A_dc_rd_data[3] .power_up = "low";

dffeas \F_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[0]~q ),
	.prn(vcc));
defparam \F_bht_ptr[0] .is_wysiwyg = "true";
defparam \F_bht_ptr[0] .power_up = "low";

dffeas \F_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[1]~q ),
	.prn(vcc));
defparam \F_bht_ptr[1] .is_wysiwyg = "true";
defparam \F_bht_ptr[1] .power_up = "low";

dffeas \F_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[2]~q ),
	.prn(vcc));
defparam \F_bht_ptr[2] .is_wysiwyg = "true";
defparam \F_bht_ptr[2] .power_up = "low";

dffeas \F_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[3]~q ),
	.prn(vcc));
defparam \F_bht_ptr[3] .is_wysiwyg = "true";
defparam \F_bht_ptr[3] .power_up = "low";

dffeas \F_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[4]~q ),
	.prn(vcc));
defparam \F_bht_ptr[4] .is_wysiwyg = "true";
defparam \F_bht_ptr[4] .power_up = "low";

dffeas \F_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[5]~q ),
	.prn(vcc));
defparam \F_bht_ptr[5] .is_wysiwyg = "true";
defparam \F_bht_ptr[5] .power_up = "low";

dffeas \F_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[6]~q ),
	.prn(vcc));
defparam \F_bht_ptr[6] .is_wysiwyg = "true";
defparam \F_bht_ptr[6] .power_up = "low";

dffeas \F_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[7]~q ),
	.prn(vcc));
defparam \F_bht_ptr[7] .is_wysiwyg = "true";
defparam \F_bht_ptr[7] .power_up = "low";

dffeas \A_dc_rd_data[1] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[1] .is_wysiwyg = "true";
defparam \A_dc_rd_data[1] .power_up = "low";

dffeas \A_dc_rd_data[4] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[4]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[4] .is_wysiwyg = "true";
defparam \A_dc_rd_data[4] .power_up = "low";

dffeas \A_dc_rd_data[20] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[20]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[20] .is_wysiwyg = "true";
defparam \A_dc_rd_data[20] .power_up = "low";

dffeas \A_dc_rd_data[12] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[12]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[12] .is_wysiwyg = "true";
defparam \A_dc_rd_data[12] .power_up = "low";

dffeas \A_dc_rd_data[28] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[28]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[28] .is_wysiwyg = "true";
defparam \A_dc_rd_data[28] .power_up = "low";

dffeas \A_dc_rd_data[16] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[16]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[16] .is_wysiwyg = "true";
defparam \A_dc_rd_data[16] .power_up = "low";

dffeas \A_dc_rd_data[8] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[8]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[8] .is_wysiwyg = "true";
defparam \A_dc_rd_data[8] .power_up = "low";

dffeas \A_dc_rd_data[24] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[24]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[24] .is_wysiwyg = "true";
defparam \A_dc_rd_data[24] .power_up = "low";

dffeas \A_dc_rd_data[2] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[2] .is_wysiwyg = "true";
defparam \A_dc_rd_data[2] .power_up = "low";

dffeas \A_dc_rd_data[18] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[18]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[18] .is_wysiwyg = "true";
defparam \A_dc_rd_data[18] .power_up = "low";

dffeas \A_dc_rd_data[10] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[10]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[10] .is_wysiwyg = "true";
defparam \A_dc_rd_data[10] .power_up = "low";

dffeas \A_dc_rd_data[26] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[26]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[26] .is_wysiwyg = "true";
defparam \A_dc_rd_data[26] .power_up = "low";

dffeas \A_dc_rd_data[5] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[5]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[5] .is_wysiwyg = "true";
defparam \A_dc_rd_data[5] .power_up = "low";

dffeas \A_dc_rd_data[21] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[21]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[21] .is_wysiwyg = "true";
defparam \A_dc_rd_data[21] .power_up = "low";

dffeas \A_dc_rd_data[13] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[13]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[13] .is_wysiwyg = "true";
defparam \A_dc_rd_data[13] .power_up = "low";

dffeas \A_dc_rd_data[29] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[29]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[29] .is_wysiwyg = "true";
defparam \A_dc_rd_data[29] .power_up = "low";

dffeas \A_dc_rd_data[23] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[23]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[23] .is_wysiwyg = "true";
defparam \A_dc_rd_data[23] .power_up = "low";

dffeas \A_dc_rd_data[15] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[15]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[15] .is_wysiwyg = "true";
defparam \A_dc_rd_data[15] .power_up = "low";

dffeas \A_dc_rd_data[31] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[31]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[31] .is_wysiwyg = "true";
defparam \A_dc_rd_data[31] .power_up = "low";

dffeas \A_dc_rd_data[11] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[11]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[11] .is_wysiwyg = "true";
defparam \A_dc_rd_data[11] .power_up = "low";

dffeas \A_dc_rd_data[27] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[27]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[27] .is_wysiwyg = "true";
defparam \A_dc_rd_data[27] .power_up = "low";

dffeas \A_dc_rd_data[9] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[9]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[9] .is_wysiwyg = "true";
defparam \A_dc_rd_data[9] .power_up = "low";

dffeas \A_dc_rd_data[25] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[25]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[25] .is_wysiwyg = "true";
defparam \A_dc_rd_data[25] .power_up = "low";

dffeas \A_dc_rd_data[6] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[6]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[6] .is_wysiwyg = "true";
defparam \A_dc_rd_data[6] .power_up = "low";

dffeas \A_dc_rd_data[22] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[22]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[22] .is_wysiwyg = "true";
defparam \A_dc_rd_data[22] .power_up = "low";

dffeas \A_dc_rd_data[14] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[14]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[14] .is_wysiwyg = "true";
defparam \A_dc_rd_data[14] .power_up = "low";

dffeas \A_dc_rd_data[30] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[30]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[30] .is_wysiwyg = "true";
defparam \A_dc_rd_data[30] .power_up = "low";

dffeas \A_dc_rd_data[19] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[19]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[19] .is_wysiwyg = "true";
defparam \A_dc_rd_data[19] .power_up = "low";

dffeas \A_dc_rd_data[17] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[17]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[17] .is_wysiwyg = "true";
defparam \A_dc_rd_data[17] .power_up = "low";

cyclonev_lcell_comb \ic_tag_clr_valid_bits~0 (
	.dataa(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ic_tag_clr_valid_bits~0 .shared_arith = "off";

cyclonev_lcell_comb \M_br_mispredict~_wirecell (
	.dataa(!\M_br_mispredict~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_mispredict~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_mispredict~_wirecell .extended_lut = "off";
defparam \M_br_mispredict~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_br_mispredict~_wirecell .shared_arith = "off";

dffeas \d_address_offset_field[2] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[0]~2_combout ),
	.q(d_address_offset_field_2),
	.prn(vcc));
defparam \d_address_offset_field[2] .is_wysiwyg = "true";
defparam \d_address_offset_field[2] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas \d_address_offset_field[0] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[0]~2_combout ),
	.q(d_address_offset_field_0),
	.prn(vcc));
defparam \d_address_offset_field[0] .is_wysiwyg = "true";
defparam \d_address_offset_field[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\d_write_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_address_line_field[0] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_0),
	.prn(vcc));
defparam \d_address_line_field[0] .is_wysiwyg = "true";
defparam \d_address_line_field[0] .power_up = "low";

dffeas \d_address_tag_field[1] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_1),
	.prn(vcc));
defparam \d_address_tag_field[1] .is_wysiwyg = "true";
defparam \d_address_tag_field[1] .power_up = "low";

dffeas \d_address_tag_field[0] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_0),
	.prn(vcc));
defparam \d_address_tag_field[0] .is_wysiwyg = "true";
defparam \d_address_tag_field[0] .power_up = "low";

dffeas \d_address_line_field[5] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_5),
	.prn(vcc));
defparam \d_address_line_field[5] .is_wysiwyg = "true";
defparam \d_address_line_field[5] .power_up = "low";

dffeas \d_address_line_field[4] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_4),
	.prn(vcc));
defparam \d_address_line_field[4] .is_wysiwyg = "true";
defparam \d_address_line_field[4] .power_up = "low";

dffeas \d_address_line_field[3] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_3),
	.prn(vcc));
defparam \d_address_line_field[3] .is_wysiwyg = "true";
defparam \d_address_line_field[3] .power_up = "low";

dffeas \d_address_line_field[2] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[2]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_2),
	.prn(vcc));
defparam \d_address_line_field[2] .is_wysiwyg = "true";
defparam \d_address_line_field[2] .power_up = "low";

dffeas \d_address_line_field[1] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[1]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_1),
	.prn(vcc));
defparam \d_address_line_field[1] .is_wysiwyg = "true";
defparam \d_address_line_field[1] .power_up = "low";

dffeas \d_address_tag_field[5] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_5),
	.prn(vcc));
defparam \d_address_tag_field[5] .is_wysiwyg = "true";
defparam \d_address_tag_field[5] .power_up = "low";

dffeas \d_address_tag_field[4] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_4),
	.prn(vcc));
defparam \d_address_tag_field[4] .is_wysiwyg = "true";
defparam \d_address_tag_field[4] .power_up = "low";

dffeas \d_address_tag_field[3] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_3),
	.prn(vcc));
defparam \d_address_tag_field[3] .is_wysiwyg = "true";
defparam \d_address_tag_field[3] .power_up = "low";

dffeas \d_address_tag_field[2] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[2]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_2),
	.prn(vcc));
defparam \d_address_tag_field[2] .is_wysiwyg = "true";
defparam \d_address_tag_field[2] .power_up = "low";

dffeas \d_address_offset_field[1] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[0]~2_combout ),
	.q(d_address_offset_field_1),
	.prn(vcc));
defparam \d_address_offset_field[1] .is_wysiwyg = "true";
defparam \d_address_offset_field[1] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \ic_fill_tag[4] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_4),
	.prn(vcc));
defparam \ic_fill_tag[4] .is_wysiwyg = "true";
defparam \ic_fill_tag[4] .power_up = "low";

dffeas \ic_fill_tag[3] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_3),
	.prn(vcc));
defparam \ic_fill_tag[3] .is_wysiwyg = "true";
defparam \ic_fill_tag[3] .power_up = "low";

dffeas \ic_fill_tag[2] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_2),
	.prn(vcc));
defparam \ic_fill_tag[2] .is_wysiwyg = "true";
defparam \ic_fill_tag[2] .power_up = "low";

dffeas \ic_fill_tag[1] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_1),
	.prn(vcc));
defparam \ic_fill_tag[1] .is_wysiwyg = "true";
defparam \ic_fill_tag[1] .power_up = "low";

dffeas \ic_fill_tag[0] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_0),
	.prn(vcc));
defparam \ic_fill_tag[0] .is_wysiwyg = "true";
defparam \ic_fill_tag[0] .power_up = "low";

dffeas \ic_fill_line[6] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_6),
	.prn(vcc));
defparam \ic_fill_line[6] .is_wysiwyg = "true";
defparam \ic_fill_line[6] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always138~0_combout ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \ic_fill_line[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_5),
	.prn(vcc));
defparam \ic_fill_line[5] .is_wysiwyg = "true";
defparam \ic_fill_line[5] .power_up = "low";

dffeas \ic_fill_line[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_4),
	.prn(vcc));
defparam \ic_fill_line[4] .is_wysiwyg = "true";
defparam \ic_fill_line[4] .power_up = "low";

dffeas \ic_fill_line[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_3),
	.prn(vcc));
defparam \ic_fill_line[3] .is_wysiwyg = "true";
defparam \ic_fill_line[3] .power_up = "low";

dffeas \ic_fill_line[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_1),
	.prn(vcc));
defparam \ic_fill_line[1] .is_wysiwyg = "true";
defparam \ic_fill_line[1] .power_up = "low";

dffeas \ic_fill_line[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_2),
	.prn(vcc));
defparam \ic_fill_line[2] .is_wysiwyg = "true";
defparam \ic_fill_line[2] .power_up = "low";

dffeas \ic_fill_line[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_0),
	.prn(vcc));
defparam \ic_fill_line[0] .is_wysiwyg = "true";
defparam \ic_fill_line[0] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[7]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \ic_fill_ap_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(ic_fill_ap_offset_0),
	.prn(vcc));
defparam \ic_fill_ap_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[0] .power_up = "low";

dffeas \ic_fill_ap_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(ic_fill_ap_offset_2),
	.prn(vcc));
defparam \ic_fill_ap_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[2] .power_up = "low";

dffeas \ic_fill_ap_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(ic_fill_ap_offset_1),
	.prn(vcc));
defparam \ic_fill_ap_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[1] .power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[20]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[12]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[28]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[16]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[8]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[24]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[18]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[10]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[26]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[5]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[21]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[13]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[29]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[23]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[15]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[31]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[11]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[27]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[9]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[25]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[6]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[22]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[14]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[30]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[19]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\d_writedata_nxt[17]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

cyclonev_lcell_comb av_addr_accepted(
	.dataa(!rst1),
	.datab(!av_begintransfer),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_addr_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam av_addr_accepted.extended_lut = "off";
defparam av_addr_accepted.lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam av_addr_accepted.shared_arith = "off";

cyclonev_lcell_comb \F_iw[14]~10 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[14]~10 .extended_lut = "off";
defparam \F_iw[14]~10 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \F_iw[14]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[16]~6 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~6 .extended_lut = "off";
defparam \F_iw[16]~6 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[16]~6 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

dffeas \E_iw[16] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[16]~q ),
	.prn(vcc));
defparam \E_iw[16] .is_wysiwyg = "true";
defparam \E_iw[16] .power_up = "low";

cyclonev_lcell_comb \F_iw[15]~7 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~7 .extended_lut = "off";
defparam \F_iw[15]~7 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[15]~7 .shared_arith = "off";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas \E_iw[15] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[15]~q ),
	.prn(vcc));
defparam \E_iw[15] .is_wysiwyg = "true";
defparam \E_iw[15] .power_up = "low";

cyclonev_lcell_comb \F_iw[13]~8 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~8 .extended_lut = "off";
defparam \F_iw[13]~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[13]~8 .shared_arith = "off";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

dffeas \E_iw[13] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[13]~q ),
	.prn(vcc));
defparam \E_iw[13] .is_wysiwyg = "true";
defparam \E_iw[13] .power_up = "low";

cyclonev_lcell_comb \E_hbreak_req~0 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_iw[15]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_hbreak_req~0 .extended_lut = "off";
defparam \E_hbreak_req~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_hbreak_req~0 .shared_arith = "off";

dffeas \E_iw[5] (
	.clk(clk_clk),
	.d(\D_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[5]~q ),
	.prn(vcc));
defparam \E_iw[5] .is_wysiwyg = "true";
defparam \E_iw[5] .power_up = "low";

cyclonev_lcell_comb \F_iw[3]~2 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~2 .extended_lut = "off";
defparam \F_iw[3]~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[3]~2 .shared_arith = "off";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

dffeas \E_iw[3] (
	.clk(clk_clk),
	.d(\D_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[3]~q ),
	.prn(vcc));
defparam \E_iw[3] .is_wysiwyg = "true";
defparam \E_iw[3] .power_up = "low";

cyclonev_lcell_comb \F_iw[1]~3 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~3 .extended_lut = "off";
defparam \F_iw[1]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[1]~3 .shared_arith = "off";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

dffeas \E_iw[1] (
	.clk(clk_clk),
	.d(\D_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[1]~q ),
	.prn(vcc));
defparam \E_iw[1] .is_wysiwyg = "true";
defparam \E_iw[1] .power_up = "low";

cyclonev_lcell_comb \F_iw[4]~4 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~4 .extended_lut = "off";
defparam \F_iw[4]~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[4]~4 .shared_arith = "off";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

dffeas \E_iw[4] (
	.clk(clk_clk),
	.d(\D_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[4]~q ),
	.prn(vcc));
defparam \E_iw[4] .is_wysiwyg = "true";
defparam \E_iw[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[2]~5 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[2]~5 .extended_lut = "off";
defparam \F_iw[2]~5 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \F_iw[2]~5 .shared_arith = "off";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas \E_iw[2] (
	.clk(clk_clk),
	.d(\D_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[2]~q ),
	.prn(vcc));
defparam \E_iw[2] .is_wysiwyg = "true";
defparam \E_iw[2] .power_up = "low";

cyclonev_lcell_comb \Equal207~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_iw[1]~q ),
	.datae(!\E_iw[4]~q ),
	.dataf(!\E_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal207~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal207~0 .extended_lut = "off";
defparam \Equal207~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \Equal207~0 .shared_arith = "off";

dffeas \E_iw[14] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[14]~q ),
	.prn(vcc));
defparam \E_iw[14] .is_wysiwyg = "true";
defparam \E_iw[14] .power_up = "low";

cyclonev_lcell_comb \F_iw[12]~11 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[12]~11 .extended_lut = "off";
defparam \F_iw[12]~11 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \F_iw[12]~11 .shared_arith = "off";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

dffeas \E_iw[12] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[12]~q ),
	.prn(vcc));
defparam \E_iw[12] .is_wysiwyg = "true";
defparam \E_iw[12] .power_up = "low";

cyclonev_lcell_comb \F_iw[11]~12 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~12 .extended_lut = "off";
defparam \F_iw[11]~12 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[11]~12 .shared_arith = "off";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

dffeas \E_iw[11] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[11]~q ),
	.prn(vcc));
defparam \E_iw[11] .is_wysiwyg = "true";
defparam \E_iw[11] .power_up = "low";

cyclonev_lcell_comb \E_hbreak_req~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_iw[12]~q ),
	.datac(!\E_iw[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_hbreak_req~1 .extended_lut = "off";
defparam \E_hbreak_req~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \E_hbreak_req~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\E_valid~0_combout ),
	.datac(!hbreak_enabled1),
	.datad(!\wait_for_one_post_bret_inst~q ),
	.datae(!\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\wait_for_one_post_bret_inst~q ),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid~1 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~0_combout ),
	.datac(!\Equal207~0_combout ),
	.datad(!\E_hbreak_req~1_combout ),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~1 .extended_lut = "off";
defparam \E_valid~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \E_valid~1 .shared_arith = "off";

dffeas M_valid_from_E(
	.clk(clk_clk),
	.d(\E_valid~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_valid_from_E~q ),
	.prn(vcc));
defparam M_valid_from_E.is_wysiwyg = "true";
defparam M_valid_from_E.power_up = "low";

dffeas A_valid(
	.clk(clk_clk),
	.d(\M_valid_from_E~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_valid~q ),
	.prn(vcc));
defparam A_valid.is_wysiwyg = "true";
defparam A_valid.power_up = "low";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\Equal169~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_div~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_ctrl_logic~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_div~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_div~0 .extended_lut = "off";
defparam \D_ctrl_div~0 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \D_ctrl_div~0 .shared_arith = "off";

dffeas E_ctrl_div(
	.clk(clk_clk),
	.d(\D_ctrl_div~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_div~q ),
	.prn(vcc));
defparam E_ctrl_div.is_wysiwyg = "true";
defparam E_ctrl_div.power_up = "low";

dffeas M_ctrl_div(
	.clk(clk_clk),
	.d(\E_ctrl_div~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_div~q ),
	.prn(vcc));
defparam M_ctrl_div.is_wysiwyg = "true";
defparam M_ctrl_div.power_up = "low";

dffeas A_ctrl_div(
	.clk(clk_clk),
	.d(\M_ctrl_div~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_div~q ),
	.prn(vcc));
defparam A_ctrl_div.is_wysiwyg = "true";
defparam A_ctrl_div.power_up = "low";

cyclonev_lcell_comb \A_div_do_sub~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\Add11~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_do_sub~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_do_sub~0 .extended_lut = "off";
defparam \A_div_do_sub~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \A_div_do_sub~0 .shared_arith = "off";

dffeas A_div_do_sub(
	.clk(clk_clk),
	.d(\A_div_do_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_do_sub~q ),
	.prn(vcc));
defparam A_div_do_sub.is_wysiwyg = "true";
defparam A_div_do_sub.power_up = "low";

dffeas A_div_accumulate_quotient_bits(
	.clk(clk_clk),
	.d(\A_div_discover_quotient_bits~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_accumulate_quotient_bits~q ),
	.prn(vcc));
defparam A_div_accumulate_quotient_bits.is_wysiwyg = "true";
defparam A_div_accumulate_quotient_bits.power_up = "low";

cyclonev_lcell_comb \A_div_discover_quotient_bits~0 (
	.dataa(!\A_div_accumulate_quotient_bits~q ),
	.datab(!\A_div_norm_cnt[5]~q ),
	.datac(!\A_div_den[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_discover_quotient_bits~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_discover_quotient_bits~0 .extended_lut = "off";
defparam \A_div_discover_quotient_bits~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \A_div_discover_quotient_bits~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[6]~28 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[6]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[6]~28 .extended_lut = "off";
defparam \F_iw[6]~28 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[6]~28 .shared_arith = "off";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_b_is_dst~0 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \F_ctrl_b_is_dst~0 .lut_mask = 64'hFFFFEFFEFFFFEFFE;
defparam \F_ctrl_b_is_dst~0 .shared_arith = "off";

dffeas D_ctrl_b_is_dst(
	.clk(clk_clk),
	.d(\F_ctrl_b_is_dst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_b_is_dst~q ),
	.prn(vcc));
defparam D_ctrl_b_is_dst.is_wysiwyg = "true";
defparam D_ctrl_b_is_dst.power_up = "low";

cyclonev_lcell_comb \F_iw[23]~14 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[23]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[23]~14 .extended_lut = "off";
defparam \F_iw[23]~14 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[23]~14 .shared_arith = "off";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cyclonev_lcell_comb \F_iw[18]~25 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~25 .extended_lut = "off";
defparam \F_iw[18]~25 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \F_iw[18]~25 .shared_arith = "off";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_implicit_dst_retaddr~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[5]~1_combout ),
	.datac(!\F_iw[3]~2_combout ),
	.datad(!\F_iw[4]~4_combout ),
	.datae(!\F_iw[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_retaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_retaddr~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_implicit_dst_retaddr~0 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_retaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_implicit_dst_retaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_retaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_retaddr.power_up = "low";

cyclonev_lcell_comb \F_op_slli~2 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_op_slli~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_op_slli~2 .extended_lut = "off";
defparam \F_op_slli~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \F_op_slli~2 .shared_arith = "off";

cyclonev_lcell_comb \F_op_slli~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(!\F_op_slli~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_op_slli~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_op_slli~0 .extended_lut = "off";
defparam \F_op_slli~0 .lut_mask = 64'hFFBFFFFFFFFFFFFF;
defparam \F_op_slli~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\F_iw[14]~10_combout ),
	.datab(!\F_iw[11]~12_combout ),
	.datac(!\F_iw[16]~6_combout ),
	.datad(!\F_iw[15]~7_combout ),
	.datae(!\F_iw[13]~8_combout ),
	.dataf(!\F_op_slli~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \F_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_eretaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_implicit_dst_eretaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_eretaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_eretaddr.power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[23]~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~0 .extended_lut = "off";
defparam \D_dst_regnum[1]~0 .lut_mask = 64'hBFFF1FFFBFFF1FFF;
defparam \D_dst_regnum[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[25]~17 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[25]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[25]~17 .extended_lut = "off";
defparam \F_iw[25]~17 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[25]~17 .shared_arith = "off";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cyclonev_lcell_comb \F_iw[20]~29 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~29 .extended_lut = "off";
defparam \F_iw[20]~29 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[20]~29 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[3]~3 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\D_iw[20]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~3 .extended_lut = "off";
defparam \D_dst_regnum[3]~3 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[3]~3 .shared_arith = "off";

cyclonev_lcell_comb F_ctrl_ignore_dst(
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[2]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_ignore_dst~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ctrl_ignore_dst.extended_lut = "off";
defparam F_ctrl_ignore_dst.lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam F_ctrl_ignore_dst.shared_arith = "off";

dffeas D_ctrl_ignore_dst(
	.clk(clk_clk),
	.d(\F_ctrl_ignore_dst~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_ignore_dst~q ),
	.prn(vcc));
defparam D_ctrl_ignore_dst.is_wysiwyg = "true";
defparam D_ctrl_ignore_dst.power_up = "low";

cyclonev_lcell_comb \F_iw[22]~15 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[22]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[22]~15 .extended_lut = "off";
defparam \F_iw[22]~15 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[22]~15 .shared_arith = "off";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cyclonev_lcell_comb \F_iw[17]~26 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[17]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[17]~26 .extended_lut = "off";
defparam \F_iw[17]~26 .lut_mask = 64'h7777777777777777;
defparam \F_iw[17]~26 .shared_arith = "off";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[0]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~1 .extended_lut = "off";
defparam \D_dst_regnum[0]~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[24]~18 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[24]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[24]~18 .extended_lut = "off";
defparam \F_iw[24]~18 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[24]~18 .shared_arith = "off";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cyclonev_lcell_comb \F_iw[19]~30 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~30 .extended_lut = "off";
defparam \F_iw[19]~30 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[19]~30 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[2]~2 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[24]~q ),
	.datac(!\D_iw[19]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~2 .extended_lut = "off";
defparam \D_dst_regnum[2]~2 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[26]~16 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[26]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[26]~16 .extended_lut = "off";
defparam \F_iw[26]~16 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[26]~16 .shared_arith = "off";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cyclonev_lcell_comb \F_iw[21]~27 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~27 .extended_lut = "off";
defparam \F_iw[21]~27 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[21]~27 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[4]~4 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[26]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~4 .extended_lut = "off";
defparam \D_dst_regnum[4]~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal297~0 (
	.dataa(!\D_dst_regnum[0]~1_combout ),
	.datab(!\D_dst_regnum[2]~2_combout ),
	.datac(!\D_dst_regnum[3]~3_combout ),
	.datad(!\D_dst_regnum[4]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal297~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal297~0 .extended_lut = "off";
defparam \Equal297~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal297~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_valid~combout ),
	.datab(!\D_ctrl_ignore_dst~q ),
	.datac(!\D_dst_regnum[1]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam D_wr_dst_reg.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_b_cmp_F~0 (
	.dataa(!\D_wr_dst_reg~combout ),
	.datab(!\D_dst_regnum[0]~1_combout ),
	.datac(!\D_dst_regnum[2]~2_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_b_cmp_F~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \D_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \D_regnum_b_cmp_F~1 (
	.dataa(!\D_dst_regnum[4]~4_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \D_regnum_b_cmp_F~1 .lut_mask = 64'h6666666666666666;
defparam \D_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_b_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\D_dst_regnum[3]~3_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datae(!\D_regnum_b_cmp_F~0_combout ),
	.dataf(!\D_regnum_b_cmp_F~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_b_cmp_F.extended_lut = "off";
defparam D_regnum_b_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_b_cmp_F.shared_arith = "off";

dffeas E_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_b_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_stall~combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_b_cmp_D.is_wysiwyg = "true";
defparam E_regnum_b_cmp_D.power_up = "low";

dffeas \E_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[2]~q ),
	.prn(vcc));
defparam \E_dst_regnum[2] .is_wysiwyg = "true";
defparam \E_dst_regnum[2] .power_up = "low";

cyclonev_lcell_comb E_hbreak_req(
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~0_combout ),
	.datac(!\Equal207~0_combout ),
	.datad(!\E_hbreak_req~1_combout ),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_hbreak_req.extended_lut = "off";
defparam E_hbreak_req.lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam E_hbreak_req.shared_arith = "off";

dffeas \D_bht_data[1] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_data[1]~q ),
	.prn(vcc));
defparam \D_bht_data[1] .is_wysiwyg = "true";
defparam \D_bht_data[1] .power_up = "low";

dffeas \E_bht_data[1] (
	.clk(clk_clk),
	.d(\D_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_data[1]~q ),
	.prn(vcc));
defparam \E_bht_data[1] .is_wysiwyg = "true";
defparam \E_bht_data[1] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_cmp~3 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~3 .extended_lut = "off";
defparam \D_ctrl_cmp~3 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \D_ctrl_cmp~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_iw[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(gnd),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'hAFFAFAAFFAAFAFFA;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\D_ctrl_cmp~3_combout ),
	.datac(!\D_ctrl_alu_subtract~0_combout ),
	.datad(!\D_ctrl_alu_subtract~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~2 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_alu_subtract~2 .shared_arith = "off";

dffeas E_ctrl_alu_subtract(
	.clk(clk_clk),
	.d(\D_ctrl_alu_subtract~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_alu_subtract~q ),
	.prn(vcc));
defparam E_ctrl_alu_subtract.is_wysiwyg = "true";
defparam E_ctrl_alu_subtract.power_up = "low";

cyclonev_lcell_comb \Equal152~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~1 .extended_lut = "off";
defparam \Equal152~1 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal152~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~3 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~3 .extended_lut = "off";
defparam \Equal152~3 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal152~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~0 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~0 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \D_ctrl_alu_signed_comparison~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~1 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\Equal152~1_combout ),
	.datac(!\Equal152~3_combout ),
	.datad(!\D_ctrl_alu_signed_comparison~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~1 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_alu_signed_comparison~1 .shared_arith = "off";

dffeas E_ctrl_alu_signed_comparison(
	.clk(clk_clk),
	.d(\D_ctrl_alu_signed_comparison~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_alu_signed_comparison~q ),
	.prn(vcc));
defparam E_ctrl_alu_signed_comparison.is_wysiwyg = "true";
defparam E_ctrl_alu_signed_comparison.power_up = "low";

cyclonev_lcell_comb \F_op_slli~3 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_op_slli~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_op_slli~3 .extended_lut = "off";
defparam \F_op_slli~3 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \F_op_slli~3 .shared_arith = "off";

cyclonev_lcell_comb \F_op_slli~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(!\F_op_slli~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_op_slli~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_op_slli~1 .extended_lut = "off";
defparam \F_op_slli~1 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \F_op_slli~1 .shared_arith = "off";

cyclonev_lcell_comb F_ctrl_src2_choose_imm(
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[2]~5_combout ),
	.datad(!\F_ctrl_b_is_dst~0_combout ),
	.datae(!\F_op_slli~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_src2_choose_imm~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ctrl_src2_choose_imm.extended_lut = "off";
defparam F_ctrl_src2_choose_imm.lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam F_ctrl_src2_choose_imm.shared_arith = "off";

dffeas D_ctrl_src2_choose_imm(
	.clk(clk_clk),
	.d(\F_ctrl_src2_choose_imm~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_src2_choose_imm~q ),
	.prn(vcc));
defparam D_ctrl_src2_choose_imm.is_wysiwyg = "true";
defparam D_ctrl_src2_choose_imm.power_up = "low";

cyclonev_lcell_comb \Equal299~0 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\D_iw[26]~q ),
	.datad(!\D_iw[25]~q ),
	.datae(!\D_iw[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal299~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal299~0 .extended_lut = "off";
defparam \Equal299~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal299~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~2 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~2 .extended_lut = "off";
defparam \D_src2_reg[29]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \D_src2_reg[29]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~30 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~30 .extended_lut = "off";
defparam \D_src2_reg[0]~30 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_src2_reg[0]~30 .shared_arith = "off";

cyclonev_lcell_comb \Equal90~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal90~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal90~0 .extended_lut = "off";
defparam \Equal90~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal90~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_ctrl_logic~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~2 (
	.dataa(!\D_iw[3]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\Equal90~0_combout ),
	.datad(!\D_ctrl_logic~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~2 .extended_lut = "off";
defparam \D_ctrl_logic~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_logic~2 .shared_arith = "off";

dffeas E_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_logic~q ),
	.prn(vcc));
defparam E_ctrl_logic.is_wysiwyg = "true";
defparam E_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \Equal103~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal103~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal103~0 .extended_lut = "off";
defparam \Equal103~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal103~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~0 .extended_lut = "off";
defparam \Equal152~0 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \Equal152~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~2 .extended_lut = "off";
defparam \D_ctrl_retaddr~2 .lut_mask = 64'hBFFFFBFFFFFFFFFF;
defparam \D_ctrl_retaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\Equal169~0_combout ),
	.datac(!\Equal103~0_combout ),
	.datad(!\Equal152~0_combout ),
	.datae(!\D_ctrl_retaddr~2_combout ),
	.dataf(!\D_ctrl_retaddr~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

dffeas E_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_retaddr~q ),
	.prn(vcc));
defparam E_ctrl_retaddr.is_wysiwyg = "true";
defparam E_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \D_ctrl_cmp~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~2 .extended_lut = "off";
defparam \D_ctrl_cmp~2 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \D_ctrl_cmp~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~0 .extended_lut = "off";
defparam \D_ctrl_cmp~0 .lut_mask = 64'hFFFFFFFFFFEBFFBE;
defparam \D_ctrl_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~1 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\D_ctrl_cmp~3_combout ),
	.datac(!\D_ctrl_cmp~2_combout ),
	.datad(!\D_ctrl_cmp~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~1 .extended_lut = "off";
defparam \D_ctrl_cmp~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_cmp~1 .shared_arith = "off";

dffeas E_ctrl_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_cmp~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_cmp~q ),
	.prn(vcc));
defparam E_ctrl_cmp.is_wysiwyg = "true";
defparam E_ctrl_cmp.power_up = "low";

cyclonev_lcell_comb \E_alu_result~0 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_ctrl_cmp~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~0 .extended_lut = "off";
defparam \E_alu_result~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\Equal169~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[1]~0 .extended_lut = "off";
defparam \D_logic_op_raw[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~2 .extended_lut = "off";
defparam \Equal152~2 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Equal152~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~4 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~4 .extended_lut = "off";
defparam \Equal152~4 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal152~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~5 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~5 .extended_lut = "off";
defparam \Equal152~5 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal152~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~0 (
	.dataa(!\Equal152~1_combout ),
	.datab(!\Equal152~2_combout ),
	.datac(!\Equal152~4_combout ),
	.datad(!\Equal152~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~0 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_alu_force_xor~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(!\D_ctrl_alu_force_xor~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~1 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~1 .lut_mask = 64'hFFFFFFFFFFB7FF7B;
defparam \D_ctrl_alu_force_xor~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_ctrl_alu_force_xor~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~2 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_alu_force_xor~2 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[1]~0 (
	.dataa(!\D_logic_op_raw[1]~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[1]~0 .extended_lut = "off";
defparam \D_logic_op[1]~0 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[1]~0 .shared_arith = "off";

dffeas \E_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_logic_op[1]~q ),
	.prn(vcc));
defparam \E_logic_op[1] .is_wysiwyg = "true";
defparam \E_logic_op[1] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\Equal169~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[0]~1 .extended_lut = "off";
defparam \D_logic_op_raw[0]~1 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[0]~1 (
	.dataa(!\D_ctrl_alu_force_xor~2_combout ),
	.datab(!\D_logic_op_raw[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[0]~1 .extended_lut = "off";
defparam \D_logic_op[0]~1 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[0]~1 .shared_arith = "off";

dffeas \E_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_logic_op[0]~q ),
	.prn(vcc));
defparam \E_logic_op[0] .is_wysiwyg = "true";
defparam \E_logic_op[0] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~31 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[31]~q ),
	.datae(!\E_src1[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~31 .extended_lut = "off";
defparam \E_alu_result~31 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~37_sumout ),
	.datac(!\E_alu_result~31_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31] .extended_lut = "off";
defparam \E_alu_result[31] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[31] .shared_arith = "off";

dffeas \M_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[31]~q ),
	.prn(vcc));
defparam \M_alu_result[31] .is_wysiwyg = "true";
defparam \M_alu_result[31] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_late_result~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~3 .extended_lut = "off";
defparam \D_ctrl_late_result~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_late_result~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mul_lsw~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\Equal169~0_combout ),
	.datae(!\Equal90~0_combout ),
	.dataf(!\D_ctrl_late_result~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mul_lsw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mul_lsw~0 .extended_lut = "off";
defparam \D_ctrl_mul_lsw~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \D_ctrl_mul_lsw~0 .shared_arith = "off";

dffeas E_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\D_ctrl_mul_lsw~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam E_ctrl_mul_lsw.is_wysiwyg = "true";
defparam E_ctrl_mul_lsw.power_up = "low";

dffeas M_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\E_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam M_ctrl_mul_lsw.is_wysiwyg = "true";
defparam M_ctrl_mul_lsw.power_up = "low";

dffeas A_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\M_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam A_ctrl_mul_lsw.is_wysiwyg = "true";
defparam A_ctrl_mul_lsw.power_up = "low";

cyclonev_lcell_comb \E_op_rdctl~0 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_iw[11]~q ),
	.datac(!\E_iw[16]~q ),
	.datad(!\E_iw[15]~q ),
	.datae(!\E_iw[13]~q ),
	.dataf(!\Equal207~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_rdctl~0 .extended_lut = "off";
defparam \E_op_rdctl~0 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \E_op_rdctl~0 .shared_arith = "off";

cyclonev_lcell_comb E_op_rdctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_rdctl.extended_lut = "off";
defparam E_op_rdctl.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam E_op_rdctl.shared_arith = "off";

dffeas M_ctrl_rdctl_inst(
	.clk(clk_clk),
	.d(\E_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_rdctl_inst~q ),
	.prn(vcc));
defparam M_ctrl_rdctl_inst.is_wysiwyg = "true";
defparam M_ctrl_rdctl_inst.power_up = "low";

cyclonev_lcell_comb \M_ctrl_mem_nxt~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_mem_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_mem_nxt~0 .extended_lut = "off";
defparam \M_ctrl_mem_nxt~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_ctrl_mem_nxt~0 .shared_arith = "off";

dffeas M_ctrl_mem(
	.clk(clk_clk),
	.d(\M_ctrl_mem_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_mem~q ),
	.prn(vcc));
defparam M_ctrl_mem.is_wysiwyg = "true";
defparam M_ctrl_mem.power_up = "low";

dffeas \A_inst_result[31] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(\M_alu_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[31]~q ),
	.prn(vcc));
defparam \A_inst_result[31] .is_wysiwyg = "true";
defparam \A_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot.is_wysiwyg = "true";
defparam E_ctrl_shift_rot.power_up = "low";

dffeas M_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\E_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_shift_rot~q ),
	.prn(vcc));
defparam M_ctrl_shift_rot.is_wysiwyg = "true";
defparam M_ctrl_shift_rot.power_up = "low";

dffeas A_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\M_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_shift_rot~q ),
	.prn(vcc));
defparam A_ctrl_shift_rot.is_wysiwyg = "true";
defparam A_ctrl_shift_rot.power_up = "low";

dffeas \E_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[4]~q ),
	.prn(vcc));
defparam \E_dst_regnum[4] .is_wysiwyg = "true";
defparam \E_dst_regnum[4] .power_up = "low";

dffeas \M_dst_regnum[4] (
	.clk(clk_clk),
	.d(\E_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[4]~q ),
	.prn(vcc));
defparam \M_dst_regnum[4] .is_wysiwyg = "true";
defparam \M_dst_regnum[4] .power_up = "low";

dffeas M_wr_dst_reg_from_E(
	.clk(clk_clk),
	.d(\E_wr_dst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_wr_dst_reg_from_E~q ),
	.prn(vcc));
defparam M_wr_dst_reg_from_E.is_wysiwyg = "true";
defparam M_wr_dst_reg_from_E.power_up = "low";

dffeas \E_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[0]~q ),
	.prn(vcc));
defparam \E_dst_regnum[0] .is_wysiwyg = "true";
defparam \E_dst_regnum[0] .power_up = "low";

dffeas \M_dst_regnum[0] (
	.clk(clk_clk),
	.d(\E_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[0]~q ),
	.prn(vcc));
defparam \M_dst_regnum[0] .is_wysiwyg = "true";
defparam \M_dst_regnum[0] .power_up = "low";

dffeas \E_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[1]~q ),
	.prn(vcc));
defparam \E_dst_regnum[1] .is_wysiwyg = "true";
defparam \E_dst_regnum[1] .power_up = "low";

dffeas \M_dst_regnum[1] (
	.clk(clk_clk),
	.d(\E_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[1]~q ),
	.prn(vcc));
defparam \M_dst_regnum[1] .is_wysiwyg = "true";
defparam \M_dst_regnum[1] .power_up = "low";

cyclonev_lcell_comb \M_regnum_b_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\M_wr_dst_reg_from_E~q ),
	.datad(!\M_dst_regnum[0]~q ),
	.datae(!\M_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \M_regnum_b_cmp_F~0 .shared_arith = "off";

dffeas \M_dst_regnum[2] (
	.clk(clk_clk),
	.d(\E_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[2]~q ),
	.prn(vcc));
defparam \M_dst_regnum[2] .is_wysiwyg = "true";
defparam \M_dst_regnum[2] .power_up = "low";

dffeas \E_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[3]~q ),
	.prn(vcc));
defparam \E_dst_regnum[3] .is_wysiwyg = "true";
defparam \E_dst_regnum[3] .power_up = "low";

dffeas \M_dst_regnum[3] (
	.clk(clk_clk),
	.d(\E_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[3]~q ),
	.prn(vcc));
defparam \M_dst_regnum[3] .is_wysiwyg = "true";
defparam \M_dst_regnum[3] .power_up = "low";

cyclonev_lcell_comb \M_regnum_b_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\M_dst_regnum[2]~q ),
	.datad(!\M_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_b_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\M_regnum_b_cmp_F~0_combout ),
	.datad(!\M_regnum_b_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_b_cmp_F.extended_lut = "off";
defparam M_regnum_b_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam M_regnum_b_cmp_F.shared_arith = "off";

dffeas A_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_b_cmp_F~combout ),
	.asdata(\M_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\A_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_b_cmp_D.is_wysiwyg = "true";
defparam A_regnum_b_cmp_D.power_up = "low";

dffeas \A_dst_regnum_from_M[4] (
	.clk(clk_clk),
	.d(\M_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[4]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[4] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[4] .power_up = "low";

dffeas A_wr_dst_reg_from_M(
	.clk(clk_clk),
	.d(\M_wr_dst_reg_from_E~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_wr_dst_reg_from_M~q ),
	.prn(vcc));
defparam A_wr_dst_reg_from_M.is_wysiwyg = "true";
defparam A_wr_dst_reg_from_M.power_up = "low";

dffeas \A_dst_regnum_from_M[0] (
	.clk(clk_clk),
	.d(\M_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[0]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[0] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[0] .power_up = "low";

dffeas \A_dst_regnum_from_M[1] (
	.clk(clk_clk),
	.d(\M_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[1]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[1] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[1] .power_up = "low";

cyclonev_lcell_comb \A_regnum_b_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\A_wr_dst_reg_from_M~q ),
	.datad(!\A_dst_regnum_from_M[0]~q ),
	.datae(!\A_dst_regnum_from_M[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \A_regnum_b_cmp_F~0 .shared_arith = "off";

dffeas \A_dst_regnum_from_M[2] (
	.clk(clk_clk),
	.d(\M_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[2]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[2] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[2] .power_up = "low";

dffeas \A_dst_regnum_from_M[3] (
	.clk(clk_clk),
	.d(\M_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[3]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[3] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[3] .power_up = "low";

cyclonev_lcell_comb \A_regnum_b_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\A_dst_regnum_from_M[2]~q ),
	.datad(!\A_dst_regnum_from_M[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_b_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\A_dst_regnum_from_M[4]~q ),
	.datac(!\A_regnum_b_cmp_F~0_combout ),
	.datad(!\A_regnum_b_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_b_cmp_F.extended_lut = "off";
defparam A_regnum_b_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam A_regnum_b_cmp_F.shared_arith = "off";

dffeas W_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_b_cmp_F~combout ),
	.asdata(\A_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(vcc),
	.q(\W_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_b_cmp_D.is_wysiwyg = "true";
defparam W_regnum_b_cmp_D.power_up = "low";

cyclonev_lcell_comb \D_src2_reg[29]~4 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\M_regnum_b_cmp_D~q ),
	.datac(!\A_regnum_b_cmp_D~q ),
	.datad(!\W_regnum_b_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~4 .extended_lut = "off";
defparam \D_src2_reg[29]~4 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \D_src2_reg[29]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~3 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\M_regnum_b_cmp_D~q ),
	.datac(!\A_regnum_b_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~3 .extended_lut = "off";
defparam \D_src2_reg[29]~3 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_src2_reg[29]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[3]~13 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~13 .extended_lut = "off";
defparam \D_src2_reg[3]~13 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_src2_reg[3]~13 .shared_arith = "off";

dffeas \A_mul_partial_prod[15] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[15]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[15] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[15] .power_up = "low";

dffeas \A_mul_partial_prod[14] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[14]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[14] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[14] .power_up = "low";

dffeas \A_mul_partial_prod[13] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[13]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[13] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[13] .power_up = "low";

dffeas \A_mul_partial_prod[12] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[12]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[12] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[12] .power_up = "low";

dffeas \A_mul_partial_prod[11] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[11]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[11] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[11] .power_up = "low";

dffeas \A_mul_partial_prod[10] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[10]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[10] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[10] .power_up = "low";

dffeas \A_mul_partial_prod[9] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[9]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[9] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[9] .power_up = "low";

dffeas \A_mul_partial_prod[8] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[8]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[8] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[8] .power_up = "low";

dffeas \A_mul_partial_prod[7] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[7]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[7] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[7] .power_up = "low";

dffeas \A_mul_partial_prod[6] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[6]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[6] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[6] .power_up = "low";

dffeas \A_mul_partial_prod[5] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[5]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[5] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[5] .power_up = "low";

dffeas \A_mul_partial_prod[4] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[4]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[4] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[4] .power_up = "low";

dffeas \A_mul_partial_prod[3] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[3]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[3] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[3] .power_up = "low";

dffeas \A_mul_partial_prod[2] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[2]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[2] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[2] .power_up = "low";

dffeas \A_mul_partial_prod[1] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[1]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[1] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[1] .power_up = "low";

dffeas \A_mul_partial_prod[0] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[0]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[0] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[0] .power_up = "low";

cyclonev_lcell_comb \Add26~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[0]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~5_sumout ),
	.cout(\Add26~6 ),
	.shareout());
defparam \Add26~5 .extended_lut = "off";
defparam \Add26~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~5 .shared_arith = "off";

cyclonev_lcell_comb \E_ld_st_dcache_management_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add24~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_dcache_management_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_dcache_management_bus~0 .extended_lut = "off";
defparam \E_ld_st_dcache_management_bus~0 .lut_mask = 64'h5FFF3FFFFFFFFFFF;
defparam \E_ld_st_dcache_management_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_bypass_or_dcache_management(
	.clk(clk_clk),
	.d(\E_ld_st_dcache_management_bus~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_bypass_or_dcache_management~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_bypass_or_dcache_management.is_wysiwyg = "true";
defparam M_ctrl_ld_st_bypass_or_dcache_management.power_up = "low";

cyclonev_lcell_comb \A_mem_stall_nxt~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_ld_st_bypass_or_dcache_management~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~0 .extended_lut = "off";
defparam \A_mem_stall_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_mem_stall_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_st_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(!\Add24~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_bus~0 .extended_lut = "off";
defparam \E_st_bus~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_st_bus~0 .shared_arith = "off";

dffeas M_ctrl_st_bypass(
	.clk(clk_clk),
	.d(\E_st_bus~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st_bypass~q ),
	.prn(vcc));
defparam M_ctrl_st_bypass.is_wysiwyg = "true";
defparam M_ctrl_st_bypass.power_up = "low";

dffeas \A_inst_result[16] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.asdata(\M_alu_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[16]~q ),
	.prn(vcc));
defparam \A_inst_result[16] .is_wysiwyg = "true";
defparam \A_inst_result[16] .power_up = "low";

dffeas \A_mul_partial_prod[16] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[16]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[16] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[16] .power_up = "low";

cyclonev_lcell_comb \Add26~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[15]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[15]~q ),
	.datag(gnd),
	.cin(\Add26~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~49_sumout ),
	.cout(\Add26~50 ),
	.shareout());
defparam \Add26~49 .extended_lut = "off";
defparam \Add26~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~49 .shared_arith = "off";

cyclonev_lcell_comb \Add26~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[16]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[16]~q ),
	.datag(gnd),
	.cin(\Add26~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~45_sumout ),
	.cout(\Add26~46 ),
	.shareout());
defparam \Add26~45 .extended_lut = "off";
defparam \Add26~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~45 .shared_arith = "off";

dffeas \A_mul_result[16] (
	.clk(clk_clk),
	.d(\Add26~45_sumout ),
	.asdata(\A_mul_partial_prod[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[16]~q ),
	.prn(vcc));
defparam \A_mul_result[16] .is_wysiwyg = "true";
defparam \A_mul_result[16] .power_up = "low";

cyclonev_lcell_comb \F_iw[7]~32 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[7]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[7]~32 .extended_lut = "off";
defparam \F_iw[7]~32 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[7]~32 .shared_arith = "off";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

dffeas \d_readdata_d1[1] (
	.clk(clk_clk),
	.d(d_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[1]~q ),
	.prn(vcc));
defparam \d_readdata_d1[1] .is_wysiwyg = "true";
defparam \d_readdata_d1[1] .power_up = "low";

dffeas \d_readdata_d1[17] (
	.clk(clk_clk),
	.d(d_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[17]~q ),
	.prn(vcc));
defparam \d_readdata_d1[17] .is_wysiwyg = "true";
defparam \d_readdata_d1[17] .power_up = "low";

dffeas \d_readdata_d1[9] (
	.clk(clk_clk),
	.d(d_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[9]~q ),
	.prn(vcc));
defparam \d_readdata_d1[9] .is_wysiwyg = "true";
defparam \d_readdata_d1[9] .power_up = "low";

dffeas \d_readdata_d1[25] (
	.clk(clk_clk),
	.d(d_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[25]~q ),
	.prn(vcc));
defparam \d_readdata_d1[25] .is_wysiwyg = "true";
defparam \d_readdata_d1[25] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_ld8_ld16~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_ld8_ld16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_ld8_ld16~0 .extended_lut = "off";
defparam \E_ctrl_ld8_ld16~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \E_ctrl_ld8_ld16~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal182~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_ctrl_ld8_ld16~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal182~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal182~0 .extended_lut = "off";
defparam \Equal182~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal182~0 .shared_arith = "off";

dffeas M_ctrl_ld8(
	.clk(clk_clk),
	.d(\Equal182~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld8~q ),
	.prn(vcc));
defparam M_ctrl_ld8.is_wysiwyg = "true";
defparam M_ctrl_ld8.power_up = "low";

cyclonev_lcell_comb \Equal185~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal185~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal185~0 .extended_lut = "off";
defparam \Equal185~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Equal185~0 .shared_arith = "off";

dffeas M_ctrl_ld16(
	.clk(clk_clk),
	.d(\Equal185~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld16.power_up = "low";

cyclonev_lcell_comb \M_ld_align_sh16~0 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\M_ctrl_ld8~q ),
	.datac(!\M_ctrl_ld16~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_sh16~0 .extended_lut = "off";
defparam \M_ld_align_sh16~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_ld_align_sh16~0 .shared_arith = "off";

dffeas A_ld_align_sh16(
	.clk(clk_clk),
	.d(\M_ld_align_sh16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_sh16~q ),
	.prn(vcc));
defparam A_ld_align_sh16.is_wysiwyg = "true";
defparam A_ld_align_sh16.power_up = "low";

dffeas \E_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_compare_op[0]~q ),
	.prn(vcc));
defparam \E_compare_op[0] .is_wysiwyg = "true";
defparam \E_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~31 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(gnd),
	.datad(!\Equal299~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~31 .extended_lut = "off";
defparam \D_src2_reg[0]~31 .lut_mask = 64'hFFBBFFBBFFBBFFBB;
defparam \D_src2_reg[0]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~17 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[29]~9_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~17 .extended_lut = "off";
defparam \E_alu_result~17 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~17_combout ),
	.datac(!\Add24~81_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29] .extended_lut = "off";
defparam \E_alu_result[29] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[29] .shared_arith = "off";

dffeas \M_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[29]~q ),
	.prn(vcc));
defparam \M_alu_result[29] .is_wysiwyg = "true";
defparam \M_alu_result[29] .power_up = "low";

dffeas \A_inst_result[29] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(\M_alu_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[29]~q ),
	.prn(vcc));
defparam \A_inst_result[29] .is_wysiwyg = "true";
defparam \A_inst_result[29] .power_up = "low";

dffeas \A_mul_partial_prod[29] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[29]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[29] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[29] .power_up = "low";

dffeas \A_mul_partial_prod[28] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[28]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[28] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[28] .power_up = "low";

dffeas \A_mul_partial_prod[27] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[27]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[27] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[27] .power_up = "low";

dffeas \A_mul_partial_prod[26] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[26]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[26] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[26] .power_up = "low";

dffeas \A_mul_partial_prod[25] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[25]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[25] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[25] .power_up = "low";

dffeas \A_mul_partial_prod[24] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[24]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[24] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[24] .power_up = "low";

dffeas \A_mul_partial_prod[23] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[23]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[23] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[23] .power_up = "low";

dffeas \A_mul_partial_prod[22] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[22]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[22] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[22] .power_up = "low";

dffeas \A_mul_partial_prod[21] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[21]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[21] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[21] .power_up = "low";

dffeas \A_mul_partial_prod[20] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[20]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[20] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[20] .power_up = "low";

dffeas \A_mul_partial_prod[19] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[19]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[19] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[19] .power_up = "low";

dffeas \A_mul_partial_prod[18] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[18]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[18] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[18] .power_up = "low";

dffeas \A_mul_partial_prod[17] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[17]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[17] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[17] .power_up = "low";

cyclonev_lcell_comb \Add26~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[17]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[17]~q ),
	.datag(gnd),
	.cin(\Add26~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~97_sumout ),
	.cout(\Add26~98 ),
	.shareout());
defparam \Add26~97 .extended_lut = "off";
defparam \Add26~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~97 .shared_arith = "off";

dffeas \A_mul_result[17] (
	.clk(clk_clk),
	.d(\Add26~97_sumout ),
	.asdata(\A_mul_partial_prod[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[17]~q ),
	.prn(vcc));
defparam \A_mul_result[17] .is_wysiwyg = "true";
defparam \A_mul_result[17] .power_up = "low";

cyclonev_lcell_comb \Add26~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[18]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[18]~q ),
	.datag(gnd),
	.cin(\Add26~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~113_sumout ),
	.cout(\Add26~114 ),
	.shareout());
defparam \Add26~113 .extended_lut = "off";
defparam \Add26~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~113 .shared_arith = "off";

dffeas \A_mul_result[18] (
	.clk(clk_clk),
	.d(\Add26~113_sumout ),
	.asdata(\A_mul_partial_prod[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[18]~q ),
	.prn(vcc));
defparam \A_mul_result[18] .is_wysiwyg = "true";
defparam \A_mul_result[18] .power_up = "low";

cyclonev_lcell_comb \Add26~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[19]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[19]~q ),
	.datag(gnd),
	.cin(\Add26~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~89_sumout ),
	.cout(\Add26~90 ),
	.shareout());
defparam \Add26~89 .extended_lut = "off";
defparam \Add26~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~89 .shared_arith = "off";

dffeas \A_mul_result[19] (
	.clk(clk_clk),
	.d(\Add26~89_sumout ),
	.asdata(\A_mul_partial_prod[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[19]~q ),
	.prn(vcc));
defparam \A_mul_result[19] .is_wysiwyg = "true";
defparam \A_mul_result[19] .power_up = "low";

cyclonev_lcell_comb \Add26~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[20]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[20]~q ),
	.datag(gnd),
	.cin(\Add26~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~109_sumout ),
	.cout(\Add26~110 ),
	.shareout());
defparam \Add26~109 .extended_lut = "off";
defparam \Add26~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~109 .shared_arith = "off";

dffeas \A_mul_result[20] (
	.clk(clk_clk),
	.d(\Add26~109_sumout ),
	.asdata(\A_mul_partial_prod[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[20]~q ),
	.prn(vcc));
defparam \A_mul_result[20] .is_wysiwyg = "true";
defparam \A_mul_result[20] .power_up = "low";

cyclonev_lcell_comb \Add26~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[21]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[21]~q ),
	.datag(gnd),
	.cin(\Add26~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~105_sumout ),
	.cout(\Add26~106 ),
	.shareout());
defparam \Add26~105 .extended_lut = "off";
defparam \Add26~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~105 .shared_arith = "off";

dffeas \A_mul_result[21] (
	.clk(clk_clk),
	.d(\Add26~105_sumout ),
	.asdata(\A_mul_partial_prod[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[21]~q ),
	.prn(vcc));
defparam \A_mul_result[21] .is_wysiwyg = "true";
defparam \A_mul_result[21] .power_up = "low";

cyclonev_lcell_comb \Add26~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[22]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[22]~q ),
	.datag(gnd),
	.cin(\Add26~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~101_sumout ),
	.cout(\Add26~102 ),
	.shareout());
defparam \Add26~101 .extended_lut = "off";
defparam \Add26~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~101 .shared_arith = "off";

dffeas \A_mul_result[22] (
	.clk(clk_clk),
	.d(\Add26~101_sumout ),
	.asdata(\A_mul_partial_prod[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[22]~q ),
	.prn(vcc));
defparam \A_mul_result[22] .is_wysiwyg = "true";
defparam \A_mul_result[22] .power_up = "low";

cyclonev_lcell_comb \Add26~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[23]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[23]~q ),
	.datag(gnd),
	.cin(\Add26~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~121_sumout ),
	.cout(\Add26~122 ),
	.shareout());
defparam \Add26~121 .extended_lut = "off";
defparam \Add26~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~121 .shared_arith = "off";

dffeas \A_mul_result[23] (
	.clk(clk_clk),
	.d(\Add26~121_sumout ),
	.asdata(\A_mul_partial_prod[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[23]~q ),
	.prn(vcc));
defparam \A_mul_result[23] .is_wysiwyg = "true";
defparam \A_mul_result[23] .power_up = "low";

cyclonev_lcell_comb \Add26~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[24]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[24]~q ),
	.datag(gnd),
	.cin(\Add26~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~117_sumout ),
	.cout(\Add26~118 ),
	.shareout());
defparam \Add26~117 .extended_lut = "off";
defparam \Add26~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~117 .shared_arith = "off";

dffeas \A_mul_result[24] (
	.clk(clk_clk),
	.d(\Add26~117_sumout ),
	.asdata(\A_mul_partial_prod[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[24]~q ),
	.prn(vcc));
defparam \A_mul_result[24] .is_wysiwyg = "true";
defparam \A_mul_result[24] .power_up = "low";

cyclonev_lcell_comb \Add26~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[25]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[25]~q ),
	.datag(gnd),
	.cin(\Add26~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~85_sumout ),
	.cout(\Add26~86 ),
	.shareout());
defparam \Add26~85 .extended_lut = "off";
defparam \Add26~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~85 .shared_arith = "off";

dffeas \A_mul_result[25] (
	.clk(clk_clk),
	.d(\Add26~85_sumout ),
	.asdata(\A_mul_partial_prod[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[25]~q ),
	.prn(vcc));
defparam \A_mul_result[25] .is_wysiwyg = "true";
defparam \A_mul_result[25] .power_up = "low";

cyclonev_lcell_comb \Add26~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[26]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[26]~q ),
	.datag(gnd),
	.cin(\Add26~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~81_sumout ),
	.cout(\Add26~82 ),
	.shareout());
defparam \Add26~81 .extended_lut = "off";
defparam \Add26~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~81 .shared_arith = "off";

dffeas \A_mul_result[26] (
	.clk(clk_clk),
	.d(\Add26~81_sumout ),
	.asdata(\A_mul_partial_prod[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[26]~q ),
	.prn(vcc));
defparam \A_mul_result[26] .is_wysiwyg = "true";
defparam \A_mul_result[26] .power_up = "low";

cyclonev_lcell_comb \Add26~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[27]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[27]~q ),
	.datag(gnd),
	.cin(\Add26~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~73_sumout ),
	.cout(\Add26~74 ),
	.shareout());
defparam \Add26~73 .extended_lut = "off";
defparam \Add26~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~73 .shared_arith = "off";

dffeas \A_mul_result[27] (
	.clk(clk_clk),
	.d(\Add26~73_sumout ),
	.asdata(\A_mul_partial_prod[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[27]~q ),
	.prn(vcc));
defparam \A_mul_result[27] .is_wysiwyg = "true";
defparam \A_mul_result[27] .power_up = "low";

cyclonev_lcell_comb \Add26~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[28]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[28]~q ),
	.datag(gnd),
	.cin(\Add26~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~69_sumout ),
	.cout(\Add26~70 ),
	.shareout());
defparam \Add26~69 .extended_lut = "off";
defparam \Add26~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~69 .shared_arith = "off";

dffeas \A_mul_result[28] (
	.clk(clk_clk),
	.d(\Add26~69_sumout ),
	.asdata(\A_mul_partial_prod[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[28]~q ),
	.prn(vcc));
defparam \A_mul_result[28] .is_wysiwyg = "true";
defparam \A_mul_result[28] .power_up = "low";

cyclonev_lcell_comb \Add26~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[29]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[29]~q ),
	.datag(gnd),
	.cin(\Add26~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~65_sumout ),
	.cout(\Add26~66 ),
	.shareout());
defparam \Add26~65 .extended_lut = "off";
defparam \Add26~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~65 .shared_arith = "off";

dffeas \A_mul_result[29] (
	.clk(clk_clk),
	.d(\Add26~65_sumout ),
	.asdata(\A_mul_partial_prod[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[29]~q ),
	.prn(vcc));
defparam \A_mul_result[29] .is_wysiwyg = "true";
defparam \A_mul_result[29] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_ld_signed~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_ld_signed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_ld_signed~0 .extended_lut = "off";
defparam \E_ctrl_ld_signed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_ld_signed~0 .shared_arith = "off";

dffeas M_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\E_ctrl_ld_signed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_signed~q ),
	.prn(vcc));
defparam M_ctrl_ld_signed.is_wysiwyg = "true";
defparam M_ctrl_ld_signed.power_up = "low";

dffeas A_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\M_ctrl_ld_signed~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_signed~q ),
	.prn(vcc));
defparam A_ctrl_ld_signed.is_wysiwyg = "true";
defparam A_ctrl_ld_signed.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_iw[13]~q ),
	.dataf(!\Equal169~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~0 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_ctrl_shift_right_arith~0 .shared_arith = "off";

dffeas E_ctrl_shift_right_arith(
	.clk(clk_clk),
	.d(\D_ctrl_shift_right_arith~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_right_arith~q ),
	.prn(vcc));
defparam E_ctrl_shift_right_arith.is_wysiwyg = "true";
defparam E_ctrl_shift_right_arith.power_up = "low";

cyclonev_lcell_comb \E_rot_fill_bit~0 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_ctrl_shift_right_arith~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_fill_bit~0 .extended_lut = "off";
defparam \E_rot_fill_bit~0 .lut_mask = 64'h7777777777777777;
defparam \E_rot_fill_bit~0 .shared_arith = "off";

dffeas M_rot_fill_bit(
	.clk(clk_clk),
	.d(\E_rot_fill_bit~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_fill_bit~q ),
	.prn(vcc));
defparam M_rot_fill_bit.is_wysiwyg = "true";
defparam M_rot_fill_bit.power_up = "low";

cyclonev_lcell_comb \F_iw[8]~24 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[8]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[8]~24 .extended_lut = "off";
defparam \F_iw[8]~24 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[8]~24 .shared_arith = "off";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

dffeas \d_readdata_d1[2] (
	.clk(clk_clk),
	.d(d_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[2]~q ),
	.prn(vcc));
defparam \d_readdata_d1[2] .is_wysiwyg = "true";
defparam \d_readdata_d1[2] .power_up = "low";

dffeas \d_readdata_d1[18] (
	.clk(clk_clk),
	.d(d_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[18]~q ),
	.prn(vcc));
defparam \d_readdata_d1[18] .is_wysiwyg = "true";
defparam \d_readdata_d1[18] .power_up = "low";

dffeas \d_readdata_d1[10] (
	.clk(clk_clk),
	.d(d_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[10]~q ),
	.prn(vcc));
defparam \d_readdata_d1[10] .is_wysiwyg = "true";
defparam \d_readdata_d1[10] .power_up = "low";

dffeas \d_readdata_d1[26] (
	.clk(clk_clk),
	.d(d_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[26]~q ),
	.prn(vcc));
defparam \d_readdata_d1[26] .is_wysiwyg = "true";
defparam \d_readdata_d1[26] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[2]~2 (
	.dataa(!\d_readdata_d1[2]~q ),
	.datab(!\d_readdata_d1[18]~q ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[2]~2 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[2]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal152~6 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal152~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal152~6 .extended_lut = "off";
defparam \Equal152~6 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \Equal152~6 .shared_arith = "off";

cyclonev_lcell_comb E_ctrl_div_signed_nxt(
	.dataa(!\Equal169~0_combout ),
	.datab(!\Equal152~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_div_signed_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_ctrl_div_signed_nxt.extended_lut = "off";
defparam E_ctrl_div_signed_nxt.lut_mask = 64'h7777777777777777;
defparam E_ctrl_div_signed_nxt.shared_arith = "off";

dffeas E_ctrl_div_signed(
	.clk(clk_clk),
	.d(\E_ctrl_div_signed_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_div_signed~q ),
	.prn(vcc));
defparam E_ctrl_div_signed.is_wysiwyg = "true";
defparam E_ctrl_div_signed.power_up = "low";

cyclonev_lcell_comb \E_div_negate_src2~0 (
	.dataa(!\E_src2[31]~q ),
	.datab(!\E_ctrl_div_signed~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_div_negate_src2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_div_negate_src2~0 .extended_lut = "off";
defparam \E_div_negate_src2~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \E_div_negate_src2~0 .shared_arith = "off";

cyclonev_lcell_comb \E_div_negate_src1~0 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_ctrl_div_signed~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_div_negate_src1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_div_negate_src1~0 .extended_lut = "off";
defparam \E_div_negate_src1~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \E_div_negate_src1~0 .shared_arith = "off";

cyclonev_lcell_comb E_div_negate_result(
	.dataa(!\E_div_negate_src2~0_combout ),
	.datab(!\E_div_negate_src1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_div_negate_result~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_div_negate_result.extended_lut = "off";
defparam E_div_negate_result.lut_mask = 64'h6666666666666666;
defparam E_div_negate_result.shared_arith = "off";

dffeas M_div_negate_result(
	.clk(clk_clk),
	.d(\E_div_negate_result~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_div_negate_result~q ),
	.prn(vcc));
defparam M_div_negate_result.is_wysiwyg = "true";
defparam M_div_negate_result.power_up = "low";

dffeas A_div_negate_result(
	.clk(clk_clk),
	.d(\M_div_negate_result~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_div_negate_result~q ),
	.prn(vcc));
defparam A_div_negate_result.is_wysiwyg = "true";
defparam A_div_negate_result.power_up = "low";

cyclonev_lcell_comb \A_div_quot_bit~0 (
	.dataa(!\Add11~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_quot_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_quot_bit~0 .extended_lut = "off";
defparam \A_div_quot_bit~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \A_div_quot_bit~0 .shared_arith = "off";

dffeas A_div_quot_bit(
	.clk(clk_clk),
	.d(\A_div_quot_bit~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_quot_bit~q ),
	.prn(vcc));
defparam A_div_quot_bit.is_wysiwyg = "true";
defparam A_div_quot_bit.power_up = "low";

cyclonev_lcell_comb \Add14~5 (
	.dataa(!\A_div_negate_result~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_last_quotient_bit~q ),
	.datae(gnd),
	.dataf(!\A_div_quot_bit~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~5_sumout ),
	.cout(\Add14~6 ),
	.shareout());
defparam \Add14~5 .extended_lut = "off";
defparam \Add14~5 .lut_mask = 64'h000055AA000055FF;
defparam \Add14~5 .shared_arith = "off";

cyclonev_lcell_comb A_div_quot_en(
	.dataa(!\A_stall~combout ),
	.datab(!\A_div_accumulate_quotient_bits~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_quot_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_div_quot_en.extended_lut = "off";
defparam A_div_quot_en.lut_mask = 64'h7777777777777777;
defparam A_div_quot_en.shared_arith = "off";

dffeas \A_div_quot[0] (
	.clk(clk_clk),
	.d(\Add14~5_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[0]~q ),
	.prn(vcc));
defparam \A_div_quot[0] .is_wysiwyg = "true";
defparam \A_div_quot[0] .power_up = "low";

cyclonev_lcell_comb \Add14~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~93_sumout ),
	.cout(\Add14~94 ),
	.shareout());
defparam \Add14~93 .extended_lut = "off";
defparam \Add14~93 .lut_mask = 64'h00000000000000FF;
defparam \Add14~93 .shared_arith = "off";

dffeas \A_div_quot[1] (
	.clk(clk_clk),
	.d(\Add14~93_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[1]~q ),
	.prn(vcc));
defparam \A_div_quot[1] .is_wysiwyg = "true";
defparam \A_div_quot[1] .power_up = "low";

cyclonev_lcell_comb \Add14~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~9_sumout ),
	.cout(\Add14~10 ),
	.shareout());
defparam \Add14~9 .extended_lut = "off";
defparam \Add14~9 .lut_mask = 64'h00000000000000FF;
defparam \Add14~9 .shared_arith = "off";

dffeas \A_div_quot[2] (
	.clk(clk_clk),
	.d(\Add14~9_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[2]~q ),
	.prn(vcc));
defparam \A_div_quot[2] .is_wysiwyg = "true";
defparam \A_div_quot[2] .power_up = "low";

dffeas d_readdatavalid_d1(
	.clk(clk_clk),
	.d(d_readdatavalid),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdatavalid_d1~q ),
	.prn(vcc));
defparam d_readdatavalid_d1.is_wysiwyg = "true";
defparam d_readdatavalid_d1.power_up = "low";

cyclonev_lcell_comb \E_ld_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add24~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_bus~0 .extended_lut = "off";
defparam \E_ld_bus~0 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \E_ld_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_bypass(
	.clk(clk_clk),
	.d(\E_ld_bus~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_bypass.power_up = "low";

dffeas A_ctrl_ld_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_ld_bypass~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_bypass~q ),
	.prn(vcc));
defparam A_ctrl_ld_bypass.is_wysiwyg = "true";
defparam A_ctrl_ld_bypass.power_up = "low";

cyclonev_lcell_comb \F_iw[10]~13 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[10]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[10]~13 .extended_lut = "off";
defparam \F_iw[10]~13 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[10]~13 .shared_arith = "off";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

dffeas \d_readdata_d1[4] (
	.clk(clk_clk),
	.d(d_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[4]~q ),
	.prn(vcc));
defparam \d_readdata_d1[4] .is_wysiwyg = "true";
defparam \d_readdata_d1[4] .power_up = "low";

dffeas \d_readdata_d1[20] (
	.clk(clk_clk),
	.d(d_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[20]~q ),
	.prn(vcc));
defparam \d_readdata_d1[20] .is_wysiwyg = "true";
defparam \d_readdata_d1[20] .power_up = "low";

dffeas \d_readdata_d1[12] (
	.clk(clk_clk),
	.d(d_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[12]~q ),
	.prn(vcc));
defparam \d_readdata_d1[12] .is_wysiwyg = "true";
defparam \d_readdata_d1[12] .power_up = "low";

dffeas \d_readdata_d1[28] (
	.clk(clk_clk),
	.d(d_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[28]~q ),
	.prn(vcc));
defparam \d_readdata_d1[28] .is_wysiwyg = "true";
defparam \d_readdata_d1[28] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[4]~0 (
	.dataa(!\d_readdata_d1[4]~q ),
	.datab(!\d_readdata_d1[20]~q ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[4]~0 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[4]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add14~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~61_sumout ),
	.cout(\Add14~62 ),
	.shareout());
defparam \Add14~61 .extended_lut = "off";
defparam \Add14~61 .lut_mask = 64'h00000000000000FF;
defparam \Add14~61 .shared_arith = "off";

dffeas \A_div_quot[3] (
	.clk(clk_clk),
	.d(\Add14~61_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[3]~q ),
	.prn(vcc));
defparam \A_div_quot[3] .is_wysiwyg = "true";
defparam \A_div_quot[3] .power_up = "low";

cyclonev_lcell_comb \Add14~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~1_sumout ),
	.cout(\Add14~2 ),
	.shareout());
defparam \Add14~1 .extended_lut = "off";
defparam \Add14~1 .lut_mask = 64'h00000000000000FF;
defparam \Add14~1 .shared_arith = "off";

dffeas \A_div_quot[4] (
	.clk(clk_clk),
	.d(\Add14~1_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[4]~q ),
	.prn(vcc));
defparam \A_div_quot[4] .is_wysiwyg = "true";
defparam \A_div_quot[4] .power_up = "low";

dffeas \A_slow_inst_result[4] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[4]~0_combout ),
	.asdata(\A_div_quot[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[4]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[4] .is_wysiwyg = "true";
defparam \A_slow_inst_result[4] .power_up = "low";

dffeas \A_inst_result[4] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\M_alu_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[4]~q ),
	.prn(vcc));
defparam \A_inst_result[4] .is_wysiwyg = "true";
defparam \A_inst_result[4] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_hi_imm16~0 (
	.dataa(!\F_iw[5]~1_combout ),
	.datab(!\F_iw[2]~5_combout ),
	.datac(!\F_iw[0]~9_combout ),
	.datad(!\F_iw[1]~3_combout ),
	.datae(!\F_iw[4]~4_combout ),
	.dataf(!\F_iw[3]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \F_ctrl_hi_imm16~0 .lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam \F_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas D_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_hi_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam D_ctrl_hi_imm16.is_wysiwyg = "true";
defparam D_ctrl_hi_imm16.power_up = "low";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~1 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datae(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~1 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~1 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \F_ctrl_unsigned_lo_imm16~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[11]~12_combout ),
	.datad(!\F_iw[13]~8_combout ),
	.datae(!\F_op_slli~0_combout ),
	.dataf(!\F_ctrl_unsigned_lo_imm16~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~0 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~0 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \F_ctrl_unsigned_lo_imm16~0 .shared_arith = "off";

dffeas D_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam D_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam D_ctrl_unsigned_lo_imm16.power_up = "low";

cyclonev_lcell_comb \Equal300~0 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal300~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal300~0 .extended_lut = "off";
defparam \Equal300~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal300~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal169~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_shift_rot_right~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \E_rot_mask[4]~0 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[4]~0 .extended_lut = "off";
defparam \E_rot_mask[4]~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[4]~0 .shared_arith = "off";

dffeas \M_rot_mask[4] (
	.clk(clk_clk),
	.d(\E_rot_mask[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[4]~q ),
	.prn(vcc));
defparam \M_rot_mask[4] .is_wysiwyg = "true";
defparam \M_rot_mask[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[9]~31 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[9]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[9]~31 .extended_lut = "off";
defparam \F_iw[9]~31 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[9]~31 .shared_arith = "off";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

dffeas \d_readdata_d1[3] (
	.clk(clk_clk),
	.d(d_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[3]~q ),
	.prn(vcc));
defparam \d_readdata_d1[3] .is_wysiwyg = "true";
defparam \d_readdata_d1[3] .power_up = "low";

dffeas \d_readdata_d1[19] (
	.clk(clk_clk),
	.d(d_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[19]~q ),
	.prn(vcc));
defparam \d_readdata_d1[19] .is_wysiwyg = "true";
defparam \d_readdata_d1[19] .power_up = "low";

dffeas \d_readdata_d1[11] (
	.clk(clk_clk),
	.d(d_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[11]~q ),
	.prn(vcc));
defparam \d_readdata_d1[11] .is_wysiwyg = "true";
defparam \d_readdata_d1[11] .power_up = "low";

dffeas \d_readdata_d1[27] (
	.clk(clk_clk),
	.d(d_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[27]~q ),
	.prn(vcc));
defparam \d_readdata_d1[27] .is_wysiwyg = "true";
defparam \d_readdata_d1[27] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[3]~15 (
	.dataa(!\d_readdata_d1[3]~q ),
	.datab(!\d_readdata_d1[19]~q ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[3]~15 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[3]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[3]~15 .shared_arith = "off";

dffeas \A_slow_inst_result[3] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[3]~15_combout ),
	.asdata(\A_div_quot[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[3]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[3] .is_wysiwyg = "true";
defparam \A_slow_inst_result[3] .power_up = "low";

dffeas \A_inst_result[3] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\M_alu_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[3]~q ),
	.prn(vcc));
defparam \A_inst_result[3] .is_wysiwyg = "true";
defparam \A_inst_result[3] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[3]~4 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[3]~4 .extended_lut = "off";
defparam \E_rot_mask[3]~4 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[3]~4 .shared_arith = "off";

dffeas \M_rot_mask[3] (
	.clk(clk_clk),
	.d(\E_rot_mask[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[3]~q ),
	.prn(vcc));
defparam \M_rot_mask[3] .is_wysiwyg = "true";
defparam \M_rot_mask[3] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_left~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal169~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_left~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_left~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_left~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \D_ctrl_shift_rot_left~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot_left(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_left~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot_left~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_left.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_left.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill2~0 .extended_lut = "off";
defparam \E_rot_sel_fill2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill2~0 .shared_arith = "off";

dffeas M_rot_sel_fill2(
	.clk(clk_clk),
	.d(\E_rot_sel_fill2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill2~q ),
	.prn(vcc));
defparam M_rot_sel_fill2.is_wysiwyg = "true";
defparam M_rot_sel_fill2.power_up = "low";

cyclonev_lcell_comb \F_ctrl_a_not_src~0 (
	.dataa(!\F_iw[5]~1_combout ),
	.datab(!\F_iw[3]~2_combout ),
	.datac(!\F_iw[1]~3_combout ),
	.datad(!\F_iw[4]~4_combout ),
	.datae(!\F_iw[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_a_not_src~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_a_not_src~0 .extended_lut = "off";
defparam \F_ctrl_a_not_src~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_a_not_src~0 .shared_arith = "off";

dffeas D_ctrl_a_not_src(
	.clk(clk_clk),
	.d(\F_ctrl_a_not_src~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_a_not_src~q ),
	.prn(vcc));
defparam D_ctrl_a_not_src.is_wysiwyg = "true";
defparam D_ctrl_a_not_src.power_up = "low";

cyclonev_lcell_comb \E_regnum_a_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\E_dst_regnum[0]~q ),
	.datad(!\E_dst_regnum[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_a_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datac(!\E_dst_regnum[3]~q ),
	.datad(!\E_dst_regnum[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_a_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\E_dst_regnum[2]~q ),
	.datac(!\E_wr_dst_reg~0_combout ),
	.datad(!\E_regnum_a_cmp_F~0_combout ),
	.datae(!\E_regnum_a_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_a_cmp_F.extended_lut = "off";
defparam E_regnum_a_cmp_F.lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam E_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_a_cmp_F~0 (
	.dataa(!\D_wr_dst_reg~combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datac(!\D_dst_regnum[0]~1_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datae(!\D_dst_regnum[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_a_cmp_F~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \D_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \D_regnum_a_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\D_dst_regnum[4]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \D_regnum_a_cmp_F~1 .lut_mask = 64'h6666666666666666;
defparam \D_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_a_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datad(!\D_dst_regnum[3]~3_combout ),
	.datae(!\D_regnum_a_cmp_F~0_combout ),
	.dataf(!\D_regnum_a_cmp_F~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_a_cmp_F.extended_lut = "off";
defparam D_regnum_a_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_a_cmp_F.shared_arith = "off";

dffeas E_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_a_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_stall~combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_a_cmp_D.is_wysiwyg = "true";
defparam E_regnum_a_cmp_D.power_up = "low";

dffeas M_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_a_cmp_F~combout ),
	.asdata(\E_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\M_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_a_cmp_D.is_wysiwyg = "true";
defparam M_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \A_regnum_a_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\A_wr_dst_reg_from_M~q ),
	.datad(!\A_dst_regnum_from_M[0]~q ),
	.datae(!\A_dst_regnum_from_M[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \A_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \A_regnum_a_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(!\A_dst_regnum_from_M[2]~q ),
	.datad(!\A_dst_regnum_from_M[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_a_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\A_dst_regnum_from_M[4]~q ),
	.datac(!\A_regnum_a_cmp_F~0_combout ),
	.datad(!\A_regnum_a_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_a_cmp_F.extended_lut = "off";
defparam A_regnum_a_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam A_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\M_wr_dst_reg_from_E~q ),
	.datad(!\M_dst_regnum[0]~q ),
	.datae(!\M_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \M_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(!\M_dst_regnum[2]~q ),
	.datad(!\M_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_a_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\M_regnum_a_cmp_F~0_combout ),
	.datad(!\M_regnum_a_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_a_cmp_F.extended_lut = "off";
defparam M_regnum_a_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam M_regnum_a_cmp_F.shared_arith = "off";

dffeas A_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_a_cmp_F~combout ),
	.asdata(\M_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\A_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_a_cmp_D.is_wysiwyg = "true";
defparam A_regnum_a_cmp_D.power_up = "low";

dffeas W_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_a_cmp_F~combout ),
	.asdata(\A_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(vcc),
	.q(\W_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_a_cmp_D.is_wysiwyg = "true";
defparam W_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \E_src1[3]~0 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\W_regnum_a_cmp_D~q ),
	.datad(!\A_regnum_a_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[3]~0 .extended_lut = "off";
defparam \E_src1[3]~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_src1[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[3]~1 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\A_regnum_a_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[3]~1 .extended_lut = "off";
defparam \E_src1[3]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_src1[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_reg[15]~11 (
	.dataa(!\M_alu_result[15]~q ),
	.datab(!\A_wr_data_unfiltered[15]~30_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\W_wr_data[15]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[15]~11 .extended_lut = "off";
defparam \D_src1_reg[15]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[31]~19 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[31]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[31]~19 .extended_lut = "off";
defparam \F_iw[31]~19 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[31]~19 .shared_arith = "off";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cyclonev_lcell_comb \F_iw[30]~20 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[30]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[30]~20 .extended_lut = "off";
defparam \F_iw[30]~20 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[30]~20 .shared_arith = "off";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cyclonev_lcell_comb \F_iw[29]~21 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[29]~21 .extended_lut = "off";
defparam \F_iw[29]~21 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[29]~21 .shared_arith = "off";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cyclonev_lcell_comb \F_iw[27]~22 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[27]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[27]~22 .extended_lut = "off";
defparam \F_iw[27]~22 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[27]~22 .shared_arith = "off";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cyclonev_lcell_comb \F_iw[28]~23 (
	.dataa(!\norm_intr_req~0_combout ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[28]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[28]~23 .extended_lut = "off";
defparam \F_iw[28]~23 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[28]~23 .shared_arith = "off";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cyclonev_lcell_comb \Equal298~0 (
	.dataa(!\D_iw[31]~q ),
	.datab(!\D_iw[30]~q ),
	.datac(!\D_iw[29]~q ),
	.datad(!\D_iw[27]~q ),
	.datae(!\D_iw[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal298~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal298~0 .extended_lut = "off";
defparam \Equal298~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal298~0 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_E(
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\E_regnum_a_cmp_D~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_E.extended_lut = "off";
defparam D_src1_hazard_E.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam D_src1_hazard_E.shared_arith = "off";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\D_src1_reg[15]~11_combout ),
	.asdata(\E_alu_result[15]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_rot~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal169~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_rot~0 .extended_lut = "off";
defparam \D_ctrl_rot~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \D_ctrl_rot~0 .shared_arith = "off";

dffeas E_ctrl_rot(
	.clk(clk_clk),
	.d(\D_ctrl_rot~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_rot~q ),
	.prn(vcc));
defparam E_ctrl_rot.is_wysiwyg = "true";
defparam E_ctrl_rot.power_up = "low";

cyclonev_lcell_comb \E_rot_pass1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass1~0 .extended_lut = "off";
defparam \E_rot_pass1~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass1~0 .shared_arith = "off";

dffeas M_rot_pass1(
	.clk(clk_clk),
	.d(\E_rot_pass1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass1~q ),
	.prn(vcc));
defparam M_rot_pass1.is_wysiwyg = "true";
defparam M_rot_pass1.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill1~0 .extended_lut = "off";
defparam \E_rot_sel_fill1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill1~0 .shared_arith = "off";

dffeas M_rot_sel_fill1(
	.clk(clk_clk),
	.d(\E_rot_sel_fill1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill1~q ),
	.prn(vcc));
defparam M_rot_sel_fill1.is_wysiwyg = "true";
defparam M_rot_sel_fill1.power_up = "low";

cyclonev_lcell_comb \E_rot_mask[6]~7 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[6]~7 .extended_lut = "off";
defparam \E_rot_mask[6]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[6]~7 .shared_arith = "off";

dffeas \M_rot_mask[6] (
	.clk(clk_clk),
	.d(\E_rot_mask[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[6]~q ),
	.prn(vcc));
defparam \M_rot_mask[6] .is_wysiwyg = "true";
defparam \M_rot_mask[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[2]~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[2]~2 .extended_lut = "off";
defparam \E_rot_mask[2]~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[2]~2 .shared_arith = "off";

dffeas \M_rot_mask[2] (
	.clk(clk_clk),
	.d(\E_rot_mask[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[2]~q ),
	.prn(vcc));
defparam \M_rot_mask[2] .is_wysiwyg = "true";
defparam \M_rot_mask[2] .power_up = "low";

dffeas \d_readdata_d1[6] (
	.clk(clk_clk),
	.d(d_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[6]~q ),
	.prn(vcc));
defparam \d_readdata_d1[6] .is_wysiwyg = "true";
defparam \d_readdata_d1[6] .power_up = "low";

dffeas \d_readdata_d1[22] (
	.clk(clk_clk),
	.d(d_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[22]~q ),
	.prn(vcc));
defparam \d_readdata_d1[22] .is_wysiwyg = "true";
defparam \d_readdata_d1[22] .power_up = "low";

dffeas \d_readdata_d1[14] (
	.clk(clk_clk),
	.d(d_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[14]~q ),
	.prn(vcc));
defparam \d_readdata_d1[14] .is_wysiwyg = "true";
defparam \d_readdata_d1[14] .power_up = "low";

dffeas \d_readdata_d1[30] (
	.clk(clk_clk),
	.d(d_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[30]~q ),
	.prn(vcc));
defparam \d_readdata_d1[30] .is_wysiwyg = "true";
defparam \d_readdata_d1[30] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[6]~10 (
	.dataa(!\d_readdata_d1[6]~q ),
	.datab(!\d_readdata_d1[22]~q ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\d_readdata_d1[30]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[6]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[6]~10 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[6]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[6]~10 .shared_arith = "off";

cyclonev_lcell_comb \Add14~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~13_sumout ),
	.cout(\Add14~14 ),
	.shareout());
defparam \Add14~13 .extended_lut = "off";
defparam \Add14~13 .lut_mask = 64'h00000000000000FF;
defparam \Add14~13 .shared_arith = "off";

dffeas \A_div_quot[5] (
	.clk(clk_clk),
	.d(\Add14~13_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[5]~q ),
	.prn(vcc));
defparam \A_div_quot[5] .is_wysiwyg = "true";
defparam \A_div_quot[5] .power_up = "low";

cyclonev_lcell_comb \Add14~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~41_sumout ),
	.cout(\Add14~42 ),
	.shareout());
defparam \Add14~41 .extended_lut = "off";
defparam \Add14~41 .lut_mask = 64'h00000000000000FF;
defparam \Add14~41 .shared_arith = "off";

dffeas \A_div_quot[6] (
	.clk(clk_clk),
	.d(\Add14~41_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[6]~q ),
	.prn(vcc));
defparam \A_div_quot[6] .is_wysiwyg = "true";
defparam \A_div_quot[6] .power_up = "low";

dffeas \A_slow_inst_result[6] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[6]~10_combout ),
	.asdata(\A_div_quot[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[6]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[6] .is_wysiwyg = "true";
defparam \A_slow_inst_result[6] .power_up = "low";

dffeas \A_inst_result[6] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\M_alu_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[6]~q ),
	.prn(vcc));
defparam \A_inst_result[6] .is_wysiwyg = "true";
defparam \A_inst_result[6] .power_up = "low";

dffeas \A_inst_result[18] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(\M_alu_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[18]~q ),
	.prn(vcc));
defparam \A_inst_result[18] .is_wysiwyg = "true";
defparam \A_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[1]~5 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[1]~5 .extended_lut = "off";
defparam \E_rot_mask[1]~5 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[1]~5 .shared_arith = "off";

dffeas \M_rot_mask[1] (
	.clk(clk_clk),
	.d(\E_rot_mask[1]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[1]~q ),
	.prn(vcc));
defparam \M_rot_mask[1] .is_wysiwyg = "true";
defparam \M_rot_mask[1] .power_up = "low";

dffeas \d_readdata_d1[5] (
	.clk(clk_clk),
	.d(d_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[5]~q ),
	.prn(vcc));
defparam \d_readdata_d1[5] .is_wysiwyg = "true";
defparam \d_readdata_d1[5] .power_up = "low";

dffeas \d_readdata_d1[21] (
	.clk(clk_clk),
	.d(d_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[21]~q ),
	.prn(vcc));
defparam \d_readdata_d1[21] .is_wysiwyg = "true";
defparam \d_readdata_d1[21] .power_up = "low";

dffeas \d_readdata_d1[13] (
	.clk(clk_clk),
	.d(d_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[13]~q ),
	.prn(vcc));
defparam \d_readdata_d1[13] .is_wysiwyg = "true";
defparam \d_readdata_d1[13] .power_up = "low";

dffeas \d_readdata_d1[29] (
	.clk(clk_clk),
	.d(d_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[29]~q ),
	.prn(vcc));
defparam \d_readdata_d1[29] .is_wysiwyg = "true";
defparam \d_readdata_d1[29] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[5]~3 (
	.dataa(!\d_readdata_d1[5]~q ),
	.datab(!\d_readdata_d1[21]~q ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[5]~3 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[5]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[5]~3 .shared_arith = "off";

dffeas \A_slow_inst_result[5] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[5]~3_combout ),
	.asdata(\A_div_quot[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[5]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[5] .is_wysiwyg = "true";
defparam \A_slow_inst_result[5] .power_up = "low";

dffeas \A_inst_result[5] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\M_alu_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[5]~q ),
	.prn(vcc));
defparam \A_inst_result[5] .is_wysiwyg = "true";
defparam \A_inst_result[5] .power_up = "low";

dffeas \A_inst_result[17] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(\M_alu_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[17]~q ),
	.prn(vcc));
defparam \A_inst_result[17] .is_wysiwyg = "true";
defparam \A_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[0]~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[0]~1 .extended_lut = "off";
defparam \E_rot_mask[0]~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[0]~1 .shared_arith = "off";

dffeas \M_rot_mask[0] (
	.clk(clk_clk),
	.d(\E_rot_mask[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[0]~q ),
	.prn(vcc));
defparam \M_rot_mask[0] .is_wysiwyg = "true";
defparam \M_rot_mask[0] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[4]~0 (
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\A_wr_data_unfiltered[4]~3_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[4]~0 .extended_lut = "off";
defparam \D_src1_reg[4]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[4]~0 .shared_arith = "off";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\D_src1_reg[4]~0_combout ),
	.asdata(\E_alu_result[4]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[1]~23 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\A_wr_data_unfiltered[1]~52_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\W_wr_data[1]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[1]~23 .extended_lut = "off";
defparam \D_src1_reg[1]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[1]~23 .shared_arith = "off";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\D_src1_reg[1]~23_combout ),
	.asdata(\E_alu_result[1]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src2[0]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h9696969696969696;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[4]~1 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_src1[2]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[4]~1 .extended_lut = "off";
defparam \E_rot_step1[4]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h6996699669966996;
defparam \Add7~1 .shared_arith = "off";

dffeas \M_rot_prestep2[8] (
	.clk(clk_clk),
	.d(\E_rot_step1[4]~1_combout ),
	.asdata(\E_rot_step1[8]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[8]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[8] .is_wysiwyg = "true";
defparam \M_rot_prestep2[8] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[20]~27 (
	.dataa(!\M_alu_result[20]~q ),
	.datab(!\A_wr_data_unfiltered[20]~60_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[20]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[20]~27 .extended_lut = "off";
defparam \D_src1_reg[20]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[20]~27 .shared_arith = "off";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\D_src1_reg[20]~27_combout ),
	.asdata(\E_alu_result[20]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[19]~22 (
	.dataa(!\M_alu_result[19]~q ),
	.datab(!\A_wr_data_unfiltered[19]~50_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[19]~22 .extended_lut = "off";
defparam \D_src1_reg[19]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[19]~22 .shared_arith = "off";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\D_src1_reg[19]~22_combout ),
	.asdata(\E_alu_result[19]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[16]~10 (
	.dataa(!\M_alu_result[16]~q ),
	.datab(!\A_wr_data_unfiltered[16]~28_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datad(!\W_wr_data[16]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[16]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[16]~10 .extended_lut = "off";
defparam \D_src1_reg[16]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[16]~10 .shared_arith = "off";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\D_src1_reg[16]~10_combout ),
	.asdata(\E_alu_result[16]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \d_readdata_d1[7] (
	.clk(clk_clk),
	.d(d_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[7]~q ),
	.prn(vcc));
defparam \d_readdata_d1[7] .is_wysiwyg = "true";
defparam \d_readdata_d1[7] .power_up = "low";

dffeas \d_readdata_d1[23] (
	.clk(clk_clk),
	.d(d_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[23]~q ),
	.prn(vcc));
defparam \d_readdata_d1[23] .is_wysiwyg = "true";
defparam \d_readdata_d1[23] .power_up = "low";

dffeas \d_readdata_d1[15] (
	.clk(clk_clk),
	.d(d_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[15]~q ),
	.prn(vcc));
defparam \d_readdata_d1[15] .is_wysiwyg = "true";
defparam \d_readdata_d1[15] .power_up = "low";

dffeas \d_readdata_d1[31] (
	.clk(clk_clk),
	.d(d_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[31]~q ),
	.prn(vcc));
defparam \d_readdata_d1[31] .is_wysiwyg = "true";
defparam \d_readdata_d1[31] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[7]~9 (
	.dataa(!\d_readdata_d1[7]~q ),
	.datab(!\d_readdata_d1[23]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[7]~9 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[7]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \Add14~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~37_sumout ),
	.cout(\Add14~38 ),
	.shareout());
defparam \Add14~37 .extended_lut = "off";
defparam \Add14~37 .lut_mask = 64'h00000000000000FF;
defparam \Add14~37 .shared_arith = "off";

dffeas \A_div_quot[7] (
	.clk(clk_clk),
	.d(\Add14~37_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[7]~q ),
	.prn(vcc));
defparam \A_div_quot[7] .is_wysiwyg = "true";
defparam \A_div_quot[7] .power_up = "low";

dffeas \A_slow_inst_result[7] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[7]~9_combout ),
	.asdata(\A_div_quot[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[7]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[7] .is_wysiwyg = "true";
defparam \A_slow_inst_result[7] .power_up = "low";

dffeas \A_inst_result[7] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\M_alu_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[7]~q ),
	.prn(vcc));
defparam \A_inst_result[7] .is_wysiwyg = "true";
defparam \A_inst_result[7] .power_up = "low";

dffeas \A_inst_result[23] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(\M_alu_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[23]~q ),
	.prn(vcc));
defparam \A_inst_result[23] .is_wysiwyg = "true";
defparam \A_inst_result[23] .power_up = "low";

dffeas \A_inst_result[15] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.asdata(\M_alu_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[15]~q ),
	.prn(vcc));
defparam \A_inst_result[15] .is_wysiwyg = "true";
defparam \A_inst_result[15] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[7]~22 (
	.dataa(!\A_inst_result[7]~q ),
	.datab(!\A_inst_result[23]~q ),
	.datac(!\A_inst_result[15]~q ),
	.datad(!\A_inst_result[31]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[7]~22 .extended_lut = "off";
defparam \A_wr_data_unfiltered[7]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[7]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_pass0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass0~0 .extended_lut = "off";
defparam \E_rot_pass0~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass0~0 .shared_arith = "off";

dffeas M_rot_pass0(
	.clk(clk_clk),
	.d(\E_rot_pass0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass0~q ),
	.prn(vcc));
defparam M_rot_pass0.is_wysiwyg = "true";
defparam M_rot_pass0.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_left~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill0~0 .extended_lut = "off";
defparam \E_rot_sel_fill0~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill0~0 .shared_arith = "off";

dffeas M_rot_sel_fill0(
	.clk(clk_clk),
	.d(\E_rot_sel_fill0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill0~q ),
	.prn(vcc));
defparam M_rot_sel_fill0.is_wysiwyg = "true";
defparam M_rot_sel_fill0.power_up = "low";

cyclonev_lcell_comb \E_rot_mask[7]~6 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[7]~6 .extended_lut = "off";
defparam \E_rot_mask[7]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[7]~6 .shared_arith = "off";

dffeas \M_rot_mask[7] (
	.clk(clk_clk),
	.d(\E_rot_mask[7]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[7]~q ),
	.prn(vcc));
defparam \M_rot_mask[7] .is_wysiwyg = "true";
defparam \M_rot_mask[7] .power_up = "low";

dffeas \d_readdata_d1[0] (
	.clk(clk_clk),
	.d(d_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[0]~q ),
	.prn(vcc));
defparam \d_readdata_d1[0] .is_wysiwyg = "true";
defparam \d_readdata_d1[0] .power_up = "low";

dffeas \d_readdata_d1[16] (
	.clk(clk_clk),
	.d(d_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[16]~q ),
	.prn(vcc));
defparam \d_readdata_d1[16] .is_wysiwyg = "true";
defparam \d_readdata_d1[16] .power_up = "low";

dffeas \d_readdata_d1[8] (
	.clk(clk_clk),
	.d(d_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[8]~q ),
	.prn(vcc));
defparam \d_readdata_d1[8] .is_wysiwyg = "true";
defparam \d_readdata_d1[8] .power_up = "low";

dffeas \d_readdata_d1[24] (
	.clk(clk_clk),
	.d(d_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[24]~q ),
	.prn(vcc));
defparam \d_readdata_d1[24] .is_wysiwyg = "true";
defparam \d_readdata_d1[24] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[0]~1 (
	.dataa(!\d_readdata_d1[0]~q ),
	.datab(!\d_readdata_d1[16]~q ),
	.datac(!\d_readdata_d1[8]~q ),
	.datad(!\d_readdata_d1[24]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[0]~1 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[0]~1 .shared_arith = "off";

dffeas \A_slow_inst_result[0] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[0]~1_combout ),
	.asdata(\A_div_quot[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[0]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[0] .is_wysiwyg = "true";
defparam \A_slow_inst_result[0] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[0]~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\M_alu_result[0]~q ),
	.datac(!\M_ctrl_mem~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[0]~0 .extended_lut = "off";
defparam \M_inst_result[0]~0 .lut_mask = 64'h5353535353535353;
defparam \M_inst_result[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_div_stall~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_ctrl_div~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_stall~0 .extended_lut = "off";
defparam \A_div_stall~0 .lut_mask = 64'h7777777777777777;
defparam \A_div_stall~0 .shared_arith = "off";

dffeas \E_iw[6] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[6]~q ),
	.prn(vcc));
defparam \E_iw[6] .is_wysiwyg = "true";
defparam \E_iw[6] .power_up = "low";

dffeas \M_iw[6] (
	.clk(clk_clk),
	.d(\E_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[6]~q ),
	.prn(vcc));
defparam \M_iw[6] .is_wysiwyg = "true";
defparam \M_iw[6] .power_up = "low";

dffeas \E_iw[7] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[7]~q ),
	.prn(vcc));
defparam \E_iw[7] .is_wysiwyg = "true";
defparam \E_iw[7] .power_up = "low";

dffeas \M_iw[7] (
	.clk(clk_clk),
	.d(\E_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[7]~q ),
	.prn(vcc));
defparam \M_iw[7] .is_wysiwyg = "true";
defparam \M_iw[7] .power_up = "low";

dffeas \E_iw[8] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[8]~q ),
	.prn(vcc));
defparam \E_iw[8] .is_wysiwyg = "true";
defparam \E_iw[8] .power_up = "low";

dffeas \M_iw[8] (
	.clk(clk_clk),
	.d(\E_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[8]~q ),
	.prn(vcc));
defparam \M_iw[8] .is_wysiwyg = "true";
defparam \M_iw[8] .power_up = "low";

cyclonev_lcell_comb E_op_wrctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_wrctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_wrctl.extended_lut = "off";
defparam E_op_wrctl.lut_mask = 64'h7777777777777777;
defparam E_op_wrctl.shared_arith = "off";

dffeas M_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\E_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam M_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam M_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb \A_ienable_reg_irq0_nxt~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_iw[6]~q ),
	.datac(!\M_iw[7]~q ),
	.datad(!\M_iw[8]~q ),
	.datae(!\M_ctrl_wrctl_inst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ienable_reg_irq0_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ienable_reg_irq0_nxt~0 .extended_lut = "off";
defparam \A_ienable_reg_irq0_nxt~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \A_ienable_reg_irq0_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \A_ienable_reg_irq0~0 (
	.dataa(!\A_div_done~q ),
	.datab(!\A_mem_stall~q ),
	.datac(!\A_mul_stall~q ),
	.datad(!\A_div_stall~0_combout ),
	.datae(!\A_ienable_reg_irq0_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ienable_reg_irq0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ienable_reg_irq0~0 .extended_lut = "off";
defparam \A_ienable_reg_irq0~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \A_ienable_reg_irq0~0 .shared_arith = "off";

dffeas A_ienable_reg_irq0(
	.clk(clk_clk),
	.d(\M_alu_result[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ienable_reg_irq0~0_combout ),
	.q(\A_ienable_reg_irq0~q ),
	.prn(vcc));
defparam A_ienable_reg_irq0.is_wysiwyg = "true";
defparam A_ienable_reg_irq0.power_up = "low";

cyclonev_lcell_comb \A_ipending_reg_irq0_nxt~0 (
	.dataa(!\A_ienable_reg_irq0~q ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[0]~q ),
	.datac(!av_readdata_9),
	.datad(!av_readdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ipending_reg_irq0_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ipending_reg_irq0_nxt~0 .extended_lut = "off";
defparam \A_ipending_reg_irq0_nxt~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \A_ipending_reg_irq0_nxt~0 .shared_arith = "off";

dffeas A_ipending_reg_irq0(
	.clk(clk_clk),
	.d(\A_ipending_reg_irq0_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_ipending_reg_irq0~q ),
	.prn(vcc));
defparam A_ipending_reg_irq0.is_wysiwyg = "true";
defparam A_ipending_reg_irq0.power_up = "low";

cyclonev_lcell_comb \D_ctrl_exception~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_ctrl_logic~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~0 .extended_lut = "off";
defparam \D_ctrl_exception~0 .lut_mask = 64'h9F6FFFFFFFFFFFFF;
defparam \D_ctrl_exception~0 .shared_arith = "off";

dffeas E_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_exception~q ),
	.prn(vcc));
defparam E_ctrl_exception.is_wysiwyg = "true";
defparam E_ctrl_exception.power_up = "low";

dffeas M_ctrl_exception(
	.clk(clk_clk),
	.d(\E_ctrl_exception~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_exception~q ),
	.prn(vcc));
defparam M_ctrl_exception.is_wysiwyg = "true";
defparam M_ctrl_exception.power_up = "low";

cyclonev_lcell_comb \D_ctrl_crst~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_ctrl_logic~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_crst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_crst~0 .extended_lut = "off";
defparam \D_ctrl_crst~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_crst~0 .shared_arith = "off";

dffeas E_ctrl_crst(
	.clk(clk_clk),
	.d(\D_ctrl_crst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_crst~q ),
	.prn(vcc));
defparam E_ctrl_crst.is_wysiwyg = "true";
defparam E_ctrl_crst.power_up = "low";

dffeas M_ctrl_crst(
	.clk(clk_clk),
	.d(\E_ctrl_crst~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_crst~q ),
	.prn(vcc));
defparam M_ctrl_crst.is_wysiwyg = "true";
defparam M_ctrl_crst.power_up = "low";

cyclonev_lcell_comb M_wrctl_estatus(
	.dataa(!\M_iw[6]~q ),
	.datab(!\M_iw[7]~q ),
	.datac(!\M_iw[8]~q ),
	.datad(!\M_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wrctl_estatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_wrctl_estatus.extended_lut = "off";
defparam M_wrctl_estatus.lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam M_wrctl_estatus.shared_arith = "off";

cyclonev_lcell_comb \A_estatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\A_status_reg_pie~q ),
	.datac(!\M_ctrl_exception~q ),
	.datad(!\M_ctrl_crst~q ),
	.datae(!\A_estatus_reg_pie~q ),
	.dataf(!\M_wrctl_estatus~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_estatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_estatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_estatus_reg_pie_inst_nxt~0 .lut_mask = 64'hFF7FFFFFFFF7FFFF;
defparam \A_estatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas A_estatus_reg_pie(
	.clk(clk_clk),
	.d(\A_estatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always138~0_combout ),
	.q(\A_estatus_reg_pie~q ),
	.prn(vcc));
defparam A_estatus_reg_pie.is_wysiwyg = "true";
defparam A_estatus_reg_pie.power_up = "low";

cyclonev_lcell_comb M_wrctl_bstatus(
	.dataa(!\M_iw[6]~q ),
	.datab(!\M_iw[7]~q ),
	.datac(!\M_iw[8]~q ),
	.datad(!\M_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wrctl_bstatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_wrctl_bstatus.extended_lut = "off";
defparam M_wrctl_bstatus.lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam M_wrctl_bstatus.shared_arith = "off";

cyclonev_lcell_comb \A_bstatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_ctrl_break~q ),
	.datab(!\M_alu_result[0]~q ),
	.datac(!\A_status_reg_pie~q ),
	.datad(!\A_bstatus_reg_pie~q ),
	.datae(!\M_wrctl_bstatus~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_bstatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_bstatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_bstatus_reg_pie_inst_nxt~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \A_bstatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas A_bstatus_reg_pie(
	.clk(clk_clk),
	.d(\A_bstatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always138~0_combout ),
	.q(\A_bstatus_reg_pie~q ),
	.prn(vcc));
defparam A_bstatus_reg_pie.is_wysiwyg = "true";
defparam A_bstatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~0 (
	.dataa(!\A_status_reg_pie~q ),
	.datab(!\A_estatus_reg_pie~q ),
	.datac(!\A_bstatus_reg_pie~q ),
	.datad(!\A_ienable_reg_irq0~q ),
	.datae(!\D_iw[6]~q ),
	.dataf(!\D_iw[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~0 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_control_reg_rddata_muxed[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~1 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\A_ipending_reg_irq0~q ),
	.datad(!\D_iw[7]~q ),
	.datae(!\D_control_reg_rddata_muxed[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~1 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~1 .lut_mask = 64'hDF8FFFFFDF8FFFFF;
defparam \D_control_reg_rddata_muxed[0]~1 .shared_arith = "off";

dffeas \E_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[0] .power_up = "low";

dffeas \M_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[0] .power_up = "low";

dffeas \A_inst_result[0] (
	.clk(clk_clk),
	.d(\M_inst_result[0]~0_combout ),
	.asdata(\M_control_reg_rddata[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_ctrl_rdctl_inst~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[0]~q ),
	.prn(vcc));
defparam \A_inst_result[0] .is_wysiwyg = "true";
defparam \A_inst_result[0] .power_up = "low";

dffeas \A_inst_result[8] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(\M_alu_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[8]~q ),
	.prn(vcc));
defparam \A_inst_result[8] .is_wysiwyg = "true";
defparam \A_inst_result[8] .power_up = "low";

dffeas \A_inst_result[24] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(\M_alu_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[24]~q ),
	.prn(vcc));
defparam \A_inst_result[24] .is_wysiwyg = "true";
defparam \A_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~4 (
	.dataa(!\A_inst_result[0]~q ),
	.datab(!\A_inst_result[16]~q ),
	.datac(!\A_inst_result[8]~q ),
	.datad(!\A_inst_result[24]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~4 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[20]~5 (
	.dataa(!\E_src1[20]~q ),
	.datab(!\E_src1[19]~q ),
	.datac(!\E_src1[18]~q ),
	.datad(!\E_src1[17]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[20]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[20]~5 .extended_lut = "off";
defparam \E_rot_step1[20]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[20]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[24]~2 (
	.dataa(!\E_src1[24]~q ),
	.datab(!\E_src1[23]~q ),
	.datac(!\E_src1[22]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[24]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[24]~2 .extended_lut = "off";
defparam \E_rot_step1[24]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[24]~2 .shared_arith = "off";

dffeas \M_rot_prestep2[24] (
	.clk(clk_clk),
	.d(\E_rot_step1[20]~5_combout ),
	.asdata(\E_rot_step1[24]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[24]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[24] .is_wysiwyg = "true";
defparam \M_rot_prestep2[24] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[12]~7 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_src1[10]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[12]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[12]~7 .extended_lut = "off";
defparam \E_rot_step1[12]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[12]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[16]~4 (
	.dataa(!\E_src1[16]~q ),
	.datab(!\E_src1[15]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[16]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[16]~4 .extended_lut = "off";
defparam \E_rot_step1[16]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[16]~4 .shared_arith = "off";

dffeas \M_rot_prestep2[16] (
	.clk(clk_clk),
	.d(\E_rot_step1[12]~7_combout ),
	.asdata(\E_rot_step1[16]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[16]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[16] .is_wysiwyg = "true";
defparam \M_rot_prestep2[16] .power_up = "low";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src2[3]~q ),
	.datae(!\E_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h9669699696696996;
defparam \Add7~2 .shared_arith = "off";

dffeas \M_rot_rn[3] (
	.clk(clk_clk),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_rn[3]~q ),
	.prn(vcc));
defparam \M_rot_rn[3] .is_wysiwyg = "true";
defparam \M_rot_rn[3] .power_up = "low";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src2[3]~q ),
	.datae(!\E_src2[4]~q ),
	.dataf(!\E_ctrl_shift_rot_right~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h6996966996696996;
defparam \Add7~3 .shared_arith = "off";

dffeas \M_rot_rn[4] (
	.clk(clk_clk),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_rn[4]~q ),
	.prn(vcc));
defparam \M_rot_rn[4] .is_wysiwyg = "true";
defparam \M_rot_rn[4] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~1 (
	.dataa(!\M_rot_prestep2[0]~q ),
	.datab(!\M_rot_prestep2[24]~q ),
	.datac(!\M_rot_prestep2[16]~q ),
	.datad(!\M_rot_prestep2[8]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~1 .extended_lut = "off";
defparam \M_rot[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~1 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[0]~q ),
	.datae(!\M_rot[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~1 .extended_lut = "off";
defparam \A_shift_rot_result~1 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~1 .shared_arith = "off";

dffeas \A_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[0] .is_wysiwyg = "true";
defparam \A_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~1 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_slow_inst_sel~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~1 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \A_wr_data_unfiltered[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~2 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~2 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~2 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_wr_data_unfiltered[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~5 (
	.dataa(!\A_slow_inst_result[0]~q ),
	.datab(!\A_wr_data_unfiltered[0]~4_combout ),
	.datac(!\A_mul_result[0]~q ),
	.datad(!\A_shift_rot_result[0]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~5 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[0]~5 .shared_arith = "off";

dffeas \W_wr_data[0] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[0]~q ),
	.prn(vcc));
defparam \W_wr_data[0] .is_wysiwyg = "true";
defparam \W_wr_data[0] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[0]~21 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\A_wr_data_unfiltered[0]~5_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\W_wr_data[0]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[0]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[0]~21 .extended_lut = "off";
defparam \D_src1_reg[0]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[0]~21 .shared_arith = "off";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\D_src1_reg[0]~21_combout ),
	.asdata(\E_alu_result[0]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[3]~27 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_src1[1]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[3]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[3]~27 .extended_lut = "off";
defparam \E_rot_step1[3]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[3]~27 .shared_arith = "off";

dffeas \M_rot_prestep2[7] (
	.clk(clk_clk),
	.d(\E_rot_step1[3]~27_combout ),
	.asdata(\E_rot_step1[7]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[7]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[7] .is_wysiwyg = "true";
defparam \M_rot_prestep2[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[27]~29 (
	.dataa(!\E_src1[27]~q ),
	.datab(!\E_src1[26]~q ),
	.datac(!\E_src1[25]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[27]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[27]~29 .extended_lut = "off";
defparam \E_rot_step1[27]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[27]~29 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[30]~12 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[30]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[30]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[30]~12 .extended_lut = "off";
defparam \E_logic_result[30]~12 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[30]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~20 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[30]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~20 .extended_lut = "off";
defparam \E_alu_result~20 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~20 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~38 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\Add24~77_sumout ),
	.datad(!\E_alu_result~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~38 .extended_lut = "off";
defparam \D_src2_reg[30]~38 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[30]~38 .shared_arith = "off";

dffeas \A_inst_result[30] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(\M_alu_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[30]~q ),
	.prn(vcc));
defparam \A_inst_result[30] .is_wysiwyg = "true";
defparam \A_inst_result[30] .power_up = "low";

dffeas \A_mul_partial_prod[30] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[30]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[30] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[30] .power_up = "low";

cyclonev_lcell_comb \Add26~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[30]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[30]~q ),
	.datag(gnd),
	.cin(\Add26~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~77_sumout ),
	.cout(\Add26~78 ),
	.shareout());
defparam \Add26~77 .extended_lut = "off";
defparam \Add26~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~77 .shared_arith = "off";

dffeas \A_mul_result[30] (
	.clk(clk_clk),
	.d(\Add26~77_sumout ),
	.asdata(\A_mul_partial_prod[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[30]~q ),
	.prn(vcc));
defparam \A_mul_result[30] .is_wysiwyg = "true";
defparam \A_mul_result[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass3~0 .extended_lut = "off";
defparam \E_rot_pass3~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass3~0 .shared_arith = "off";

dffeas M_rot_pass3(
	.clk(clk_clk),
	.d(\E_rot_pass3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass3~q ),
	.prn(vcc));
defparam M_rot_pass3.is_wysiwyg = "true";
defparam M_rot_pass3.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill3~0 .extended_lut = "off";
defparam \E_rot_sel_fill3~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill3~0 .shared_arith = "off";

dffeas M_rot_sel_fill3(
	.clk(clk_clk),
	.d(\E_rot_sel_fill3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill3~q ),
	.prn(vcc));
defparam M_rot_sel_fill3.is_wysiwyg = "true";
defparam M_rot_sel_fill3.power_up = "low";

cyclonev_lcell_comb \E_rot_step1[26]~11 (
	.dataa(!\E_src1[26]~q ),
	.datab(!\E_src1[25]~q ),
	.datac(!\E_src1[24]~q ),
	.datad(!\E_src1[23]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[26]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[26]~11 .extended_lut = "off";
defparam \E_rot_step1[26]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[26]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[30]~8 (
	.dataa(!\E_src1[30]~q ),
	.datab(!\E_src1[29]~q ),
	.datac(!\E_src1[28]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[30]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[30]~8 .extended_lut = "off";
defparam \E_rot_step1[30]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[30]~8 .shared_arith = "off";

dffeas \M_rot_prestep2[30] (
	.clk(clk_clk),
	.d(\E_rot_step1[26]~11_combout ),
	.asdata(\E_rot_step1[30]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[30]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[30] .is_wysiwyg = "true";
defparam \M_rot_prestep2[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[2]~9 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_src1[0]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[2]~9 .extended_lut = "off";
defparam \E_rot_step1[2]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[2]~9 .shared_arith = "off";

dffeas \M_rot_prestep2[6] (
	.clk(clk_clk),
	.d(\E_rot_step1[2]~9_combout ),
	.asdata(\E_rot_step1[6]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[6]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[6] .is_wysiwyg = "true";
defparam \M_rot_prestep2[6] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~19 (
	.dataa(!\M_rot_prestep2[30]~q ),
	.datab(!\M_rot_prestep2[22]~q ),
	.datac(!\M_rot_prestep2[14]~q ),
	.datad(!\M_rot_prestep2[6]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~19 .extended_lut = "off";
defparam \M_rot[6]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~19 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~19 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[6]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~19 .extended_lut = "off";
defparam \A_shift_rot_result~19 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~19 .shared_arith = "off";

dffeas \A_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[30] .is_wysiwyg = "true";
defparam \A_shift_rot_result[30] .power_up = "low";

dffeas M_ctrl_ld8_ld16(
	.clk(clk_clk),
	.d(\E_ctrl_ld8_ld16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld8_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld8_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld8_ld16.power_up = "low";

dffeas A_ld_align_byte2_byte3_fill(
	.clk(clk_clk),
	.d(\M_ctrl_ld8_ld16~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_byte2_byte3_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte2_byte3_fill.is_wysiwyg = "true";
defparam A_ld_align_byte2_byte3_fill.power_up = "low";

dffeas \A_mem_baddr[1] (
	.clk(clk_clk),
	.d(\M_alu_result[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[1]~q ),
	.prn(vcc));
defparam \A_mem_baddr[1] .is_wysiwyg = "true";
defparam \A_mem_baddr[1] .power_up = "low";

dffeas \A_mem_baddr[0] (
	.clk(clk_clk),
	.d(\M_alu_result[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[0]~q ),
	.prn(vcc));
defparam \A_mem_baddr[0] .is_wysiwyg = "true";
defparam \A_mem_baddr[0] .power_up = "low";

dffeas A_ctrl_ld16(
	.clk(clk_clk),
	.d(\M_ctrl_ld16~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld16~q ),
	.prn(vcc));
defparam A_ctrl_ld16.is_wysiwyg = "true";
defparam A_ctrl_ld16.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_data_sign_bit~0 (
	.dataa(!\A_mem_baddr[0]~q ),
	.datab(!\A_ctrl_ld16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_sign_bit~0 .extended_lut = "off";
defparam \A_slow_ld_data_sign_bit~0 .lut_mask = 64'h7777777777777777;
defparam \A_slow_ld_data_sign_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_ld_data_fill_bit~0 (
	.dataa(!\A_mem_baddr[1]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[23]~q ),
	.datae(!\A_slow_ld_data_sign_bit~0_combout ),
	.dataf(!\A_ctrl_ld_signed~q ),
	.datag(!\d_readdata_d1[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_fill_bit~0 .extended_lut = "on";
defparam \A_slow_ld_data_fill_bit~0 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_ld_data_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[30]~19 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\A_slow_ld_data_fill_bit~0_combout ),
	.datac(!\d_readdata_d1[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[30]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[30]~19 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[30]~19 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[30]~19 .shared_arith = "off";

cyclonev_lcell_comb \Add14~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~33_sumout ),
	.cout(\Add14~34 ),
	.shareout());
defparam \Add14~33 .extended_lut = "off";
defparam \Add14~33 .lut_mask = 64'h00000000000000FF;
defparam \Add14~33 .shared_arith = "off";

dffeas \A_div_quot[8] (
	.clk(clk_clk),
	.d(\Add14~33_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[8]~q ),
	.prn(vcc));
defparam \A_div_quot[8] .is_wysiwyg = "true";
defparam \A_div_quot[8] .power_up = "low";

cyclonev_lcell_comb \Add14~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~29_sumout ),
	.cout(\Add14~30 ),
	.shareout());
defparam \Add14~29 .extended_lut = "off";
defparam \Add14~29 .lut_mask = 64'h00000000000000FF;
defparam \Add14~29 .shared_arith = "off";

dffeas \A_div_quot[9] (
	.clk(clk_clk),
	.d(\Add14~29_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[9]~q ),
	.prn(vcc));
defparam \A_div_quot[9] .is_wysiwyg = "true";
defparam \A_div_quot[9] .power_up = "low";

cyclonev_lcell_comb \Add14~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~25_sumout ),
	.cout(\Add14~26 ),
	.shareout());
defparam \Add14~25 .extended_lut = "off";
defparam \Add14~25 .lut_mask = 64'h00000000000000FF;
defparam \Add14~25 .shared_arith = "off";

dffeas \A_div_quot[10] (
	.clk(clk_clk),
	.d(\Add14~25_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[10]~q ),
	.prn(vcc));
defparam \A_div_quot[10] .is_wysiwyg = "true";
defparam \A_div_quot[10] .power_up = "low";

cyclonev_lcell_comb \Add14~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~21_sumout ),
	.cout(\Add14~22 ),
	.shareout());
defparam \Add14~21 .extended_lut = "off";
defparam \Add14~21 .lut_mask = 64'h00000000000000FF;
defparam \Add14~21 .shared_arith = "off";

dffeas \A_div_quot[11] (
	.clk(clk_clk),
	.d(\Add14~21_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[11]~q ),
	.prn(vcc));
defparam \A_div_quot[11] .is_wysiwyg = "true";
defparam \A_div_quot[11] .power_up = "low";

cyclonev_lcell_comb \Add14~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~17_sumout ),
	.cout(\Add14~18 ),
	.shareout());
defparam \Add14~17 .extended_lut = "off";
defparam \Add14~17 .lut_mask = 64'h00000000000000FF;
defparam \Add14~17 .shared_arith = "off";

dffeas \A_div_quot[12] (
	.clk(clk_clk),
	.d(\Add14~17_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[12]~q ),
	.prn(vcc));
defparam \A_div_quot[12] .is_wysiwyg = "true";
defparam \A_div_quot[12] .power_up = "low";

cyclonev_lcell_comb \Add14~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~57_sumout ),
	.cout(\Add14~58 ),
	.shareout());
defparam \Add14~57 .extended_lut = "off";
defparam \Add14~57 .lut_mask = 64'h00000000000000FF;
defparam \Add14~57 .shared_arith = "off";

dffeas \A_div_quot[13] (
	.clk(clk_clk),
	.d(\Add14~57_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[13]~q ),
	.prn(vcc));
defparam \A_div_quot[13] .is_wysiwyg = "true";
defparam \A_div_quot[13] .power_up = "low";

cyclonev_lcell_comb \Add14~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~53_sumout ),
	.cout(\Add14~54 ),
	.shareout());
defparam \Add14~53 .extended_lut = "off";
defparam \Add14~53 .lut_mask = 64'h00000000000000FF;
defparam \Add14~53 .shared_arith = "off";

dffeas \A_div_quot[14] (
	.clk(clk_clk),
	.d(\Add14~53_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[14]~q ),
	.prn(vcc));
defparam \A_div_quot[14] .is_wysiwyg = "true";
defparam \A_div_quot[14] .power_up = "low";

cyclonev_lcell_comb \Add14~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~49_sumout ),
	.cout(\Add14~50 ),
	.shareout());
defparam \Add14~49 .extended_lut = "off";
defparam \Add14~49 .lut_mask = 64'h00000000000000FF;
defparam \Add14~49 .shared_arith = "off";

dffeas \A_div_quot[15] (
	.clk(clk_clk),
	.d(\Add14~49_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[15]~q ),
	.prn(vcc));
defparam \A_div_quot[15] .is_wysiwyg = "true";
defparam \A_div_quot[15] .power_up = "low";

cyclonev_lcell_comb \Add14~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~45_sumout ),
	.cout(\Add14~46 ),
	.shareout());
defparam \Add14~45 .extended_lut = "off";
defparam \Add14~45 .lut_mask = 64'h00000000000000FF;
defparam \Add14~45 .shared_arith = "off";

dffeas \A_div_quot[16] (
	.clk(clk_clk),
	.d(\Add14~45_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[16]~q ),
	.prn(vcc));
defparam \A_div_quot[16] .is_wysiwyg = "true";
defparam \A_div_quot[16] .power_up = "low";

cyclonev_lcell_comb \Add14~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~97_sumout ),
	.cout(\Add14~98 ),
	.shareout());
defparam \Add14~97 .extended_lut = "off";
defparam \Add14~97 .lut_mask = 64'h00000000000000FF;
defparam \Add14~97 .shared_arith = "off";

dffeas \A_div_quot[17] (
	.clk(clk_clk),
	.d(\Add14~97_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[17]~q ),
	.prn(vcc));
defparam \A_div_quot[17] .is_wysiwyg = "true";
defparam \A_div_quot[17] .power_up = "low";

cyclonev_lcell_comb \Add14~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~113_sumout ),
	.cout(\Add14~114 ),
	.shareout());
defparam \Add14~113 .extended_lut = "off";
defparam \Add14~113 .lut_mask = 64'h00000000000000FF;
defparam \Add14~113 .shared_arith = "off";

dffeas \A_div_quot[18] (
	.clk(clk_clk),
	.d(\Add14~113_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[18]~q ),
	.prn(vcc));
defparam \A_div_quot[18] .is_wysiwyg = "true";
defparam \A_div_quot[18] .power_up = "low";

cyclonev_lcell_comb \Add14~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~89_sumout ),
	.cout(\Add14~90 ),
	.shareout());
defparam \Add14~89 .extended_lut = "off";
defparam \Add14~89 .lut_mask = 64'h00000000000000FF;
defparam \Add14~89 .shared_arith = "off";

dffeas \A_div_quot[19] (
	.clk(clk_clk),
	.d(\Add14~89_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[19]~q ),
	.prn(vcc));
defparam \A_div_quot[19] .is_wysiwyg = "true";
defparam \A_div_quot[19] .power_up = "low";

cyclonev_lcell_comb \Add14~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~109_sumout ),
	.cout(\Add14~110 ),
	.shareout());
defparam \Add14~109 .extended_lut = "off";
defparam \Add14~109 .lut_mask = 64'h00000000000000FF;
defparam \Add14~109 .shared_arith = "off";

dffeas \A_div_quot[20] (
	.clk(clk_clk),
	.d(\Add14~109_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[20]~q ),
	.prn(vcc));
defparam \A_div_quot[20] .is_wysiwyg = "true";
defparam \A_div_quot[20] .power_up = "low";

cyclonev_lcell_comb \Add14~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~105_sumout ),
	.cout(\Add14~106 ),
	.shareout());
defparam \Add14~105 .extended_lut = "off";
defparam \Add14~105 .lut_mask = 64'h00000000000000FF;
defparam \Add14~105 .shared_arith = "off";

dffeas \A_div_quot[21] (
	.clk(clk_clk),
	.d(\Add14~105_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[21]~q ),
	.prn(vcc));
defparam \A_div_quot[21] .is_wysiwyg = "true";
defparam \A_div_quot[21] .power_up = "low";

cyclonev_lcell_comb \Add14~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~101_sumout ),
	.cout(\Add14~102 ),
	.shareout());
defparam \Add14~101 .extended_lut = "off";
defparam \Add14~101 .lut_mask = 64'h00000000000000FF;
defparam \Add14~101 .shared_arith = "off";

dffeas \A_div_quot[22] (
	.clk(clk_clk),
	.d(\Add14~101_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[22]~q ),
	.prn(vcc));
defparam \A_div_quot[22] .is_wysiwyg = "true";
defparam \A_div_quot[22] .power_up = "low";

cyclonev_lcell_comb \Add14~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~121_sumout ),
	.cout(\Add14~122 ),
	.shareout());
defparam \Add14~121 .extended_lut = "off";
defparam \Add14~121 .lut_mask = 64'h00000000000000FF;
defparam \Add14~121 .shared_arith = "off";

dffeas \A_div_quot[23] (
	.clk(clk_clk),
	.d(\Add14~121_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[23]~q ),
	.prn(vcc));
defparam \A_div_quot[23] .is_wysiwyg = "true";
defparam \A_div_quot[23] .power_up = "low";

cyclonev_lcell_comb \Add14~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~117_sumout ),
	.cout(\Add14~118 ),
	.shareout());
defparam \Add14~117 .extended_lut = "off";
defparam \Add14~117 .lut_mask = 64'h00000000000000FF;
defparam \Add14~117 .shared_arith = "off";

dffeas \A_div_quot[24] (
	.clk(clk_clk),
	.d(\Add14~117_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[24]~q ),
	.prn(vcc));
defparam \A_div_quot[24] .is_wysiwyg = "true";
defparam \A_div_quot[24] .power_up = "low";

cyclonev_lcell_comb \Add14~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~85_sumout ),
	.cout(\Add14~86 ),
	.shareout());
defparam \Add14~85 .extended_lut = "off";
defparam \Add14~85 .lut_mask = 64'h00000000000000FF;
defparam \Add14~85 .shared_arith = "off";

dffeas \A_div_quot[25] (
	.clk(clk_clk),
	.d(\Add14~85_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[25]~q ),
	.prn(vcc));
defparam \A_div_quot[25] .is_wysiwyg = "true";
defparam \A_div_quot[25] .power_up = "low";

cyclonev_lcell_comb \Add14~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~81_sumout ),
	.cout(\Add14~82 ),
	.shareout());
defparam \Add14~81 .extended_lut = "off";
defparam \Add14~81 .lut_mask = 64'h00000000000000FF;
defparam \Add14~81 .shared_arith = "off";

dffeas \A_div_quot[26] (
	.clk(clk_clk),
	.d(\Add14~81_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[26]~q ),
	.prn(vcc));
defparam \A_div_quot[26] .is_wysiwyg = "true";
defparam \A_div_quot[26] .power_up = "low";

cyclonev_lcell_comb \Add14~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~73_sumout ),
	.cout(\Add14~74 ),
	.shareout());
defparam \Add14~73 .extended_lut = "off";
defparam \Add14~73 .lut_mask = 64'h00000000000000FF;
defparam \Add14~73 .shared_arith = "off";

dffeas \A_div_quot[27] (
	.clk(clk_clk),
	.d(\Add14~73_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[27]~q ),
	.prn(vcc));
defparam \A_div_quot[27] .is_wysiwyg = "true";
defparam \A_div_quot[27] .power_up = "low";

cyclonev_lcell_comb \Add14~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~69_sumout ),
	.cout(\Add14~70 ),
	.shareout());
defparam \Add14~69 .extended_lut = "off";
defparam \Add14~69 .lut_mask = 64'h00000000000000FF;
defparam \Add14~69 .shared_arith = "off";

dffeas \A_div_quot[28] (
	.clk(clk_clk),
	.d(\Add14~69_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[28]~q ),
	.prn(vcc));
defparam \A_div_quot[28] .is_wysiwyg = "true";
defparam \A_div_quot[28] .power_up = "low";

cyclonev_lcell_comb \Add14~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~65_sumout ),
	.cout(\Add14~66 ),
	.shareout());
defparam \Add14~65 .extended_lut = "off";
defparam \Add14~65 .lut_mask = 64'h00000000000000FF;
defparam \Add14~65 .shared_arith = "off";

dffeas \A_div_quot[29] (
	.clk(clk_clk),
	.d(\Add14~65_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[29]~q ),
	.prn(vcc));
defparam \A_div_quot[29] .is_wysiwyg = "true";
defparam \A_div_quot[29] .power_up = "low";

cyclonev_lcell_comb \Add14~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~77_sumout ),
	.cout(\Add14~78 ),
	.shareout());
defparam \Add14~77 .extended_lut = "off";
defparam \Add14~77 .lut_mask = 64'h00000000000000FF;
defparam \Add14~77 .shared_arith = "off";

dffeas \A_div_quot[30] (
	.clk(clk_clk),
	.d(\Add14~77_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[30]~q ),
	.prn(vcc));
defparam \A_div_quot[30] .is_wysiwyg = "true";
defparam \A_div_quot[30] .power_up = "low";

dffeas \A_slow_inst_result[30] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[30]~19_combout ),
	.asdata(\A_div_quot[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[30]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[30] .is_wysiwyg = "true";
defparam \A_slow_inst_result[30] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[30]~43 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[30]~q ),
	.dataf(!\A_slow_inst_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[30]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[30]~43 .extended_lut = "off";
defparam \A_wr_data_unfiltered[30]~43 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[30]~43 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[30]~44 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[30]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[30]~q ),
	.datae(!\A_wr_data_unfiltered[30]~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[30]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[30]~44 .extended_lut = "off";
defparam \A_wr_data_unfiltered[30]~44 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[30]~44 .shared_arith = "off";

dffeas \W_wr_data[30] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[30]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[30]~q ),
	.prn(vcc));
defparam \W_wr_data[30] .is_wysiwyg = "true";
defparam \W_wr_data[30] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[30]~39 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\A_wr_data_unfiltered[30]~44_combout ),
	.dataf(!\M_alu_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~39 .extended_lut = "off";
defparam \D_src2_reg[30]~39 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[30]~39 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~8 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\Equal300~0_combout ),
	.datac(!\D_iw[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~8 .extended_lut = "off";
defparam \D_src2[30]~8 .lut_mask = 64'h4747474747474747;
defparam \D_src2[30]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~9 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[30]~38_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datae(!\D_src2_reg[30]~39_combout ),
	.dataf(!\D_src2[30]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~9 .extended_lut = "off";
defparam \D_src2[30]~9 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[30]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[18]~1 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[18]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[18]~1 .extended_lut = "off";
defparam \E_src2[18]~1 .lut_mask = 64'h7777777777777777;
defparam \E_src2[18]~1 .shared_arith = "off";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\D_src2[30]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclonev_lcell_comb \Add24~85 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~q ),
	.datag(gnd),
	.cin(\Add24~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~85_sumout ),
	.cout(\Add24~86 ),
	.shareout());
defparam \Add24~85 .extended_lut = "off";
defparam \Add24~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~85 .shared_arith = "off";

cyclonev_lcell_comb \Add24~81 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~q ),
	.datag(gnd),
	.cin(\Add24~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~81_sumout ),
	.cout(\Add24~82 ),
	.shareout());
defparam \Add24~81 .extended_lut = "off";
defparam \Add24~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~81 .shared_arith = "off";

cyclonev_lcell_comb \Add24~77 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(\Add24~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~77_sumout ),
	.cout(\Add24~78 ),
	.shareout());
defparam \Add24~77 .extended_lut = "off";
defparam \Add24~77 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~77 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~77_sumout ),
	.datac(!\E_alu_result~20_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30] .extended_lut = "off";
defparam \E_alu_result[30] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[30] .shared_arith = "off";

dffeas \M_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[30]~q ),
	.prn(vcc));
defparam \M_alu_result[30] .is_wysiwyg = "true";
defparam \M_alu_result[30] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[30]~18 (
	.dataa(!\M_alu_result[30]~q ),
	.datab(!\A_wr_data_unfiltered[30]~44_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[30]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[30]~18 .extended_lut = "off";
defparam \D_src1_reg[30]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[30]~18 .shared_arith = "off";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\D_src1_reg[30]~18_combout ),
	.asdata(\E_alu_result[30]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[31]~26 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_src1[30]~q ),
	.datac(!\E_src1[29]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[31]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[31]~26 .extended_lut = "off";
defparam \E_rot_step1[31]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[31]~26 .shared_arith = "off";

dffeas \M_rot_prestep2[31] (
	.clk(clk_clk),
	.d(\E_rot_step1[27]~29_combout ),
	.asdata(\E_rot_step1[31]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[31]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[31] .is_wysiwyg = "true";
defparam \M_rot_prestep2[31] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[19]~31 (
	.dataa(!\E_src1[19]~q ),
	.datab(!\E_src1[18]~q ),
	.datac(!\E_src1[17]~q ),
	.datad(!\E_src1[16]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[19]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[19]~31 .extended_lut = "off";
defparam \E_rot_step1[19]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[19]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[23]~28 (
	.dataa(!\E_src1[23]~q ),
	.datab(!\E_src1[22]~q ),
	.datac(!\E_src1[21]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[23]~28 .extended_lut = "off";
defparam \E_rot_step1[23]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[23]~28 .shared_arith = "off";

dffeas \M_rot_prestep2[23] (
	.clk(clk_clk),
	.d(\E_rot_step1[19]~31_combout ),
	.asdata(\E_rot_step1[23]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[23]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[23] .is_wysiwyg = "true";
defparam \M_rot_prestep2[23] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[11]~25 (
	.dataa(!\E_src1[11]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_src1[9]~q ),
	.datad(!\E_src1[8]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[11]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[11]~25 .extended_lut = "off";
defparam \E_rot_step1[11]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[11]~25 .shared_arith = "off";

dffeas \M_rot_prestep2[15] (
	.clk(clk_clk),
	.d(\E_rot_step1[11]~25_combout ),
	.asdata(\E_rot_step1[15]~30_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[15]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[15] .is_wysiwyg = "true";
defparam \M_rot_prestep2[15] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~9 (
	.dataa(!\M_rot_prestep2[7]~q ),
	.datab(!\M_rot_prestep2[31]~q ),
	.datac(!\M_rot_prestep2[23]~q ),
	.datad(!\M_rot_prestep2[15]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~9 .extended_lut = "off";
defparam \M_rot[7]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~9 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[7]~q ),
	.datae(!\M_rot[7]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~9 .extended_lut = "off";
defparam \A_shift_rot_result~9 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~9 .shared_arith = "off";

dffeas \A_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[7] .is_wysiwyg = "true";
defparam \A_shift_rot_result[7] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[7]~23 (
	.dataa(!\A_slow_inst_result[7]~q ),
	.datab(!\A_wr_data_unfiltered[7]~22_combout ),
	.datac(!\A_mul_result[7]~q ),
	.datad(!\A_shift_rot_result[7]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[7]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[7]~23 .extended_lut = "off";
defparam \A_wr_data_unfiltered[7]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[7]~23 .shared_arith = "off";

dffeas \W_wr_data[7] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[7]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[7]~q ),
	.prn(vcc));
defparam \W_wr_data[7] .is_wysiwyg = "true";
defparam \W_wr_data[7] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[7]~19 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\A_wr_data_unfiltered[7]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~19 .extended_lut = "off";
defparam \D_src2_reg[7]~19 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[7]~19 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[7]~20 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[7]~19_combout ),
	.datad(!\E_alu_result[7]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~20 .extended_lut = "off";
defparam \D_src2_reg[7]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[0]~0 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[0]~0 .extended_lut = "off";
defparam \E_src2[0]~0 .lut_mask = 64'h7777777777777777;
defparam \E_src2[0]~0 .shared_arith = "off";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(\D_src2_reg[7]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cyclonev_lcell_comb \Add24~134 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add24~134_cout ),
	.shareout());
defparam \Add24~134 .extended_lut = "off";
defparam \Add24~134 .lut_mask = 64'h0000000000005555;
defparam \Add24~134 .shared_arith = "off";

cyclonev_lcell_comb \Add24~73 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~q ),
	.datag(gnd),
	.cin(\Add24~134_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~73_sumout ),
	.cout(\Add24~74 ),
	.shareout());
defparam \Add24~73 .extended_lut = "off";
defparam \Add24~73 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~73 .shared_arith = "off";

cyclonev_lcell_comb \Add24~69 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~q ),
	.datag(gnd),
	.cin(\Add24~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~69_sumout ),
	.cout(\Add24~70 ),
	.shareout());
defparam \Add24~69 .extended_lut = "off";
defparam \Add24~69 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~69 .shared_arith = "off";

cyclonev_lcell_comb \Add24~25 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~q ),
	.datag(gnd),
	.cin(\Add24~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~25_sumout ),
	.cout(\Add24~26 ),
	.shareout());
defparam \Add24~25 .extended_lut = "off";
defparam \Add24~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~25 .shared_arith = "off";

cyclonev_lcell_comb \Add24~29 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~q ),
	.datag(gnd),
	.cin(\Add24~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~29_sumout ),
	.cout(\Add24~30 ),
	.shareout());
defparam \Add24~29 .extended_lut = "off";
defparam \Add24~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~29 .shared_arith = "off";

cyclonev_lcell_comb \Add24~33 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~q ),
	.datag(gnd),
	.cin(\Add24~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~33_sumout ),
	.cout(\Add24~34 ),
	.shareout());
defparam \Add24~33 .extended_lut = "off";
defparam \Add24~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~33 .shared_arith = "off";

cyclonev_lcell_comb \Add24~17 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(\Add24~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~17_sumout ),
	.cout(\Add24~18 ),
	.shareout());
defparam \Add24~17 .extended_lut = "off";
defparam \Add24~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~17 .shared_arith = "off";

cyclonev_lcell_comb \Add24~21 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(\Add24~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~21_sumout ),
	.cout(\Add24~22 ),
	.shareout());
defparam \Add24~21 .extended_lut = "off";
defparam \Add24~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~21 .shared_arith = "off";

cyclonev_lcell_comb \Add24~9 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~q ),
	.datag(gnd),
	.cin(\Add24~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~9_sumout ),
	.cout(\Add24~10 ),
	.shareout());
defparam \Add24~9 .extended_lut = "off";
defparam \Add24~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~9 (
	.dataa(!\E_src2[7]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~9 .extended_lut = "off";
defparam \E_alu_result~9 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~9 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_jmp_indirect_nxt~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\Equal169~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_jmp_indirect_nxt~0 .extended_lut = "off";
defparam \E_ctrl_jmp_indirect_nxt~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \E_ctrl_jmp_indirect_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid_jmp_indirect~0 (
	.dataa(!\D_valid~combout ),
	.datab(!\E_ctrl_jmp_indirect_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid_jmp_indirect~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid_jmp_indirect~0 .extended_lut = "off";
defparam \E_valid_jmp_indirect~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid_jmp_indirect~0 .shared_arith = "off";

dffeas E_valid_jmp_indirect(
	.clk(clk_clk),
	.d(\E_valid_jmp_indirect~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_valid_jmp_indirect~q ),
	.prn(vcc));
defparam E_valid_jmp_indirect.is_wysiwyg = "true";
defparam E_valid_jmp_indirect.power_up = "low";

dffeas E_ctrl_jmp_indirect(
	.clk(clk_clk),
	.d(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_jmp_indirect~q ),
	.prn(vcc));
defparam E_ctrl_jmp_indirect.is_wysiwyg = "true";
defparam E_ctrl_jmp_indirect.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[0]~0 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[0]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \M_pipe_flush_waddr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr[0]~1 (
	.dataa(!\E_ctrl_break~q ),
	.datab(!\E_ctrl_exception~q ),
	.datac(!\M_pipe_flush_waddr[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[0]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr[0]~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_pipe_flush_waddr[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[5]~5 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\E_extra_pc[5]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[5]~5 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[5]~5 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[5]~5 .shared_arith = "off";

dffeas \D_pc[5] (
	.clk(clk_clk),
	.d(\F_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[5]~q ),
	.prn(vcc));
defparam \D_pc[5] .is_wysiwyg = "true";
defparam \D_pc[5] .power_up = "low";

dffeas \E_pc[5] (
	.clk(clk_clk),
	.d(\D_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[5]~q ),
	.prn(vcc));
defparam \E_pc[5] .is_wysiwyg = "true";
defparam \E_pc[5] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[0]~2 (
	.dataa(!\E_ctrl_crst~q ),
	.datab(!\M_pipe_flush_waddr[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[0]~2 .extended_lut = "off";
defparam \M_pipe_flush_waddr[0]~2 .lut_mask = 64'h7777777777777777;
defparam \M_pipe_flush_waddr[0]~2 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[5] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[5]~5_combout ),
	.asdata(\E_pc[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[5]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[5] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[5] .power_up = "low";

dffeas \D_pc[12] (
	.clk(clk_clk),
	.d(\F_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[12]~q ),
	.prn(vcc));
defparam \D_pc[12] .is_wysiwyg = "true";
defparam \D_pc[12] .power_up = "low";

dffeas \D_pc[11] (
	.clk(clk_clk),
	.d(\F_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[11]~q ),
	.prn(vcc));
defparam \D_pc[11] .is_wysiwyg = "true";
defparam \D_pc[11] .power_up = "low";

dffeas \D_pc[10] (
	.clk(clk_clk),
	.d(\F_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[10]~q ),
	.prn(vcc));
defparam \D_pc[10] .is_wysiwyg = "true";
defparam \D_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datae(gnd),
	.dataf(!\Add3~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[0] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[0]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[0] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[0] .power_up = "low";

dffeas \D_pc_plus_one[0] (
	.clk(clk_clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[0]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[0] .is_wysiwyg = "true";
defparam \D_pc_plus_one[0] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_br_cond_nxt~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_br_cond_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_br_cond_nxt~0 .extended_lut = "off";
defparam \E_ctrl_br_cond_nxt~0 .lut_mask = 64'hAFFF3FFFFFFFFFFF;
defparam \E_ctrl_br_cond_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb D_br_pred_not_taken(
	.dataa(!\D_bht_data[1]~q ),
	.datab(!\E_ctrl_br_cond_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_not_taken~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_br_pred_not_taken.extended_lut = "off";
defparam D_br_pred_not_taken.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam D_br_pred_not_taken.shared_arith = "off";

dffeas \E_extra_pc[0] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[0]~q ),
	.asdata(\D_pc_plus_one[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[0]~q ),
	.prn(vcc));
defparam \E_extra_pc[0] .is_wysiwyg = "true";
defparam \E_extra_pc[0] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[0]~11 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_extra_pc[0]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[0]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[0]~11 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[0]~11 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[0]~11 .shared_arith = "off";

dffeas \D_pc[0] (
	.clk(clk_clk),
	.d(\F_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[0]~q ),
	.prn(vcc));
defparam \D_pc[0] .is_wysiwyg = "true";
defparam \D_pc[0] .power_up = "low";

dffeas \E_pc[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[0]~q ),
	.prn(vcc));
defparam \E_pc[0] .is_wysiwyg = "true";
defparam \E_pc[0] .power_up = "low";

dffeas \M_pipe_flush_waddr[0] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[0]~11_combout ),
	.asdata(\E_pc[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[0]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[0] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[0] .power_up = "low";

cyclonev_lcell_comb \F_ic_valid~4 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.datad(!\F_pc[0]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_pc[2]~q ),
	.datag(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~4 .extended_lut = "on";
defparam \F_ic_valid~4 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_valid~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\F_pc[2]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_ic_valid~4_combout ),
	.datag(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~0 .extended_lut = "on";
defparam \F_ic_valid~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_hit~0 (
	.dataa(!\F_pc[10]~q ),
	.datab(!\F_pc[11]~q ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~0 .extended_lut = "off";
defparam \F_ic_hit~0 .lut_mask = 64'h6996699669966996;
defparam \F_ic_hit~0 .shared_arith = "off";

dffeas \D_pc[14] (
	.clk(clk_clk),
	.d(\F_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[14]~q ),
	.prn(vcc));
defparam \D_pc[14] .is_wysiwyg = "true";
defparam \D_pc[14] .power_up = "low";

dffeas \D_pc[13] (
	.clk(clk_clk),
	.d(\F_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[13]~q ),
	.prn(vcc));
defparam \D_pc[13] .is_wysiwyg = "true";
defparam \D_pc[13] .power_up = "low";

cyclonev_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout());
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h00000000000000FF;
defparam \Add3~49 .shared_arith = "off";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h00000000000000FF;
defparam \Add3~45 .shared_arith = "off";

dffeas \D_pc_plus_one[13] (
	.clk(clk_clk),
	.d(\Add3~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[13]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[13] .is_wysiwyg = "true";
defparam \D_pc_plus_one[13] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datae(gnd),
	.dataf(!\Add3~57_sumout ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datae(gnd),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datae(gnd),
	.dataf(!\Add3~9_sumout ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datae(gnd),
	.dataf(!\Add3~37_sumout ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datae(gnd),
	.dataf(!\Add3~33_sumout ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datae(gnd),
	.dataf(!\Add3~29_sumout ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datae(gnd),
	.dataf(!\Add3~25_sumout ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datae(gnd),
	.dataf(!\Add3~21_sumout ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datae(gnd),
	.dataf(!\Add3~17_sumout ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000000000000000;
defparam \Add0~41 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[10] (
	.clk(clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[10]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[10] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[10] .power_up = "low";

cyclonev_lcell_comb \Add1~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_br_taken_waddr_partial[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~22_cout ),
	.shareout());
defparam \Add1~22 .extended_lut = "off";
defparam \Add1~22 .lut_mask = 64'h00000000000000FF;
defparam \Add1~22 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[10]~q ),
	.datae(gnd),
	.dataf(!\D_iw[18]~q ),
	.datag(gnd),
	.cin(\Add1~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[11]~q ),
	.datae(gnd),
	.dataf(!\D_iw[19]~q ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[12]~q ),
	.datae(gnd),
	.dataf(!\D_iw[20]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[13]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~8 (
	.dataa(!\D_pc[13]~q ),
	.datab(!\Add1~9_sumout ),
	.datac(!\Add3~45_sumout ),
	.datad(!\D_iw[19]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~8 .extended_lut = "off";
defparam \F_pc_nxt~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~8 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~9 (
	.dataa(!\E_src1[15]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~9 .extended_lut = "off";
defparam \F_pc_nxt~9 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~9 .shared_arith = "off";

dffeas \E_extra_pc[13] (
	.clk(clk_clk),
	.d(\Add1~9_sumout ),
	.asdata(\D_pc_plus_one[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[13]~q ),
	.prn(vcc));
defparam \E_extra_pc[13] .is_wysiwyg = "true";
defparam \E_extra_pc[13] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[13]~10 (
	.dataa(!\E_src1[15]~q ),
	.datab(!\E_extra_pc[13]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[13]~10 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[13]~10 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \M_pipe_flush_waddr_nxt[13]~10 .shared_arith = "off";

dffeas \E_pc[13] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[13]~q ),
	.prn(vcc));
defparam \E_pc[13] .is_wysiwyg = "true";
defparam \E_pc[13] .power_up = "low";

dffeas \M_pipe_flush_waddr[13] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[13]~10_combout ),
	.asdata(\E_pc[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[13]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[13] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[13] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_nxt~9_combout ),
	.asdata(\M_pipe_flush_waddr[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[13]~q ),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h00000000000000FF;
defparam \Add3~41 .shared_arith = "off";

dffeas \D_pc_plus_one[14] (
	.clk(clk_clk),
	.d(\Add3~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[14]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[14] .is_wysiwyg = "true";
defparam \D_pc_plus_one[14] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[14]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~6 (
	.dataa(!\D_pc[14]~q ),
	.datab(!\Add1~5_sumout ),
	.datac(!\Add3~41_sumout ),
	.datad(!\D_iw[20]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~6 .extended_lut = "off";
defparam \F_pc_nxt~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~7 (
	.dataa(!\E_src1[16]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~7 .extended_lut = "off";
defparam \F_pc_nxt~7 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~7 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr[12]~3 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_break~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_crst~q ),
	.datae(!\E_ctrl_jmp_indirect~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[12]~3 .extended_lut = "off";
defparam \M_pipe_flush_waddr[12]~3 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \M_pipe_flush_waddr[12]~3 .shared_arith = "off";

dffeas \E_extra_pc[14] (
	.clk(clk_clk),
	.d(\Add1~5_sumout ),
	.asdata(\D_pc_plus_one[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[14]~q ),
	.prn(vcc));
defparam \E_extra_pc[14] .is_wysiwyg = "true";
defparam \E_extra_pc[14] .power_up = "low";

dffeas \E_pc[14] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[14]~q ),
	.prn(vcc));
defparam \E_pc[14] .is_wysiwyg = "true";
defparam \E_pc[14] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[14]~14 (
	.dataa(!\E_ctrl_crst~q ),
	.datab(!\M_pipe_flush_waddr[0]~0_combout ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_src1[16]~q ),
	.datae(!\M_pipe_flush_waddr[12]~3_combout ),
	.dataf(!\E_extra_pc[14]~q ),
	.datag(!\E_pc[14]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[14]~14 .extended_lut = "on";
defparam \M_pipe_flush_waddr_nxt[14]~14 .lut_mask = 64'hFFB8BF8FFFB8BF8F;
defparam \M_pipe_flush_waddr_nxt[14]~14 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr[14]~5 (
	.dataa(!\M_pipe_flush_waddr_nxt[14]~14_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[14]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[14]~5 .extended_lut = "off";
defparam \M_pipe_flush_waddr[14]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pipe_flush_waddr[14]~5 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[14] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr[14]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[14]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[14] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[14] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[14]~_wirecell (
	.dataa(!\M_pipe_flush_waddr[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[14]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[14]~_wirecell .extended_lut = "off";
defparam \M_pipe_flush_waddr[14]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pipe_flush_waddr[14]~_wirecell .shared_arith = "off";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_nxt~7_combout ),
	.asdata(\M_pipe_flush_waddr[14]~_wirecell_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[14]~q ),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

cyclonev_lcell_comb \F_ic_hit~1 (
	.dataa(!\F_pc[14]~q ),
	.datab(!\F_pc[13]~q ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~1 .extended_lut = "off";
defparam \F_ic_hit~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_hit~1 .shared_arith = "off";

cyclonev_lcell_comb F_issue(
	.dataa(!\F_kill~1_combout ),
	.datab(!\F_pc[12]~q ),
	.datac(!\F_ic_valid~0_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datae(!\F_ic_hit~0_combout ),
	.dataf(!\F_ic_hit~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_issue~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_issue.extended_lut = "off";
defparam F_issue.lut_mask = 64'hBFEFFFFFFFFFFFFF;
defparam F_issue.shared_arith = "off";

dffeas D_issue(
	.clk(clk_clk),
	.d(\F_issue~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_issue~q ),
	.prn(vcc));
defparam D_issue.is_wysiwyg = "true";
defparam D_issue.power_up = "low";

cyclonev_lcell_comb \F_ctrl_br~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[2]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br~0 .extended_lut = "off";
defparam \F_ctrl_br~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \F_ctrl_br~0 .shared_arith = "off";

dffeas D_ctrl_br(
	.clk(clk_clk),
	.d(\F_ctrl_br~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_br~q ),
	.prn(vcc));
defparam D_ctrl_br.is_wysiwyg = "true";
defparam D_ctrl_br.power_up = "low";

cyclonev_lcell_comb \F_ctrl_br_uncond~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[5]~1_combout ),
	.datac(!\F_iw[3]~2_combout ),
	.datad(!\F_iw[1]~3_combout ),
	.datae(!\F_iw[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br_uncond~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br_uncond~0 .extended_lut = "off";
defparam \F_ctrl_br_uncond~0 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \F_ctrl_br_uncond~0 .shared_arith = "off";

dffeas D_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\F_ctrl_br_uncond~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_br_uncond~q ),
	.prn(vcc));
defparam D_ctrl_br_uncond.is_wysiwyg = "true";
defparam D_ctrl_br_uncond.power_up = "low";

cyclonev_lcell_comb \D_br_pred_taken~0 (
	.dataa(!\D_bht_data[1]~q ),
	.datab(!\D_ctrl_br~q ),
	.datac(!\D_ctrl_br_uncond~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_taken~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_br_pred_taken~0 .extended_lut = "off";
defparam \D_br_pred_taken~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_br_pred_taken~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal169~0_combout ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~2 .extended_lut = "off";
defparam \F_kill~2 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \F_kill~2 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~0 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_issue~q ),
	.datac(!\Equal103~0_combout ),
	.datad(!\D_br_pred_taken~0_combout ),
	.datae(!\F_kill~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~0 .extended_lut = "off";
defparam \F_kill~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \F_kill~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~1 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_iw_valid~q ),
	.datac(!\D_kill~q ),
	.datad(!\E_valid_jmp_indirect~q ),
	.datae(!\F_kill~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~1 .extended_lut = "off";
defparam \F_kill~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \F_kill~1 .shared_arith = "off";

dffeas D_kill(
	.clk(clk_clk),
	.d(\F_kill~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_kill~q ),
	.prn(vcc));
defparam D_kill.is_wysiwyg = "true";
defparam D_kill.power_up = "low";

cyclonev_lcell_comb \F_pc[14]~1 (
	.dataa(!\D_iw_valid~q ),
	.datab(!\D_kill~q ),
	.datac(!\D_issue~q ),
	.datad(!\D_bht_data[1]~q ),
	.datae(!\D_ctrl_br~q ),
	.dataf(!\D_ctrl_br_uncond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc[14]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc[14]~1 .extended_lut = "off";
defparam \F_pc[14]~1 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \F_pc[14]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~0 (
	.dataa(!\D_pc[0]~q ),
	.datab(!\D_br_taken_waddr_partial[0]~q ),
	.datac(!\Add3~5_sumout ),
	.datad(!\D_iw[6]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~0 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~1 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~1 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[0]~1 .shared_arith = "off";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[0]~q ),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

cyclonev_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout());
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h00000000000000FF;
defparam \Add3~57 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[1] (
	.clk(clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[1]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[1] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[1] .power_up = "low";

dffeas \D_pc_plus_one[1] (
	.clk(clk_clk),
	.d(\Add3~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[1]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[1] .is_wysiwyg = "true";
defparam \D_pc_plus_one[1] .power_up = "low";

dffeas \E_extra_pc[1] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[1]~q ),
	.asdata(\D_pc_plus_one[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[1]~q ),
	.prn(vcc));
defparam \E_extra_pc[1] .is_wysiwyg = "true";
defparam \E_extra_pc[1] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[1]~12 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\E_extra_pc[1]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[1]~12 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[1]~12 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[1]~12 .shared_arith = "off";

dffeas \D_pc[1] (
	.clk(clk_clk),
	.d(\F_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[1]~q ),
	.prn(vcc));
defparam \D_pc[1] .is_wysiwyg = "true";
defparam \D_pc[1] .power_up = "low";

dffeas \E_pc[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[1]~q ),
	.prn(vcc));
defparam \E_pc[1] .is_wysiwyg = "true";
defparam \E_pc[1] .power_up = "low";

dffeas \M_pipe_flush_waddr[1] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[1]~12_combout ),
	.asdata(\E_pc[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[1]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[1] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[1] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~2 (
	.dataa(!\D_pc[1]~q ),
	.datab(!\D_br_taken_waddr_partial[1]~q ),
	.datac(!\Add3~57_sumout ),
	.datad(!\D_iw[7]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~2 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~3 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[1]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~3 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[1]~3 .shared_arith = "off";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[1]~q ),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[2] (
	.clk(clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[2]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[2] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[2] .power_up = "low";

dffeas \D_pc_plus_one[2] (
	.clk(clk_clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[2]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[2] .is_wysiwyg = "true";
defparam \D_pc_plus_one[2] .power_up = "low";

dffeas \E_extra_pc[2] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[2]~q ),
	.asdata(\D_pc_plus_one[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[2]~q ),
	.prn(vcc));
defparam \E_extra_pc[2] .is_wysiwyg = "true";
defparam \E_extra_pc[2] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[2]~13 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_extra_pc[2]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[2]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[2]~13 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[2]~13 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[2]~13 .shared_arith = "off";

dffeas \D_pc[2] (
	.clk(clk_clk),
	.d(\F_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[2]~q ),
	.prn(vcc));
defparam \D_pc[2] .is_wysiwyg = "true";
defparam \D_pc[2] .power_up = "low";

dffeas \E_pc[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[2]~q ),
	.prn(vcc));
defparam \E_pc[2] .is_wysiwyg = "true";
defparam \E_pc[2] .power_up = "low";

dffeas \M_pipe_flush_waddr[2] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[2]~13_combout ),
	.asdata(\E_pc[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[2]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[2] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~4 (
	.dataa(!\D_pc[2]~q ),
	.datab(!\D_br_taken_waddr_partial[2]~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\D_iw[8]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~4 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~5 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[2]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~5 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[2]~5 .shared_arith = "off";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[2]~q ),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[3] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[3]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[3] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[3] .power_up = "low";

dffeas \D_pc_plus_one[3] (
	.clk(clk_clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[3]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[3] .is_wysiwyg = "true";
defparam \D_pc_plus_one[3] .power_up = "low";

dffeas \E_extra_pc[3] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[3]~q ),
	.asdata(\D_pc_plus_one[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[3]~q ),
	.prn(vcc));
defparam \E_extra_pc[3] .is_wysiwyg = "true";
defparam \E_extra_pc[3] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[3]~7 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\E_extra_pc[3]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[3]~7 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[3]~7 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \M_pipe_flush_waddr_nxt[3]~7 .shared_arith = "off";

dffeas \D_pc[3] (
	.clk(clk_clk),
	.d(\F_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[3]~q ),
	.prn(vcc));
defparam \D_pc[3] .is_wysiwyg = "true";
defparam \D_pc[3] .power_up = "low";

dffeas \E_pc[3] (
	.clk(clk_clk),
	.d(\D_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[3]~q ),
	.prn(vcc));
defparam \E_pc[3] .is_wysiwyg = "true";
defparam \E_pc[3] .power_up = "low";

dffeas \M_pipe_flush_waddr[3] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[3]~7_combout ),
	.asdata(\E_pc[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[3]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[3] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[3] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~12 (
	.dataa(!\D_pc[3]~q ),
	.datab(!\D_br_taken_waddr_partial[3]~q ),
	.datac(!\Add3~9_sumout ),
	.datad(!\D_iw[9]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~12 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[0]~12 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~13 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[3]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[0]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~13 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~13 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[0]~13 .shared_arith = "off";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[0]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[3]~q ),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h00000000000000FF;
defparam \Add3~37 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[4] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[4]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[4] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[4] .power_up = "low";

dffeas \D_pc_plus_one[4] (
	.clk(clk_clk),
	.d(\Add3~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[4]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[4] .is_wysiwyg = "true";
defparam \D_pc_plus_one[4] .power_up = "low";

dffeas \E_extra_pc[4] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[4]~q ),
	.asdata(\D_pc_plus_one[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[4]~q ),
	.prn(vcc));
defparam \E_extra_pc[4] .is_wysiwyg = "true";
defparam \E_extra_pc[4] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[4]~4 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\E_extra_pc[4]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[4]~4 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[4]~4 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[4]~4 .shared_arith = "off";

dffeas \D_pc[4] (
	.clk(clk_clk),
	.d(\F_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[4]~q ),
	.prn(vcc));
defparam \D_pc[4] .is_wysiwyg = "true";
defparam \D_pc[4] .power_up = "low";

dffeas \E_pc[4] (
	.clk(clk_clk),
	.d(\D_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[4]~q ),
	.prn(vcc));
defparam \E_pc[4] .is_wysiwyg = "true";
defparam \E_pc[4] .power_up = "low";

dffeas \M_pipe_flush_waddr[4] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[4]~4_combout ),
	.asdata(\E_pc[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[4]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[4] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[4] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~8 (
	.dataa(!\D_pc[4]~q ),
	.datab(!\D_br_taken_waddr_partial[4]~q ),
	.datac(!\Add3~37_sumout ),
	.datad(!\D_iw[10]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~8 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~9 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[4]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[1]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~9 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[1]~9 .shared_arith = "off";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[1]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[4]~q ),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h00000000000000FF;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h00000000000000FF;
defparam \Add3~29 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[6]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[6] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[6] .power_up = "low";

dffeas \D_pc_plus_one[6] (
	.clk(clk_clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[6]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[6] .is_wysiwyg = "true";
defparam \D_pc_plus_one[6] .power_up = "low";

dffeas \E_extra_pc[6] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[6]~q ),
	.asdata(\D_pc_plus_one[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[6]~q ),
	.prn(vcc));
defparam \E_extra_pc[6] .is_wysiwyg = "true";
defparam \E_extra_pc[6] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[6]~3 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\E_extra_pc[6]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[6]~3 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[6]~3 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[6]~3 .shared_arith = "off";

dffeas \D_pc[6] (
	.clk(clk_clk),
	.d(\F_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[6]~q ),
	.prn(vcc));
defparam \D_pc[6] .is_wysiwyg = "true";
defparam \D_pc[6] .power_up = "low";

dffeas \E_pc[6] (
	.clk(clk_clk),
	.d(\D_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[6]~q ),
	.prn(vcc));
defparam \E_pc[6] .is_wysiwyg = "true";
defparam \E_pc[6] .power_up = "low";

dffeas \M_pipe_flush_waddr[6] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[6]~3_combout ),
	.asdata(\E_pc[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[6]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[6] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[6] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~6 (
	.dataa(!\D_pc[6]~q ),
	.datab(!\D_br_taken_waddr_partial[6]~q ),
	.datac(!\Add3~29_sumout ),
	.datad(!\D_iw[12]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~6 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~7 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~7 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[3]~7 .shared_arith = "off";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[6]~q ),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[7] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[7]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[7] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[7] .power_up = "low";

dffeas \D_pc_plus_one[7] (
	.clk(clk_clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[7]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[7] .is_wysiwyg = "true";
defparam \D_pc_plus_one[7] .power_up = "low";

dffeas \E_extra_pc[7] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[7]~q ),
	.asdata(\D_pc_plus_one[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[7]~q ),
	.prn(vcc));
defparam \E_extra_pc[7] .is_wysiwyg = "true";
defparam \E_extra_pc[7] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[7]~1 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\E_extra_pc[7]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[7]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[7]~1 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[7]~1 .shared_arith = "off";

dffeas \D_pc[7] (
	.clk(clk_clk),
	.d(\F_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[7]~q ),
	.prn(vcc));
defparam \D_pc[7] .is_wysiwyg = "true";
defparam \D_pc[7] .power_up = "low";

dffeas \E_pc[7] (
	.clk(clk_clk),
	.d(\D_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[7]~q ),
	.prn(vcc));
defparam \E_pc[7] .is_wysiwyg = "true";
defparam \E_pc[7] .power_up = "low";

dffeas \M_pipe_flush_waddr[7] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[7]~1_combout ),
	.asdata(\E_pc[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[7]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[7] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~2 (
	.dataa(!\D_pc[7]~q ),
	.datab(!\D_br_taken_waddr_partial[7]~q ),
	.datac(!\Add3~25_sumout ),
	.datad(!\D_iw[13]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~2 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~3 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[4]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~3 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[4]~3 .shared_arith = "off";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[7]~q ),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[8] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[8]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[8] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[8] .power_up = "low";

dffeas \D_pc_plus_one[8] (
	.clk(clk_clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[8]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[8] .is_wysiwyg = "true";
defparam \D_pc_plus_one[8] .power_up = "low";

dffeas \E_extra_pc[8] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[8]~q ),
	.asdata(\D_pc_plus_one[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[8]~q ),
	.prn(vcc));
defparam \E_extra_pc[8] .is_wysiwyg = "true";
defparam \E_extra_pc[8] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[8]~2 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\E_extra_pc[8]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[8]~2 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[8]~2 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[8]~2 .shared_arith = "off";

dffeas \D_pc[8] (
	.clk(clk_clk),
	.d(\F_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[8]~q ),
	.prn(vcc));
defparam \D_pc[8] .is_wysiwyg = "true";
defparam \D_pc[8] .power_up = "low";

dffeas \E_pc[8] (
	.clk(clk_clk),
	.d(\D_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[8]~q ),
	.prn(vcc));
defparam \E_pc[8] .is_wysiwyg = "true";
defparam \E_pc[8] .power_up = "low";

dffeas \M_pipe_flush_waddr[8] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[8]~2_combout ),
	.asdata(\E_pc[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[8]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[8] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~4 (
	.dataa(!\D_pc[8]~q ),
	.datab(!\D_br_taken_waddr_partial[8]~q ),
	.datac(!\Add3~21_sumout ),
	.datad(!\D_iw[14]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~4 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~5 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[8]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[5]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~5 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[5]~5 .shared_arith = "off";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[8]~q ),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[9] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[9]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[9] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[9] .power_up = "low";

dffeas \D_pc_plus_one[9] (
	.clk(clk_clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[9]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[9] .is_wysiwyg = "true";
defparam \D_pc_plus_one[9] .power_up = "low";

dffeas \E_extra_pc[9] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[9]~q ),
	.asdata(\D_pc_plus_one[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[9]~q ),
	.prn(vcc));
defparam \E_extra_pc[9] .is_wysiwyg = "true";
defparam \E_extra_pc[9] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[9]~0 (
	.dataa(!\E_src1[11]~q ),
	.datab(!\E_extra_pc[9]~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_jmp_indirect~q ),
	.datae(!\M_pipe_flush_waddr[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[9]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[9]~0 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \M_pipe_flush_waddr_nxt[9]~0 .shared_arith = "off";

dffeas \D_pc[9] (
	.clk(clk_clk),
	.d(\F_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[9]~q ),
	.prn(vcc));
defparam \D_pc[9] .is_wysiwyg = "true";
defparam \D_pc[9] .power_up = "low";

dffeas \E_pc[9] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[9]~q ),
	.prn(vcc));
defparam \E_pc[9] .is_wysiwyg = "true";
defparam \E_pc[9] .power_up = "low";

dffeas \M_pipe_flush_waddr[9] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[9]~0_combout ),
	.asdata(\E_pc[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[9]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[9] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[9] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[6]~0 (
	.dataa(!\D_pc[9]~q ),
	.datab(!\D_br_taken_waddr_partial[9]~q ),
	.datac(!\Add3~17_sumout ),
	.datad(!\D_iw[15]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[6]~0 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[6]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[6]~1 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[9]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[6]~1 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[6]~1 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[6]~1 .shared_arith = "off";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[9]~q ),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

dffeas \D_pc_plus_one[10] (
	.clk(clk_clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[10]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[10] .is_wysiwyg = "true";
defparam \D_pc_plus_one[10] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt~2 (
	.dataa(!\D_pc[10]~q ),
	.datab(!\Add1~1_sumout ),
	.datac(!\Add3~13_sumout ),
	.datad(!\D_iw[16]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~2 .extended_lut = "off";
defparam \F_pc_nxt~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~3 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~3 .extended_lut = "off";
defparam \F_pc_nxt~3 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~3 .shared_arith = "off";

dffeas \E_extra_pc[10] (
	.clk(clk_clk),
	.d(\Add1~1_sumout ),
	.asdata(\D_pc_plus_one[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[10]~q ),
	.prn(vcc));
defparam \E_extra_pc[10] .is_wysiwyg = "true";
defparam \E_extra_pc[10] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[10]~8 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_extra_pc[10]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[10]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[10]~8 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[10]~8 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[10]~8 .shared_arith = "off";

dffeas \E_pc[10] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[10]~q ),
	.prn(vcc));
defparam \E_pc[10] .is_wysiwyg = "true";
defparam \E_pc[10] .power_up = "low";

dffeas \M_pipe_flush_waddr[10] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[10]~8_combout ),
	.asdata(\E_pc[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[10]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[10] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[10] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_nxt~3_combout ),
	.asdata(\M_pipe_flush_waddr[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[10]~q ),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout());
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h00000000000000FF;
defparam \Add3~53 .shared_arith = "off";

dffeas \D_pc_plus_one[11] (
	.clk(clk_clk),
	.d(\Add3~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[11]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[11] .is_wysiwyg = "true";
defparam \D_pc_plus_one[11] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt~4 (
	.dataa(!\D_pc[11]~q ),
	.datab(!\Add1~17_sumout ),
	.datac(!\Add3~53_sumout ),
	.datad(!\D_iw[17]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~4 .extended_lut = "off";
defparam \F_pc_nxt~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~5 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~5 .extended_lut = "off";
defparam \F_pc_nxt~5 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~5 .shared_arith = "off";

dffeas \E_extra_pc[11] (
	.clk(clk_clk),
	.d(\Add1~17_sumout ),
	.asdata(\D_pc_plus_one[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[11]~q ),
	.prn(vcc));
defparam \E_extra_pc[11] .is_wysiwyg = "true";
defparam \E_extra_pc[11] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[11]~9 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_extra_pc[11]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[11]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[11]~9 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[11]~9 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[11]~9 .shared_arith = "off";

dffeas \E_pc[11] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[11]~q ),
	.prn(vcc));
defparam \E_pc[11] .is_wysiwyg = "true";
defparam \E_pc[11] .power_up = "low";

dffeas \M_pipe_flush_waddr[11] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[11]~9_combout ),
	.asdata(\E_pc[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[11]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[11] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[11] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_nxt~5_combout ),
	.asdata(\M_pipe_flush_waddr[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[11]~q ),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \D_pc_plus_one[12] (
	.clk(clk_clk),
	.d(\Add3~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[12]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[12] .is_wysiwyg = "true";
defparam \D_pc_plus_one[12] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt~0 (
	.dataa(!\D_pc[12]~q ),
	.datab(!\Add1~13_sumout ),
	.datac(!\Add3~49_sumout ),
	.datad(!\D_iw[18]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~0 .extended_lut = "off";
defparam \F_pc_nxt~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~1 (
	.dataa(!\E_src1[14]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~1 .extended_lut = "off";
defparam \F_pc_nxt~1 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~1 .shared_arith = "off";

dffeas \E_pc[12] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[12]~q ),
	.prn(vcc));
defparam \E_pc[12] .is_wysiwyg = "true";
defparam \E_pc[12] .power_up = "low";

dffeas \E_extra_pc[12] (
	.clk(clk_clk),
	.d(\Add1~13_sumout ),
	.asdata(\D_pc_plus_one[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[12]~q ),
	.prn(vcc));
defparam \E_extra_pc[12] .is_wysiwyg = "true";
defparam \E_extra_pc[12] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[12]~6 (
	.dataa(!\E_pc[12]~q ),
	.datab(!\E_extra_pc[12]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_ctrl_crst~q ),
	.datae(!\M_pipe_flush_waddr[0]~0_combout ),
	.dataf(!\M_pipe_flush_waddr[12]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[12]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[12]~6 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[12]~6 .lut_mask = 64'hFFFEFFFFFFFFFFFE;
defparam \M_pipe_flush_waddr_nxt[12]~6 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[12] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[12]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[12]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[12] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[12] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[12]~_wirecell (
	.dataa(!\M_pipe_flush_waddr[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[12]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[12]~_wirecell .extended_lut = "off";
defparam \M_pipe_flush_waddr[12]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pipe_flush_waddr[12]~_wirecell .shared_arith = "off";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_nxt~1_combout ),
	.asdata(\M_pipe_flush_waddr[12]~_wirecell_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[12]~q ),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

cyclonev_lcell_comb \F_ic_hit~2 (
	.dataa(!\F_pc[12]~q ),
	.datab(!\F_ic_valid~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\F_ic_hit~0_combout ),
	.datae(!\F_ic_hit~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~2 .extended_lut = "off";
defparam \F_ic_hit~2 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \F_ic_hit~2 .shared_arith = "off";

dffeas D_iw_valid(
	.clk(clk_clk),
	.d(\F_ic_hit~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw_valid~q ),
	.prn(vcc));
defparam D_iw_valid.is_wysiwyg = "true";
defparam D_iw_valid.power_up = "low";

cyclonev_lcell_comb \F_pc[14]~0 (
	.dataa(!\D_iw_valid~q ),
	.datab(!\D_kill~q ),
	.datac(!\D_ctrl_a_not_src~q ),
	.datad(!\D_issue~q ),
	.datae(!\D_br_pred_taken~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc[14]~0 .extended_lut = "off";
defparam \F_pc[14]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_pc[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~10 (
	.dataa(!\D_pc[5]~q ),
	.datab(!\D_br_taken_waddr_partial[5]~q ),
	.datac(!\Add3~33_sumout ),
	.datad(!\D_iw[11]~q ),
	.datae(!\F_pc[14]~0_combout ),
	.dataf(!\F_pc[14]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~10 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~11 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[5]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[2]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~11 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[2]~11 .shared_arith = "off";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[5]~q ),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \D_br_taken_waddr_partial[5] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[5]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[5] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[5] .power_up = "low";

dffeas \D_pc_plus_one[5] (
	.clk(clk_clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[5]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[5] .is_wysiwyg = "true";
defparam \D_pc_plus_one[5] .power_up = "low";

dffeas \E_extra_pc[5] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[5]~q ),
	.asdata(\D_pc_plus_one[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[5]~q ),
	.prn(vcc));
defparam \E_extra_pc[5] .is_wysiwyg = "true";
defparam \E_extra_pc[5] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[7] (
	.dataa(!\Add24~9_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~9_combout ),
	.datae(!\E_extra_pc[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7] .extended_lut = "off";
defparam \E_alu_result[7] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[7] .shared_arith = "off";

dffeas \M_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[7]~q ),
	.prn(vcc));
defparam \M_alu_result[7] .is_wysiwyg = "true";
defparam \M_alu_result[7] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[7]~8 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\A_wr_data_unfiltered[7]~23_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[7]~8 .extended_lut = "off";
defparam \D_src1_reg[7]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[7]~8 .shared_arith = "off";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\D_src1_reg[7]~8_combout ),
	.asdata(\E_alu_result[7]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[7]~24 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src1[5]~q ),
	.datad(!\E_src1[4]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[7]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[7]~24 .extended_lut = "off";
defparam \E_rot_step1[7]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[7]~24 .shared_arith = "off";

dffeas \M_rot_prestep2[11] (
	.clk(clk_clk),
	.d(\E_rot_step1[7]~24_combout ),
	.asdata(\E_rot_step1[11]~25_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[11]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[11] .is_wysiwyg = "true";
defparam \M_rot_prestep2[11] .power_up = "low";

dffeas \M_rot_prestep2[3] (
	.clk(clk_clk),
	.d(\E_rot_step1[31]~26_combout ),
	.asdata(\E_rot_step1[3]~27_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[3]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[3] .is_wysiwyg = "true";
defparam \M_rot_prestep2[3] .power_up = "low";

dffeas \M_rot_prestep2[27] (
	.clk(clk_clk),
	.d(\E_rot_step1[23]~28_combout ),
	.asdata(\E_rot_step1[27]~29_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[27]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[27] .is_wysiwyg = "true";
defparam \M_rot_prestep2[27] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~5 (
	.dataa(!\M_rot_prestep2[11]~q ),
	.datab(!\M_rot_prestep2[3]~q ),
	.datac(!\M_rot_prestep2[27]~q ),
	.datad(!\M_rot_prestep2[19]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~5 .extended_lut = "off";
defparam \M_rot[3]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~5 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[3]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~5 .extended_lut = "off";
defparam \A_shift_rot_result~5 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~5 .shared_arith = "off";

dffeas \A_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[11] .is_wysiwyg = "true";
defparam \A_shift_rot_result[11] .power_up = "low";

dffeas \A_inst_result[11] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.asdata(\M_alu_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[11]~q ),
	.prn(vcc));
defparam \A_inst_result[11] .is_wysiwyg = "true";
defparam \A_inst_result[11] .power_up = "low";

dffeas \A_inst_result[27] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(\M_alu_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[27]~q ),
	.prn(vcc));
defparam \A_inst_result[27] .is_wysiwyg = "true";
defparam \A_inst_result[27] .power_up = "low";

dffeas A_ld_align_byte1_fill(
	.clk(clk_clk),
	.d(\M_ctrl_ld8~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_byte1_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte1_fill.is_wysiwyg = "true";
defparam A_ld_align_byte1_fill.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result[15]~0 (
	.dataa(!\A_ctrl_div~q ),
	.datab(!\A_ld_align_sh16~q ),
	.datac(!\A_ld_align_byte1_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result[15]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result[15]~0 .extended_lut = "off";
defparam \A_slow_inst_result[15]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_slow_inst_result[15]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result[15]~1 (
	.dataa(!\A_ctrl_div~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result[15]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result[15]~1 .extended_lut = "off";
defparam \A_slow_inst_result[15]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_slow_inst_result[15]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[11]~5 (
	.dataa(!\d_readdata_d1[11]~q ),
	.datab(!\d_readdata_d1[27]~q ),
	.datac(!\A_div_quot[11]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[11]~5 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[11]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[11]~5 .shared_arith = "off";

dffeas \A_slow_inst_result[11] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[11]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[11]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[11] .is_wysiwyg = "true";
defparam \A_slow_inst_result[11] .power_up = "low";

cyclonev_lcell_comb A_data_ram_ld_align_fill_bit(
	.dataa(!\A_data_ram_ld_align_sign_bit~q ),
	.datab(!\A_ctrl_ld_signed~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_data_ram_ld_align_fill_bit~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_data_ram_ld_align_fill_bit.extended_lut = "off";
defparam A_data_ram_ld_align_fill_bit.lut_mask = 64'h7777777777777777;
defparam A_data_ram_ld_align_fill_bit.shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~10 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_ld_align_byte1_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~10 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~10 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \A_wr_data_unfiltered[8]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~11 (
	.dataa(!\A_slow_inst_sel~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~11 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~11 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_wr_data_unfiltered[8]~11 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~14 (
	.dataa(!\A_inst_result[11]~q ),
	.datab(!\A_inst_result[27]~q ),
	.datac(!\A_slow_inst_result[11]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~14 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[11]~14 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~15 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[11]~q ),
	.datad(!\A_shift_rot_result[11]~q ),
	.datae(!\A_wr_data_unfiltered[11]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~15 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[11]~15 .shared_arith = "off";

dffeas \W_wr_data[11] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[11]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[11]~q ),
	.prn(vcc));
defparam \W_wr_data[11] .is_wysiwyg = "true";
defparam \W_wr_data[11] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[11]~4 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\A_wr_data_unfiltered[11]~15_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\W_wr_data[11]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[11]~4 .extended_lut = "off";
defparam \D_src1_reg[11]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[11]~4 .shared_arith = "off";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\D_src1_reg[11]~4_combout ),
	.asdata(\E_alu_result[11]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

cyclonev_lcell_comb \Add24~1 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~q ),
	.datag(gnd),
	.cin(\Add24~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~1_sumout ),
	.cout(\Add24~2 ),
	.shareout());
defparam \Add24~1 .extended_lut = "off";
defparam \Add24~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~1 .shared_arith = "off";

cyclonev_lcell_comb \Add24~5 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~q ),
	.datag(gnd),
	.cin(\Add24~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~5_sumout ),
	.cout(\Add24~6 ),
	.shareout());
defparam \Add24~5 .extended_lut = "off";
defparam \Add24~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~5 .shared_arith = "off";

cyclonev_lcell_comb \Add24~13 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(\Add24~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~13_sumout ),
	.cout(\Add24~14 ),
	.shareout());
defparam \Add24~13 .extended_lut = "off";
defparam \Add24~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~13 .shared_arith = "off";

cyclonev_lcell_comb \Add24~45 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(\Add24~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~45_sumout ),
	.cout(\Add24~46 ),
	.shareout());
defparam \Add24~45 .extended_lut = "off";
defparam \Add24~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~45 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[11]~1 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[11]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[11]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[11]~1 .extended_lut = "off";
defparam \E_logic_result[11]~1 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[11]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~5 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[11]~1_combout ),
	.datad(!\E_extra_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~5 .extended_lut = "off";
defparam \E_alu_result[11]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[11]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~45_sumout ),
	.datac(!\E_alu_result[11]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11] .extended_lut = "off";
defparam \E_alu_result[11] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[11] .shared_arith = "off";

dffeas \M_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[11]~q ),
	.prn(vcc));
defparam \M_alu_result[11] .is_wysiwyg = "true";
defparam \M_alu_result[11] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[11]~15 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[11]~q ),
	.datae(!\A_shift_rot_result[11]~q ),
	.dataf(!\A_wr_data_unfiltered[11]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~15 .extended_lut = "off";
defparam \D_src2_reg[11]~15 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[11]~15 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[11]~92 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[11]~q ),
	.dataf(!\D_src2_reg[11]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~92 .extended_lut = "off";
defparam \D_src2_reg[11]~92 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[11]~92 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[11]~123 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\D_src2_reg[11]~92_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[11]~5_combout ),
	.datag(!\Add24~45_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~123_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~123 .extended_lut = "on";
defparam \D_src2_reg[11]~123 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[11]~123 .shared_arith = "off";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(\D_src2_reg[11]~123_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cyclonev_lcell_comb \Add24~41 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(\Add24~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~41_sumout ),
	.cout(\Add24~42 ),
	.shareout());
defparam \Add24~41 .extended_lut = "off";
defparam \Add24~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~41 .shared_arith = "off";

cyclonev_lcell_comb \Add24~61 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~q ),
	.datag(gnd),
	.cin(\Add24~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~61_sumout ),
	.cout(\Add24~62 ),
	.shareout());
defparam \Add24~61 .extended_lut = "off";
defparam \Add24~61 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~61 .shared_arith = "off";

cyclonev_lcell_comb \Add24~57 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(\Add24~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~57_sumout ),
	.cout(\Add24~58 ),
	.shareout());
defparam \Add24~57 .extended_lut = "off";
defparam \Add24~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~57 .shared_arith = "off";

cyclonev_lcell_comb \Add24~53 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~q ),
	.datag(gnd),
	.cin(\Add24~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~53_sumout ),
	.cout(\Add24~54 ),
	.shareout());
defparam \Add24~53 .extended_lut = "off";
defparam \Add24~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~53 .shared_arith = "off";

cyclonev_lcell_comb \Add24~49 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(\Add24~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~49_sumout ),
	.cout(\Add24~50 ),
	.shareout());
defparam \Add24~49 .extended_lut = "off";
defparam \Add24~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~49 .shared_arith = "off";

cyclonev_lcell_comb \Add24~105 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(\Add24~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~105_sumout ),
	.cout(\Add24~106 ),
	.shareout());
defparam \Add24~105 .extended_lut = "off";
defparam \Add24~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~105 .shared_arith = "off";

cyclonev_lcell_comb \Add24~121 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(\Add24~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~121_sumout ),
	.cout(\Add24~122 ),
	.shareout());
defparam \Add24~121 .extended_lut = "off";
defparam \Add24~121 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~121 .shared_arith = "off";

cyclonev_lcell_comb \Add24~101 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(\Add24~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~101_sumout ),
	.cout(\Add24~102 ),
	.shareout());
defparam \Add24~101 .extended_lut = "off";
defparam \Add24~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~101 .shared_arith = "off";

cyclonev_lcell_comb \Add24~117 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(\Add24~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~117_sumout ),
	.cout(\Add24~118 ),
	.shareout());
defparam \Add24~117 .extended_lut = "off";
defparam \Add24~117 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~117 .shared_arith = "off";

cyclonev_lcell_comb \Add24~113 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~q ),
	.datag(gnd),
	.cin(\Add24~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~113_sumout ),
	.cout(\Add24~114 ),
	.shareout());
defparam \Add24~113 .extended_lut = "off";
defparam \Add24~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~113 .shared_arith = "off";

cyclonev_lcell_comb \Add24~109 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~q ),
	.datag(gnd),
	.cin(\Add24~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~109_sumout ),
	.cout(\Add24~110 ),
	.shareout());
defparam \Add24~109 .extended_lut = "off";
defparam \Add24~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~109 .shared_arith = "off";

cyclonev_lcell_comb \Add24~129 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(\Add24~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~129_sumout ),
	.cout(\Add24~130 ),
	.shareout());
defparam \Add24~129 .extended_lut = "off";
defparam \Add24~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~129 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~30_combout ),
	.datac(!\Add24~129_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23] .extended_lut = "off";
defparam \E_alu_result[23] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[23] .shared_arith = "off";

dffeas \M_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[23]~q ),
	.prn(vcc));
defparam \M_alu_result[23] .is_wysiwyg = "true";
defparam \M_alu_result[23] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~30 (
	.dataa(!\M_rot_prestep2[23]~q ),
	.datab(!\M_rot_prestep2[15]~q ),
	.datac(!\M_rot_prestep2[7]~q ),
	.datad(!\M_rot_prestep2[31]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~30 .extended_lut = "off";
defparam \M_rot[7]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~30 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~30 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[7]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~30 .extended_lut = "off";
defparam \A_shift_rot_result~30 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~30 .shared_arith = "off";

dffeas \A_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[23] .is_wysiwyg = "true";
defparam \A_shift_rot_result[23] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[23]~30 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[23]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[23]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[23]~30 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[23]~30 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[23]~30 .shared_arith = "off";

dffeas \A_slow_inst_result[23] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[23]~30_combout ),
	.asdata(\A_div_quot[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[23]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[23] .is_wysiwyg = "true";
defparam \A_slow_inst_result[23] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[23]~65 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[23]~q ),
	.dataf(!\A_slow_inst_result[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[23]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[23]~65 .extended_lut = "off";
defparam \A_wr_data_unfiltered[23]~65 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[23]~65 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[23]~66 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[23]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[23]~q ),
	.datae(!\A_wr_data_unfiltered[23]~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[23]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[23]~66 .extended_lut = "off";
defparam \A_wr_data_unfiltered[23]~66 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[23]~66 .shared_arith = "off";

dffeas \W_wr_data[23] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[23]~66_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[23]~q ),
	.prn(vcc));
defparam \W_wr_data[23] .is_wysiwyg = "true";
defparam \W_wr_data[23] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[23]~30 (
	.dataa(!\M_alu_result[23]~q ),
	.datab(!\A_wr_data_unfiltered[23]~66_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[23]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[23]~30 .extended_lut = "off";
defparam \D_src1_reg[23]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[23]~30 .shared_arith = "off";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\D_src1_reg[23]~30_combout ),
	.asdata(\E_alu_result[23]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~30 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[23]~q ),
	.datae(!\E_src1[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~30 .extended_lut = "off";
defparam \E_alu_result~30 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~58 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~30_combout ),
	.datad(!\Add24~129_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~58 .extended_lut = "off";
defparam \D_src2_reg[23]~58 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[23]~58 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~59 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\A_wr_data_unfiltered[23]~66_combout ),
	.dataf(!\M_alu_result[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~59 .extended_lut = "off";
defparam \D_src2_reg[23]~59 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[23]~59 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~26 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~26 .extended_lut = "off";
defparam \D_src2[23]~26 .lut_mask = 64'h5353535353535353;
defparam \D_src2[23]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~27 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[23]~58_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datae(!\D_src2_reg[23]~59_combout ),
	.dataf(!\D_src2[23]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~27 .extended_lut = "off";
defparam \D_src2[23]~27 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[23]~27 .shared_arith = "off";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\D_src2[23]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclonev_lcell_comb \Add24~125 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~q ),
	.datag(gnd),
	.cin(\Add24~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~125_sumout ),
	.cout(\Add24~126 ),
	.shareout());
defparam \Add24~125 .extended_lut = "off";
defparam \Add24~125 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~125 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~29_combout ),
	.datac(!\Add24~125_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24] .extended_lut = "off";
defparam \E_alu_result[24] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[24] .shared_arith = "off";

dffeas \M_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[24]~q ),
	.prn(vcc));
defparam \M_alu_result[24] .is_wysiwyg = "true";
defparam \M_alu_result[24] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~29 (
	.dataa(!\M_rot_prestep2[24]~q ),
	.datab(!\M_rot_prestep2[16]~q ),
	.datac(!\M_rot_prestep2[8]~q ),
	.datad(!\M_rot_prestep2[0]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~29 .extended_lut = "off";
defparam \M_rot[0]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~29 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~29 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[0]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~29 .extended_lut = "off";
defparam \A_shift_rot_result~29 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~29 .shared_arith = "off";

dffeas \A_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[24] .is_wysiwyg = "true";
defparam \A_shift_rot_result[24] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[24]~29 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[24]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[24]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[24]~29 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[24]~29 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[24]~29 .shared_arith = "off";

dffeas \A_slow_inst_result[24] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[24]~29_combout ),
	.asdata(\A_div_quot[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[24]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[24] .is_wysiwyg = "true";
defparam \A_slow_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[24]~63 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[24]~q ),
	.dataf(!\A_slow_inst_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[24]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[24]~63 .extended_lut = "off";
defparam \A_wr_data_unfiltered[24]~63 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[24]~63 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[24]~64 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[24]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[24]~q ),
	.datae(!\A_wr_data_unfiltered[24]~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[24]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[24]~64 .extended_lut = "off";
defparam \A_wr_data_unfiltered[24]~64 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[24]~64 .shared_arith = "off";

dffeas \W_wr_data[24] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[24]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[24]~q ),
	.prn(vcc));
defparam \W_wr_data[24] .is_wysiwyg = "true";
defparam \W_wr_data[24] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[24]~29 (
	.dataa(!\M_alu_result[24]~q ),
	.datab(!\A_wr_data_unfiltered[24]~64_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[24]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[24]~29 .extended_lut = "off";
defparam \D_src1_reg[24]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[24]~29 .shared_arith = "off";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\D_src1_reg[24]~29_combout ),
	.asdata(\E_alu_result[24]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~29 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[24]~q ),
	.datae(!\E_src1[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~29 .extended_lut = "off";
defparam \E_alu_result~29 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~56 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~29_combout ),
	.datad(!\Add24~125_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~56 .extended_lut = "off";
defparam \D_src2_reg[24]~56 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[24]~56 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~57 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\A_wr_data_unfiltered[24]~64_combout ),
	.dataf(!\M_alu_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~57 .extended_lut = "off";
defparam \D_src2_reg[24]~57 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[24]~57 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~24 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~24 .extended_lut = "off";
defparam \D_src2[24]~24 .lut_mask = 64'h5353535353535353;
defparam \D_src2[24]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~25 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[24]~56_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datae(!\D_src2_reg[24]~57_combout ),
	.dataf(!\D_src2[24]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~25 .extended_lut = "off";
defparam \D_src2[24]~25 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[24]~25 .shared_arith = "off";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\D_src2[24]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclonev_lcell_comb \Add24~97 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(\Add24~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~97_sumout ),
	.cout(\Add24~98 ),
	.shareout());
defparam \Add24~97 .extended_lut = "off";
defparam \Add24~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~97 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~22_combout ),
	.datac(!\Add24~97_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25] .extended_lut = "off";
defparam \E_alu_result[25] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[25] .shared_arith = "off";

dffeas \M_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[25]~q ),
	.prn(vcc));
defparam \M_alu_result[25] .is_wysiwyg = "true";
defparam \M_alu_result[25] .power_up = "low";

dffeas \A_inst_result[25] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(\M_alu_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[25]~q ),
	.prn(vcc));
defparam \A_inst_result[25] .is_wysiwyg = "true";
defparam \A_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[21]~21 (
	.dataa(!\E_src1[21]~q ),
	.datab(!\E_src1[20]~q ),
	.datac(!\E_src1[19]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[21]~21 .extended_lut = "off";
defparam \E_rot_step1[21]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[25]~18 (
	.dataa(!\E_src1[25]~q ),
	.datab(!\E_src1[24]~q ),
	.datac(!\E_src1[23]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[25]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[25]~18 .extended_lut = "off";
defparam \E_rot_step1[25]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[25]~18 .shared_arith = "off";

dffeas \M_rot_prestep2[25] (
	.clk(clk_clk),
	.d(\E_rot_step1[21]~21_combout ),
	.asdata(\E_rot_step1[25]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[25]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[25] .is_wysiwyg = "true";
defparam \M_rot_prestep2[25] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[29]~19 (
	.dataa(!\E_src1[29]~q ),
	.datab(!\E_src1[28]~q ),
	.datac(!\E_src1[27]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[29]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[29]~19 .extended_lut = "off";
defparam \E_rot_step1[29]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[29]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[1]~16 (
	.dataa(!\E_src1[1]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_src1[31]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[1]~16 .extended_lut = "off";
defparam \E_rot_step1[1]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[1]~16 .shared_arith = "off";

dffeas \M_rot_prestep2[1] (
	.clk(clk_clk),
	.d(\E_rot_step1[29]~19_combout ),
	.asdata(\E_rot_step1[1]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[1]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[1] .is_wysiwyg = "true";
defparam \M_rot_prestep2[1] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~21 (
	.dataa(!\M_rot_prestep2[25]~q ),
	.datab(!\M_rot_prestep2[17]~q ),
	.datac(!\M_rot_prestep2[9]~q ),
	.datad(!\M_rot_prestep2[1]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~21 .extended_lut = "off";
defparam \M_rot[1]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~21 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~21 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[1]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~21 .extended_lut = "off";
defparam \A_shift_rot_result~21 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~21 .shared_arith = "off";

dffeas \A_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[25] .is_wysiwyg = "true";
defparam \A_shift_rot_result[25] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[25]~21 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\A_slow_ld_data_fill_bit~0_combout ),
	.datac(!\d_readdata_d1[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[25]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[25]~21 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[25]~21 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[25]~21 .shared_arith = "off";

dffeas \A_slow_inst_result[25] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[25]~21_combout ),
	.asdata(\A_div_quot[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[25]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[25] .is_wysiwyg = "true";
defparam \A_slow_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[25]~47 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[25]~q ),
	.dataf(!\A_slow_inst_result[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[25]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[25]~47 .extended_lut = "off";
defparam \A_wr_data_unfiltered[25]~47 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[25]~47 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[25]~48 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[25]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[25]~q ),
	.datae(!\A_wr_data_unfiltered[25]~47_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[25]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[25]~48 .extended_lut = "off";
defparam \A_wr_data_unfiltered[25]~48 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[25]~48 .shared_arith = "off";

dffeas \W_wr_data[25] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[25]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[25]~q ),
	.prn(vcc));
defparam \W_wr_data[25] .is_wysiwyg = "true";
defparam \W_wr_data[25] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[25]~20 (
	.dataa(!\M_alu_result[25]~q ),
	.datab(!\A_wr_data_unfiltered[25]~48_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[25]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[25]~20 .extended_lut = "off";
defparam \D_src1_reg[25]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[25]~20 .shared_arith = "off";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\D_src1_reg[25]~20_combout ),
	.asdata(\E_alu_result[25]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~22 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[25]~q ),
	.datae(!\E_src1[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~22 .extended_lut = "off";
defparam \E_alu_result~22 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~42 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~22_combout ),
	.datad(!\Add24~97_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~42 .extended_lut = "off";
defparam \D_src2_reg[25]~42 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[25]~42 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~43 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\A_wr_data_unfiltered[25]~48_combout ),
	.dataf(!\M_alu_result[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~43 .extended_lut = "off";
defparam \D_src2_reg[25]~43 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[25]~43 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~12 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~12 .extended_lut = "off";
defparam \D_src2[25]~12 .lut_mask = 64'h5353535353535353;
defparam \D_src2[25]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~13 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[25]~42_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datae(!\D_src2_reg[25]~43_combout ),
	.dataf(!\D_src2[25]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~13 .extended_lut = "off";
defparam \D_src2[25]~13 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[25]~13 .shared_arith = "off";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\D_src2[25]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclonev_lcell_comb \Add24~93 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(\Add24~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~93_sumout ),
	.cout(\Add24~94 ),
	.shareout());
defparam \Add24~93 .extended_lut = "off";
defparam \Add24~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~93 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~21_combout ),
	.datac(!\Add24~93_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26] .extended_lut = "off";
defparam \E_alu_result[26] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[26] .shared_arith = "off";

dffeas \M_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[26]~q ),
	.prn(vcc));
defparam \M_alu_result[26] .is_wysiwyg = "true";
defparam \M_alu_result[26] .power_up = "low";

dffeas \A_inst_result[26] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(\M_alu_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[26]~q ),
	.prn(vcc));
defparam \A_inst_result[26] .is_wysiwyg = "true";
defparam \A_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[22]~10 (
	.dataa(!\E_src1[22]~q ),
	.datab(!\E_src1[21]~q ),
	.datac(!\E_src1[20]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[22]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[22]~10 .extended_lut = "off";
defparam \E_rot_step1[22]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[22]~10 .shared_arith = "off";

dffeas \M_rot_prestep2[26] (
	.clk(clk_clk),
	.d(\E_rot_step1[22]~10_combout ),
	.asdata(\E_rot_step1[26]~11_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[26]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[26] .is_wysiwyg = "true";
defparam \M_rot_prestep2[26] .power_up = "low";

dffeas \M_rot_prestep2[2] (
	.clk(clk_clk),
	.d(\E_rot_step1[30]~8_combout ),
	.asdata(\E_rot_step1[2]~9_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[2]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[2] .is_wysiwyg = "true";
defparam \M_rot_prestep2[2] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~20 (
	.dataa(!\M_rot_prestep2[26]~q ),
	.datab(!\M_rot_prestep2[18]~q ),
	.datac(!\M_rot_prestep2[10]~q ),
	.datad(!\M_rot_prestep2[2]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~20 .extended_lut = "off";
defparam \M_rot[2]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~20 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~20 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[2]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~20 .extended_lut = "off";
defparam \A_shift_rot_result~20 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~20 .shared_arith = "off";

dffeas \A_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[26] .is_wysiwyg = "true";
defparam \A_shift_rot_result[26] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[26]~20 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[26]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[26]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[26]~20 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[26]~20 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[26]~20 .shared_arith = "off";

dffeas \A_slow_inst_result[26] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[26]~20_combout ),
	.asdata(\A_div_quot[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[26]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[26] .is_wysiwyg = "true";
defparam \A_slow_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[26]~45 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[26]~q ),
	.dataf(!\A_slow_inst_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[26]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[26]~45 .extended_lut = "off";
defparam \A_wr_data_unfiltered[26]~45 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[26]~45 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[26]~46 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[26]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[26]~q ),
	.datae(!\A_wr_data_unfiltered[26]~45_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[26]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[26]~46 .extended_lut = "off";
defparam \A_wr_data_unfiltered[26]~46 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[26]~46 .shared_arith = "off";

dffeas \W_wr_data[26] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[26]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[26]~q ),
	.prn(vcc));
defparam \W_wr_data[26] .is_wysiwyg = "true";
defparam \W_wr_data[26] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[26]~19 (
	.dataa(!\M_alu_result[26]~q ),
	.datab(!\A_wr_data_unfiltered[26]~46_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[26]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[26]~19 .extended_lut = "off";
defparam \D_src1_reg[26]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[26]~19 .shared_arith = "off";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\D_src1_reg[26]~19_combout ),
	.asdata(\E_alu_result[26]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~21 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[26]~q ),
	.datae(!\E_src1[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~21 .extended_lut = "off";
defparam \E_alu_result~21 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~21 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~40 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~21_combout ),
	.datad(!\Add24~93_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~40 .extended_lut = "off";
defparam \D_src2_reg[26]~40 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[26]~40 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~41 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\A_wr_data_unfiltered[26]~46_combout ),
	.dataf(!\M_alu_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~41 .extended_lut = "off";
defparam \D_src2_reg[26]~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[26]~41 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~10 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~10 .extended_lut = "off";
defparam \D_src2[26]~10 .lut_mask = 64'h5353535353535353;
defparam \D_src2[26]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~11 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[26]~40_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datae(!\D_src2_reg[26]~41_combout ),
	.dataf(!\D_src2[26]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~11 .extended_lut = "off";
defparam \D_src2[26]~11 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[26]~11 .shared_arith = "off";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\D_src2[26]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclonev_lcell_comb \Add24~89 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~q ),
	.datag(gnd),
	.cin(\Add24~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~89_sumout ),
	.cout(\Add24~90 ),
	.shareout());
defparam \Add24~89 .extended_lut = "off";
defparam \Add24~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add24~89 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~19_combout ),
	.datac(!\Add24~89_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27] .extended_lut = "off";
defparam \E_alu_result[27] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[27] .shared_arith = "off";

dffeas \M_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[27]~q ),
	.prn(vcc));
defparam \M_alu_result[27] .is_wysiwyg = "true";
defparam \M_alu_result[27] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~18 (
	.dataa(!\M_rot_prestep2[27]~q ),
	.datab(!\M_rot_prestep2[19]~q ),
	.datac(!\M_rot_prestep2[11]~q ),
	.datad(!\M_rot_prestep2[3]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~18 .extended_lut = "off";
defparam \M_rot[3]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~18 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~18 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[3]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~18 .extended_lut = "off";
defparam \A_shift_rot_result~18 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~18 .shared_arith = "off";

dffeas \A_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[27] .is_wysiwyg = "true";
defparam \A_shift_rot_result[27] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[27]~18 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[27]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[27]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[27]~18 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[27]~18 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[27]~18 .shared_arith = "off";

dffeas \A_slow_inst_result[27] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[27]~18_combout ),
	.asdata(\A_div_quot[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[27]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[27] .is_wysiwyg = "true";
defparam \A_slow_inst_result[27] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[27]~41 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[27]~q ),
	.dataf(!\A_slow_inst_result[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[27]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[27]~41 .extended_lut = "off";
defparam \A_wr_data_unfiltered[27]~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[27]~41 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[27]~42 (
	.dataa(!\A_inst_result[27]~q ),
	.datab(!\A_ctrl_mul_lsw~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[27]~q ),
	.datae(!\A_wr_data_unfiltered[27]~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[27]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[27]~42 .extended_lut = "off";
defparam \A_wr_data_unfiltered[27]~42 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \A_wr_data_unfiltered[27]~42 .shared_arith = "off";

dffeas \W_wr_data[27] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[27]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[27]~q ),
	.prn(vcc));
defparam \W_wr_data[27] .is_wysiwyg = "true";
defparam \W_wr_data[27] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[27]~17 (
	.dataa(!\M_alu_result[27]~q ),
	.datab(!\A_wr_data_unfiltered[27]~42_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[27]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[27]~17 .extended_lut = "off";
defparam \D_src1_reg[27]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[27]~17 .shared_arith = "off";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\D_src1_reg[27]~17_combout ),
	.asdata(\E_alu_result[27]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[27]~11 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[27]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[27]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[27]~11 .extended_lut = "off";
defparam \E_logic_result[27]~11 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[27]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~19 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[27]~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~19 .extended_lut = "off";
defparam \E_alu_result~19 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~19 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~36 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~19_combout ),
	.datad(!\Add24~89_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~36 .extended_lut = "off";
defparam \D_src2_reg[27]~36 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[27]~36 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~37 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\A_wr_data_unfiltered[27]~42_combout ),
	.dataf(!\M_alu_result[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~37 .extended_lut = "off";
defparam \D_src2_reg[27]~37 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[27]~37 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~6 (
	.dataa(!\D_iw[17]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~6 .extended_lut = "off";
defparam \D_src2[27]~6 .lut_mask = 64'h5353535353535353;
defparam \D_src2[27]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~7 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[27]~36_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\D_src2_reg[27]~37_combout ),
	.dataf(!\D_src2[27]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~7 .extended_lut = "off";
defparam \D_src2[27]~7 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[27]~7 .shared_arith = "off";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\D_src2[27]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[28]~34 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~18_combout ),
	.datad(!\Add24~85_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~34 .extended_lut = "off";
defparam \D_src2_reg[28]~34 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[28]~34 .shared_arith = "off";

dffeas \A_inst_result[28] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(\M_alu_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[28]~q ),
	.prn(vcc));
defparam \A_inst_result[28] .is_wysiwyg = "true";
defparam \A_inst_result[28] .power_up = "low";

dffeas \M_rot_prestep2[28] (
	.clk(clk_clk),
	.d(\E_rot_step1[24]~2_combout ),
	.asdata(\E_rot_step1[28]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[28]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[28] .is_wysiwyg = "true";
defparam \M_rot_prestep2[28] .power_up = "low";

dffeas \M_rot_prestep2[20] (
	.clk(clk_clk),
	.d(\E_rot_step1[16]~4_combout ),
	.asdata(\E_rot_step1[20]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[20]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[20] .is_wysiwyg = "true";
defparam \M_rot_prestep2[20] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[0]~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\E_src1[31]~q ),
	.datac(!\E_src1[30]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[0]~0 .extended_lut = "off";
defparam \E_rot_step1[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[0]~0 .shared_arith = "off";

dffeas \M_rot_prestep2[4] (
	.clk(clk_clk),
	.d(\E_rot_step1[0]~0_combout ),
	.asdata(\E_rot_step1[4]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[4]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[4] .is_wysiwyg = "true";
defparam \M_rot_prestep2[4] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~17 (
	.dataa(!\M_rot_prestep2[28]~q ),
	.datab(!\M_rot_prestep2[20]~q ),
	.datac(!\M_rot_prestep2[12]~q ),
	.datad(!\M_rot_prestep2[4]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~17 .extended_lut = "off";
defparam \M_rot[4]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~17 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~17 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[4]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~17 .extended_lut = "off";
defparam \A_shift_rot_result~17 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~17 .shared_arith = "off";

dffeas \A_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[28] .is_wysiwyg = "true";
defparam \A_shift_rot_result[28] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[28]~17 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[28]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[28]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[28]~17 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[28]~17 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[28]~17 .shared_arith = "off";

dffeas \A_slow_inst_result[28] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[28]~17_combout ),
	.asdata(\A_div_quot[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[28]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[28] .is_wysiwyg = "true";
defparam \A_slow_inst_result[28] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[28]~39 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[28]~q ),
	.dataf(!\A_slow_inst_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[28]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[28]~39 .extended_lut = "off";
defparam \A_wr_data_unfiltered[28]~39 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[28]~39 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[28]~40 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[28]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[28]~q ),
	.datae(!\A_wr_data_unfiltered[28]~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[28]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[28]~40 .extended_lut = "off";
defparam \A_wr_data_unfiltered[28]~40 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[28]~40 .shared_arith = "off";

dffeas \W_wr_data[28] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[28]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[28]~q ),
	.prn(vcc));
defparam \W_wr_data[28] .is_wysiwyg = "true";
defparam \W_wr_data[28] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[28]~35 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\A_wr_data_unfiltered[28]~40_combout ),
	.dataf(!\M_alu_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~35 .extended_lut = "off";
defparam \D_src2_reg[28]~35 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[28]~35 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~4 (
	.dataa(!\D_iw[18]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~4 .extended_lut = "off";
defparam \D_src2[28]~4 .lut_mask = 64'h5353535353535353;
defparam \D_src2[28]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~5 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[28]~34_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datae(!\D_src2_reg[28]~35_combout ),
	.dataf(!\D_src2[28]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~5 .extended_lut = "off";
defparam \D_src2[28]~5 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[28]~5 .shared_arith = "off";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\D_src2[28]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[28]~10 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[28]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[28]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[28]~10 .extended_lut = "off";
defparam \E_logic_result[28]~10 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[28]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~18 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[28]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~18 .extended_lut = "off";
defparam \E_alu_result~18 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~18_combout ),
	.datac(!\Add24~85_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28] .extended_lut = "off";
defparam \E_alu_result[28] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[28] .shared_arith = "off";

dffeas \M_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[28]~q ),
	.prn(vcc));
defparam \M_alu_result[28] .is_wysiwyg = "true";
defparam \M_alu_result[28] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[28]~16 (
	.dataa(!\M_alu_result[28]~q ),
	.datab(!\A_wr_data_unfiltered[28]~40_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[28]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[28]~16 .extended_lut = "off";
defparam \D_src1_reg[28]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[28]~16 .shared_arith = "off";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\D_src1_reg[28]~16_combout ),
	.asdata(\E_alu_result[28]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[28]~3 (
	.dataa(!\E_src1[28]~q ),
	.datab(!\E_src1[27]~q ),
	.datac(!\E_src1[26]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[28]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[28]~3 .extended_lut = "off";
defparam \E_rot_step1[28]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[28]~3 .shared_arith = "off";

dffeas \M_rot_prestep2[0] (
	.clk(clk_clk),
	.d(\E_rot_step1[28]~3_combout ),
	.asdata(\E_rot_step1[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[0]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[0] .is_wysiwyg = "true";
defparam \M_rot_prestep2[0] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~8 (
	.dataa(!\M_rot_prestep2[8]~q ),
	.datab(!\M_rot_prestep2[0]~q ),
	.datac(!\M_rot_prestep2[24]~q ),
	.datad(!\M_rot_prestep2[16]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~8 .extended_lut = "off";
defparam \M_rot[0]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~8 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[0]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~8 .extended_lut = "off";
defparam \A_shift_rot_result~8 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~8 .shared_arith = "off";

dffeas \A_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[8] .is_wysiwyg = "true";
defparam \A_shift_rot_result[8] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[8]~8 (
	.dataa(!\d_readdata_d1[8]~q ),
	.datab(!\d_readdata_d1[24]~q ),
	.datac(!\A_div_quot[8]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[8]~8 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[8]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[8]~8 .shared_arith = "off";

dffeas \A_slow_inst_result[8] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[8]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[8]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[8] .is_wysiwyg = "true";
defparam \A_slow_inst_result[8] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~20 (
	.dataa(!\A_inst_result[8]~q ),
	.datab(!\A_inst_result[24]~q ),
	.datac(!\A_slow_inst_result[8]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~20 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[8]~20 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~21 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[8]~q ),
	.datad(!\A_shift_rot_result[8]~q ),
	.datae(!\A_wr_data_unfiltered[8]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~21 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[8]~21 .shared_arith = "off";

dffeas \W_wr_data[8] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[8]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[8]~q ),
	.prn(vcc));
defparam \W_wr_data[8] .is_wysiwyg = "true";
defparam \W_wr_data[8] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[8]~18 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[8]~q ),
	.datae(!\A_shift_rot_result[8]~q ),
	.dataf(!\A_wr_data_unfiltered[8]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~18 .extended_lut = "off";
defparam \D_src2_reg[8]~18 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[8]~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[8]~95 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[8]~q ),
	.dataf(!\D_src2_reg[8]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~95 .extended_lut = "off";
defparam \D_src2_reg[8]~95 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[8]~95 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[8]~4 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[8]~4 .extended_lut = "off";
defparam \E_logic_result[8]~4 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[8]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~8 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[8]~4_combout ),
	.datad(!\E_extra_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~8 .extended_lut = "off";
defparam \E_alu_result[8]~8 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[8]~111 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\D_src2_reg[8]~95_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[8]~8_combout ),
	.datag(!\Add24~1_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~111_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~111 .extended_lut = "on";
defparam \D_src2_reg[8]~111 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[8]~111 .shared_arith = "off";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(\D_src2_reg[8]~111_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[8] (
	.dataa(!\Add24~1_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[8]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8] .extended_lut = "off";
defparam \E_alu_result[8] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[8] .shared_arith = "off";

dffeas \M_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[8]~q ),
	.prn(vcc));
defparam \M_alu_result[8] .is_wysiwyg = "true";
defparam \M_alu_result[8] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[8]~7 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\A_wr_data_unfiltered[8]~21_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\W_wr_data[8]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[8]~7 .extended_lut = "off";
defparam \D_src1_reg[8]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[8]~7 .shared_arith = "off";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\D_src1_reg[8]~7_combout ),
	.asdata(\E_alu_result[8]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[8]~6 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_src1[6]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[8]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[8]~6 .extended_lut = "off";
defparam \E_rot_step1[8]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[8]~6 .shared_arith = "off";

dffeas \M_rot_prestep2[12] (
	.clk(clk_clk),
	.d(\E_rot_step1[8]~6_combout ),
	.asdata(\E_rot_step1[12]~7_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[12]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[12] .is_wysiwyg = "true";
defparam \M_rot_prestep2[12] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~4 (
	.dataa(!\M_rot_prestep2[12]~q ),
	.datab(!\M_rot_prestep2[4]~q ),
	.datac(!\M_rot_prestep2[28]~q ),
	.datad(!\M_rot_prestep2[20]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~4 .extended_lut = "off";
defparam \M_rot[4]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~4 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~4 .extended_lut = "off";
defparam \A_shift_rot_result~4 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~4 .shared_arith = "off";

dffeas \A_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[12] .is_wysiwyg = "true";
defparam \A_shift_rot_result[12] .power_up = "low";

dffeas \A_inst_result[12] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.asdata(\M_alu_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[12]~q ),
	.prn(vcc));
defparam \A_inst_result[12] .is_wysiwyg = "true";
defparam \A_inst_result[12] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[12]~4 (
	.dataa(!\d_readdata_d1[12]~q ),
	.datab(!\d_readdata_d1[28]~q ),
	.datac(!\A_div_quot[12]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[12]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[12]~4 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[12]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[12]~4 .shared_arith = "off";

dffeas \A_slow_inst_result[12] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[12]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[12]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[12] .is_wysiwyg = "true";
defparam \A_slow_inst_result[12] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[12]~12 (
	.dataa(!\A_inst_result[12]~q ),
	.datab(!\A_inst_result[28]~q ),
	.datac(!\A_slow_inst_result[12]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[12]~12 .extended_lut = "off";
defparam \A_wr_data_unfiltered[12]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[12]~13 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[12]~q ),
	.datad(!\A_shift_rot_result[12]~q ),
	.datae(!\A_wr_data_unfiltered[12]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[12]~13 .extended_lut = "off";
defparam \A_wr_data_unfiltered[12]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[12]~13 .shared_arith = "off";

dffeas \W_wr_data[12] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[12]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[12]~q ),
	.prn(vcc));
defparam \W_wr_data[12] .is_wysiwyg = "true";
defparam \W_wr_data[12] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[12]~14 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[12]~q ),
	.datae(!\A_shift_rot_result[12]~q ),
	.dataf(!\A_wr_data_unfiltered[12]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~14 .extended_lut = "off";
defparam \D_src2_reg[12]~14 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[12]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[12]~91 (
	.dataa(!\M_alu_result[12]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[12]~q ),
	.dataf(!\D_src2_reg[12]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~91 .extended_lut = "off";
defparam \D_src2_reg[12]~91 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[12]~91 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[12]~0 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[12]~q ),
	.datad(!\E_src1[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[12]~0 .extended_lut = "off";
defparam \E_logic_result[12]~0 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[12]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~4 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[12]~0_combout ),
	.datad(!\E_extra_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~4 .extended_lut = "off";
defparam \E_alu_result[12]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[12]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[12]~127 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\D_src2_reg[12]~91_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[12]~4_combout ),
	.datag(!\Add24~41_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~127_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~127 .extended_lut = "on";
defparam \D_src2_reg[12]~127 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[12]~127 .shared_arith = "off";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(\D_src2_reg[12]~127_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[12] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~41_sumout ),
	.datac(!\E_alu_result[12]~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12] .extended_lut = "off";
defparam \E_alu_result[12] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[12] .shared_arith = "off";

dffeas \M_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[12]~q ),
	.prn(vcc));
defparam \M_alu_result[12] .is_wysiwyg = "true";
defparam \M_alu_result[12] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[12]~3 (
	.dataa(!\M_alu_result[12]~q ),
	.datab(!\A_wr_data_unfiltered[12]~13_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\W_wr_data[12]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[12]~3 .extended_lut = "off";
defparam \D_src1_reg[12]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[12]~3 .shared_arith = "off";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\D_src1_reg[12]~3_combout ),
	.asdata(\E_alu_result[12]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[13]~23 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_src1[11]~q ),
	.datad(!\E_src1[10]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[13]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[13]~23 .extended_lut = "off";
defparam \E_rot_step1[13]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[13]~23 .shared_arith = "off";

dffeas \M_rot_prestep2[17] (
	.clk(clk_clk),
	.d(\E_rot_step1[13]~23_combout ),
	.asdata(\E_rot_step1[17]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[17]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[17] .is_wysiwyg = "true";
defparam \M_rot_prestep2[17] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~24 (
	.dataa(!\M_rot_prestep2[17]~q ),
	.datab(!\M_rot_prestep2[9]~q ),
	.datac(!\M_rot_prestep2[1]~q ),
	.datad(!\M_rot_prestep2[25]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~24 .extended_lut = "off";
defparam \M_rot[1]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~24 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~24 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[1]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~24 .extended_lut = "off";
defparam \A_shift_rot_result~24 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~24 .shared_arith = "off";

dffeas \A_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[17] .is_wysiwyg = "true";
defparam \A_shift_rot_result[17] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[17]~24 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\A_slow_ld_data_fill_bit~0_combout ),
	.datac(!\d_readdata_d1[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[17]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[17]~24 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[17]~24 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[17]~24 .shared_arith = "off";

dffeas \A_slow_inst_result[17] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[17]~24_combout ),
	.asdata(\A_div_quot[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[17]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[17] .is_wysiwyg = "true";
defparam \A_slow_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[17]~53 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[17]~q ),
	.dataf(!\A_slow_inst_result[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[17]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[17]~53 .extended_lut = "off";
defparam \A_wr_data_unfiltered[17]~53 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[17]~53 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[17]~54 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_wr_data_unfiltered[22]~26_combout ),
	.datac(!\A_mul_result[17]~q ),
	.datad(!\A_inst_result[17]~q ),
	.datae(!\A_wr_data_unfiltered[17]~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[17]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[17]~54 .extended_lut = "off";
defparam \A_wr_data_unfiltered[17]~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[17]~54 .shared_arith = "off";

dffeas \W_wr_data[17] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[17]~54_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[17]~q ),
	.prn(vcc));
defparam \W_wr_data[17] .is_wysiwyg = "true";
defparam \W_wr_data[17] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[17]~47 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\W_wr_data[17]~q ),
	.datad(!\A_wr_data_unfiltered[17]~54_combout ),
	.datae(!\M_alu_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~47 .extended_lut = "off";
defparam \D_src2_reg[17]~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[17]~47 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[17]~48 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\E_alu_result~24_combout ),
	.datad(!\Add24~105_sumout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~48 .extended_lut = "off";
defparam \D_src2_reg[17]~48 .lut_mask = 64'hFFFFF7D5FFFFF7D5;
defparam \D_src2_reg[17]~48 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~15 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\Equal300~0_combout ),
	.datac(!\D_iw[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~15 .extended_lut = "off";
defparam \D_src2[17]~15 .lut_mask = 64'h4747474747474747;
defparam \D_src2[17]~15 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~16 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_ctrl_src2_choose_imm~q ),
	.datad(!\D_src2_reg[17]~47_combout ),
	.datae(!\D_src2_reg[17]~48_combout ),
	.dataf(!\D_src2[17]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~16 .extended_lut = "off";
defparam \D_src2[17]~16 .lut_mask = 64'hFFFFDEFFFFFFFFFF;
defparam \D_src2[17]~16 .shared_arith = "off";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\D_src2[17]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~24 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[17]~q ),
	.datae(!\E_src1[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~24 .extended_lut = "off";
defparam \E_alu_result~24 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~24 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~24_combout ),
	.datac(!\Add24~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17] .extended_lut = "off";
defparam \E_alu_result[17] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[17] .shared_arith = "off";

dffeas \M_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[17]~q ),
	.prn(vcc));
defparam \M_alu_result[17] .is_wysiwyg = "true";
defparam \M_alu_result[17] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[17]~24 (
	.dataa(!\M_alu_result[17]~q ),
	.datab(!\A_wr_data_unfiltered[17]~54_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datad(!\W_wr_data[17]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[17]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[17]~24 .extended_lut = "off";
defparam \D_src1_reg[17]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[17]~24 .shared_arith = "off";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\D_src1_reg[17]~24_combout ),
	.asdata(\E_alu_result[17]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[17]~20 (
	.dataa(!\E_src1[17]~q ),
	.datab(!\E_src1[16]~q ),
	.datac(!\E_src1[15]~q ),
	.datad(!\E_src1[14]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[17]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[17]~20 .extended_lut = "off";
defparam \E_rot_step1[17]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[17]~20 .shared_arith = "off";

dffeas \M_rot_prestep2[21] (
	.clk(clk_clk),
	.d(\E_rot_step1[17]~20_combout ),
	.asdata(\E_rot_step1[21]~21_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[21]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[21] .is_wysiwyg = "true";
defparam \M_rot_prestep2[21] .power_up = "low";

dffeas \M_rot_prestep2[5] (
	.clk(clk_clk),
	.d(\E_rot_step1[1]~16_combout ),
	.asdata(\E_rot_step1[5]~17_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[5]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[5] .is_wysiwyg = "true";
defparam \M_rot_prestep2[5] .power_up = "low";

dffeas \M_rot_prestep2[29] (
	.clk(clk_clk),
	.d(\E_rot_step1[25]~18_combout ),
	.asdata(\E_rot_step1[29]~19_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[29]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[29] .is_wysiwyg = "true";
defparam \M_rot_prestep2[29] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~26 (
	.dataa(!\M_rot_prestep2[21]~q ),
	.datab(!\M_rot_prestep2[13]~q ),
	.datac(!\M_rot_prestep2[5]~q ),
	.datad(!\M_rot_prestep2[29]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~26 .extended_lut = "off";
defparam \M_rot[5]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~26 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~26 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[5]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~26 .extended_lut = "off";
defparam \A_shift_rot_result~26 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~26 .shared_arith = "off";

dffeas \A_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[21] .is_wysiwyg = "true";
defparam \A_shift_rot_result[21] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[21]~26 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[21]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[21]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[21]~26 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[21]~26 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[21]~26 .shared_arith = "off";

dffeas \A_slow_inst_result[21] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[21]~26_combout ),
	.asdata(\A_div_quot[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[21]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[21] .is_wysiwyg = "true";
defparam \A_slow_inst_result[21] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[21]~57 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[21]~q ),
	.dataf(!\A_slow_inst_result[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[21]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[21]~57 .extended_lut = "off";
defparam \A_wr_data_unfiltered[21]~57 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[21]~57 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[21]~58 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[21]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[21]~q ),
	.datae(!\A_wr_data_unfiltered[21]~57_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[21]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[21]~58 .extended_lut = "off";
defparam \A_wr_data_unfiltered[21]~58 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[21]~58 .shared_arith = "off";

dffeas \W_wr_data[21] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[21]~58_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[21]~q ),
	.prn(vcc));
defparam \W_wr_data[21] .is_wysiwyg = "true";
defparam \W_wr_data[21] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[21]~26 (
	.dataa(!\M_alu_result[21]~q ),
	.datab(!\A_wr_data_unfiltered[21]~58_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[21]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[21]~26 .extended_lut = "off";
defparam \D_src1_reg[21]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[21]~26 .shared_arith = "off";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\D_src1_reg[21]~26_combout ),
	.asdata(\E_alu_result[21]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[21]~51 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~26_combout ),
	.datad(!\Add24~113_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~51 .extended_lut = "off";
defparam \D_src2_reg[21]~51 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[21]~51 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~52 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\A_wr_data_unfiltered[21]~58_combout ),
	.dataf(!\M_alu_result[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~52 .extended_lut = "off";
defparam \D_src2_reg[21]~52 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[21]~52 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~19 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~19 .extended_lut = "off";
defparam \D_src2[21]~19 .lut_mask = 64'h5353535353535353;
defparam \D_src2[21]~19 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~20 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[21]~51_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datae(!\D_src2_reg[21]~52_combout ),
	.dataf(!\D_src2[21]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~20 .extended_lut = "off";
defparam \D_src2[21]~20 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[21]~20 .shared_arith = "off";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\D_src2[21]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[21]~14 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[21]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[21]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[21]~14 .extended_lut = "off";
defparam \E_logic_result[21]~14 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[21]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~26 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[21]~14_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~26 .extended_lut = "off";
defparam \E_alu_result~26 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~26 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~26_combout ),
	.datac(!\Add24~113_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21] .extended_lut = "off";
defparam \E_alu_result[21] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[21] .shared_arith = "off";

dffeas \M_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[21]~q ),
	.prn(vcc));
defparam \M_alu_result[21] .is_wysiwyg = "true";
defparam \M_alu_result[21] .power_up = "low";

dffeas \A_inst_result[21] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(\M_alu_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[21]~q ),
	.prn(vcc));
defparam \A_inst_result[21] .is_wysiwyg = "true";
defparam \A_inst_result[21] .power_up = "low";

dffeas \A_inst_result[13] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.asdata(\M_alu_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[13]~q ),
	.prn(vcc));
defparam \A_inst_result[13] .is_wysiwyg = "true";
defparam \A_inst_result[13] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[5]~8 (
	.dataa(!\A_inst_result[5]~q ),
	.datab(!\A_inst_result[21]~q ),
	.datac(!\A_inst_result[13]~q ),
	.datad(!\A_inst_result[29]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[5]~8 .extended_lut = "off";
defparam \A_wr_data_unfiltered[5]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[5]~8 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[5]~3 (
	.dataa(!\M_rot_prestep2[5]~q ),
	.datab(!\M_rot_prestep2[29]~q ),
	.datac(!\M_rot_prestep2[21]~q ),
	.datad(!\M_rot_prestep2[13]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~3 .extended_lut = "off";
defparam \M_rot[5]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~3 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[5]~q ),
	.datae(!\M_rot[5]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~3 .extended_lut = "off";
defparam \A_shift_rot_result~3 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~3 .shared_arith = "off";

dffeas \A_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[5] .is_wysiwyg = "true";
defparam \A_shift_rot_result[5] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[5]~9 (
	.dataa(!\A_slow_inst_result[5]~q ),
	.datab(!\A_wr_data_unfiltered[5]~8_combout ),
	.datac(!\A_mul_result[5]~q ),
	.datad(!\A_shift_rot_result[5]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[5]~9 .extended_lut = "off";
defparam \A_wr_data_unfiltered[5]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[5]~9 .shared_arith = "off";

dffeas \W_wr_data[5] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[5]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[5]~q ),
	.prn(vcc));
defparam \W_wr_data[5] .is_wysiwyg = "true";
defparam \W_wr_data[5] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[5]~11 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\A_wr_data_unfiltered[5]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~11 .extended_lut = "off";
defparam \D_src2_reg[5]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[5]~11 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~12 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[5]~11_combout ),
	.datad(!\E_alu_result[5]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~12 .extended_lut = "off";
defparam \D_src2_reg[5]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[5]~12 .shared_arith = "off";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(\D_src2_reg[5]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~3 (
	.dataa(!\E_src2[5]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~3 .extended_lut = "off";
defparam \E_alu_result~3 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5] (
	.dataa(!\Add24~17_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~3_combout ),
	.datae(!\E_extra_pc[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5] .extended_lut = "off";
defparam \E_alu_result[5] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[5] .shared_arith = "off";

dffeas \M_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[5]~q ),
	.prn(vcc));
defparam \M_alu_result[5] .is_wysiwyg = "true";
defparam \M_alu_result[5] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[5]~2 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\A_wr_data_unfiltered[5]~9_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[5]~2 .extended_lut = "off";
defparam \D_src1_reg[5]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[5]~2 .shared_arith = "off";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\D_src1_reg[5]~2_combout ),
	.asdata(\E_alu_result[5]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[5]~17 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src1[3]~q ),
	.datad(!\E_src1[2]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[5]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[5]~17 .extended_lut = "off";
defparam \E_rot_step1[5]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[5]~17 .shared_arith = "off";

dffeas \M_rot_prestep2[9] (
	.clk(clk_clk),
	.d(\E_rot_step1[5]~17_combout ),
	.asdata(\E_rot_step1[9]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[9]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[9] .is_wysiwyg = "true";
defparam \M_rot_prestep2[9] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~7 (
	.dataa(!\M_rot_prestep2[9]~q ),
	.datab(!\M_rot_prestep2[1]~q ),
	.datac(!\M_rot_prestep2[25]~q ),
	.datad(!\M_rot_prestep2[17]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~7 .extended_lut = "off";
defparam \M_rot[1]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~7 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[1]~q ),
	.datae(!\M_rot[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~7 .extended_lut = "off";
defparam \A_shift_rot_result~7 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~7 .shared_arith = "off";

dffeas \A_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[9] .is_wysiwyg = "true";
defparam \A_shift_rot_result[9] .power_up = "low";

dffeas \A_inst_result[9] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(\M_alu_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[9]~q ),
	.prn(vcc));
defparam \A_inst_result[9] .is_wysiwyg = "true";
defparam \A_inst_result[9] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[9]~7 (
	.dataa(!\d_readdata_d1[9]~q ),
	.datab(!\d_readdata_d1[25]~q ),
	.datac(!\A_div_quot[9]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[9]~7 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[9]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[9]~7 .shared_arith = "off";

dffeas \A_slow_inst_result[9] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[9]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[9]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[9] .is_wysiwyg = "true";
defparam \A_slow_inst_result[9] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[9]~18 (
	.dataa(!\A_inst_result[9]~q ),
	.datab(!\A_inst_result[25]~q ),
	.datac(!\A_slow_inst_result[9]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[9]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[9]~18 .extended_lut = "off";
defparam \A_wr_data_unfiltered[9]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[9]~18 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[9]~19 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[9]~q ),
	.datad(!\A_shift_rot_result[9]~q ),
	.datae(!\A_wr_data_unfiltered[9]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[9]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[9]~19 .extended_lut = "off";
defparam \A_wr_data_unfiltered[9]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[9]~19 .shared_arith = "off";

dffeas \W_wr_data[9] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[9]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[9]~q ),
	.prn(vcc));
defparam \W_wr_data[9] .is_wysiwyg = "true";
defparam \W_wr_data[9] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[9]~17 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[9]~q ),
	.datae(!\A_shift_rot_result[9]~q ),
	.dataf(!\A_wr_data_unfiltered[9]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~17 .extended_lut = "off";
defparam \D_src2_reg[9]~17 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[9]~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~94 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[9]~q ),
	.dataf(!\D_src2_reg[9]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~94 .extended_lut = "off";
defparam \D_src2_reg[9]~94 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[9]~94 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[9]~3 (
	.dataa(!\E_src2[9]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[9]~3 .extended_lut = "off";
defparam \E_logic_result[9]~3 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[9]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~7 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[9]~3_combout ),
	.datad(!\E_extra_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~7 .extended_lut = "off";
defparam \E_alu_result[9]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~115 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\D_src2_reg[9]~94_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[9]~7_combout ),
	.datag(!\Add24~5_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~115_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~115 .extended_lut = "on";
defparam \D_src2_reg[9]~115 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[9]~115 .shared_arith = "off";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(\D_src2_reg[9]~115_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[9] (
	.dataa(!\Add24~5_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[9]~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9] .extended_lut = "off";
defparam \E_alu_result[9] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[9] .shared_arith = "off";

dffeas \M_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[9]~q ),
	.prn(vcc));
defparam \M_alu_result[9] .is_wysiwyg = "true";
defparam \M_alu_result[9] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[9]~6 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\A_wr_data_unfiltered[9]~19_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\W_wr_data[9]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[9]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[9]~6 .extended_lut = "off";
defparam \D_src1_reg[9]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[9]~6 .shared_arith = "off";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\D_src1_reg[9]~6_combout ),
	.asdata(\E_alu_result[9]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[9]~22 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src1[7]~q ),
	.datad(!\E_src1[6]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[9]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[9]~22 .extended_lut = "off";
defparam \E_rot_step1[9]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[9]~22 .shared_arith = "off";

dffeas \M_rot_prestep2[13] (
	.clk(clk_clk),
	.d(\E_rot_step1[9]~22_combout ),
	.asdata(\E_rot_step1[13]~23_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[13]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[13] .is_wysiwyg = "true";
defparam \M_rot_prestep2[13] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~14 (
	.dataa(!\M_rot_prestep2[13]~q ),
	.datab(!\M_rot_prestep2[5]~q ),
	.datac(!\M_rot_prestep2[29]~q ),
	.datad(!\M_rot_prestep2[21]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~14 .extended_lut = "off";
defparam \M_rot[5]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~14 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~14 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[5]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~14 .extended_lut = "off";
defparam \A_shift_rot_result~14 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~14 .shared_arith = "off";

dffeas \A_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[13] .is_wysiwyg = "true";
defparam \A_shift_rot_result[13] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[13]~14 (
	.dataa(!\d_readdata_d1[13]~q ),
	.datab(!\d_readdata_d1[29]~q ),
	.datac(!\A_div_quot[13]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[13]~14 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[13]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[13]~14 .shared_arith = "off";

dffeas \A_slow_inst_result[13] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[13]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[13]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[13] .is_wysiwyg = "true";
defparam \A_slow_inst_result[13] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[13]~33 (
	.dataa(!\A_inst_result[13]~q ),
	.datab(!\A_inst_result[29]~q ),
	.datac(!\A_slow_inst_result[13]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[13]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[13]~33 .extended_lut = "off";
defparam \A_wr_data_unfiltered[13]~33 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[13]~33 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[13]~34 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[13]~q ),
	.datad(!\A_shift_rot_result[13]~q ),
	.datae(!\A_wr_data_unfiltered[13]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[13]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[13]~34 .extended_lut = "off";
defparam \A_wr_data_unfiltered[13]~34 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[13]~34 .shared_arith = "off";

dffeas \W_wr_data[13] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[13]~34_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[13]~q ),
	.prn(vcc));
defparam \W_wr_data[13] .is_wysiwyg = "true";
defparam \W_wr_data[13] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[13]~27 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[13]~q ),
	.datae(!\A_shift_rot_result[13]~q ),
	.dataf(!\A_wr_data_unfiltered[13]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~27 .extended_lut = "off";
defparam \D_src2_reg[13]~27 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[13]~27 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[13]~98 (
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[13]~q ),
	.dataf(!\D_src2_reg[13]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~98 .extended_lut = "off";
defparam \D_src2_reg[13]~98 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[13]~98 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[13]~8 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[13]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[13]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[13]~8 .extended_lut = "off";
defparam \E_logic_result[13]~8 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[13]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13]~14 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[13]~8_combout ),
	.datad(!\E_extra_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~14 .extended_lut = "off";
defparam \E_alu_result[13]~14 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[13]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[13]~99 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\D_src2_reg[13]~98_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[13]~14_combout ),
	.datag(!\Add24~61_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~99_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~99 .extended_lut = "on";
defparam \D_src2_reg[13]~99 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[13]~99 .shared_arith = "off";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(\D_src2_reg[13]~99_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[13] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~61_sumout ),
	.datac(!\E_alu_result[13]~14_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13] .extended_lut = "off";
defparam \E_alu_result[13] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[13] .shared_arith = "off";

dffeas \M_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[13]~q ),
	.prn(vcc));
defparam \M_alu_result[13] .is_wysiwyg = "true";
defparam \M_alu_result[13] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[13]~13 (
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\A_wr_data_unfiltered[13]~34_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\W_wr_data[13]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[13]~13 .extended_lut = "off";
defparam \D_src1_reg[13]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[13]~13 .shared_arith = "off";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\D_src1_reg[13]~13_combout ),
	.asdata(\E_alu_result[13]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[14]~12 (
	.dataa(!\E_src1[14]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[14]~12 .extended_lut = "off";
defparam \E_rot_step1[14]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[14]~12 .shared_arith = "off";

dffeas \M_rot_prestep2[18] (
	.clk(clk_clk),
	.d(\E_rot_step1[14]~12_combout ),
	.asdata(\E_rot_step1[18]~13_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[18]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[18] .is_wysiwyg = "true";
defparam \M_rot_prestep2[18] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~28 (
	.dataa(!\M_rot_prestep2[18]~q ),
	.datab(!\M_rot_prestep2[10]~q ),
	.datac(!\M_rot_prestep2[2]~q ),
	.datad(!\M_rot_prestep2[26]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~28 .extended_lut = "off";
defparam \M_rot[2]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~28 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~28 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[2]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~28 .extended_lut = "off";
defparam \A_shift_rot_result~28 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~28 .shared_arith = "off";

dffeas \A_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[18] .is_wysiwyg = "true";
defparam \A_shift_rot_result[18] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[18]~28 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[18]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[18]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[18]~28 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[18]~28 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[18]~28 .shared_arith = "off";

dffeas \A_slow_inst_result[18] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[18]~28_combout ),
	.asdata(\A_div_quot[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[18]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[18] .is_wysiwyg = "true";
defparam \A_slow_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[18]~61 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[18]~q ),
	.dataf(!\A_slow_inst_result[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[18]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[18]~61 .extended_lut = "off";
defparam \A_wr_data_unfiltered[18]~61 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[18]~61 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[18]~62 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[18]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[18]~q ),
	.datae(!\A_wr_data_unfiltered[18]~61_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[18]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[18]~62 .extended_lut = "off";
defparam \A_wr_data_unfiltered[18]~62 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[18]~62 .shared_arith = "off";

dffeas \W_wr_data[18] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[18]~62_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[18]~q ),
	.prn(vcc));
defparam \W_wr_data[18] .is_wysiwyg = "true";
defparam \W_wr_data[18] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[18]~54 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\W_wr_data[18]~q ),
	.datad(!\A_wr_data_unfiltered[18]~62_combout ),
	.datae(!\M_alu_result[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~54 .extended_lut = "off";
defparam \D_src2_reg[18]~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[18]~54 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~55 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\E_alu_result~28_combout ),
	.datad(!\Add24~121_sumout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~55 .extended_lut = "off";
defparam \D_src2_reg[18]~55 .lut_mask = 64'hFFFFF7D5FFFFF7D5;
defparam \D_src2_reg[18]~55 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~22 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~22 .extended_lut = "off";
defparam \D_src2[18]~22 .lut_mask = 64'h5353535353535353;
defparam \D_src2[18]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~23 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_ctrl_src2_choose_imm~q ),
	.datad(!\D_src2_reg[18]~54_combout ),
	.datae(!\D_src2_reg[18]~55_combout ),
	.dataf(!\D_src2[18]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~23 .extended_lut = "off";
defparam \D_src2[18]~23 .lut_mask = 64'hFFFFDEFFFFFFFFFF;
defparam \D_src2[18]~23 .shared_arith = "off";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\D_src2[18]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~28 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[18]~q ),
	.datae(!\E_src1[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~28 .extended_lut = "off";
defparam \E_alu_result~28 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~28 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~28_combout ),
	.datac(!\Add24~121_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18] .extended_lut = "off";
defparam \E_alu_result[18] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[18] .shared_arith = "off";

dffeas \M_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[18]~q ),
	.prn(vcc));
defparam \M_alu_result[18] .is_wysiwyg = "true";
defparam \M_alu_result[18] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[18]~28 (
	.dataa(!\M_alu_result[18]~q ),
	.datab(!\A_wr_data_unfiltered[18]~62_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datad(!\W_wr_data[18]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[18]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[18]~28 .extended_lut = "off";
defparam \D_src1_reg[18]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[18]~28 .shared_arith = "off";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\D_src1_reg[18]~28_combout ),
	.asdata(\E_alu_result[18]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[18]~13 (
	.dataa(!\E_src1[18]~q ),
	.datab(!\E_src1[17]~q ),
	.datac(!\E_src1[16]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[18]~13 .extended_lut = "off";
defparam \E_rot_step1[18]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[18]~13 .shared_arith = "off";

dffeas \M_rot_prestep2[22] (
	.clk(clk_clk),
	.d(\E_rot_step1[18]~13_combout ),
	.asdata(\E_rot_step1[22]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[22]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[22] .is_wysiwyg = "true";
defparam \M_rot_prestep2[22] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~25 (
	.dataa(!\M_rot_prestep2[22]~q ),
	.datab(!\M_rot_prestep2[14]~q ),
	.datac(!\M_rot_prestep2[6]~q ),
	.datad(!\M_rot_prestep2[30]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~25 .extended_lut = "off";
defparam \M_rot[6]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~25 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~25 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[6]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~25 .extended_lut = "off";
defparam \A_shift_rot_result~25 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~25 .shared_arith = "off";

dffeas \A_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[22] .is_wysiwyg = "true";
defparam \A_shift_rot_result[22] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[22]~25 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\A_slow_ld_data_fill_bit~0_combout ),
	.datac(!\d_readdata_d1[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[22]~25 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[22]~25 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[22]~25 .shared_arith = "off";

dffeas \A_slow_inst_result[22] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[22]~25_combout ),
	.asdata(\A_div_quot[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[22]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[22] .is_wysiwyg = "true";
defparam \A_slow_inst_result[22] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~55 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[22]~q ),
	.dataf(!\A_slow_inst_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~55 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~55 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[22]~55 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~56 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[22]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[22]~q ),
	.datae(!\A_wr_data_unfiltered[22]~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~56 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~56 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[22]~56 .shared_arith = "off";

dffeas \W_wr_data[22] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[22]~56_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[22]~q ),
	.prn(vcc));
defparam \W_wr_data[22] .is_wysiwyg = "true";
defparam \W_wr_data[22] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[22]~25 (
	.dataa(!\M_alu_result[22]~q ),
	.datab(!\A_wr_data_unfiltered[22]~56_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[22]~25 .extended_lut = "off";
defparam \D_src1_reg[22]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[22]~25 .shared_arith = "off";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\D_src1_reg[22]~25_combout ),
	.asdata(\E_alu_result[22]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[22]~49 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~25_combout ),
	.datad(!\Add24~109_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~49 .extended_lut = "off";
defparam \D_src2_reg[22]~49 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[22]~49 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~50 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\A_wr_data_unfiltered[22]~56_combout ),
	.dataf(!\M_alu_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~50 .extended_lut = "off";
defparam \D_src2_reg[22]~50 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[22]~50 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~17 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\Equal300~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~17 .extended_lut = "off";
defparam \D_src2[22]~17 .lut_mask = 64'h5353535353535353;
defparam \D_src2[22]~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~18 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[22]~49_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datae(!\D_src2_reg[22]~50_combout ),
	.dataf(!\D_src2[22]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~18 .extended_lut = "off";
defparam \D_src2[22]~18 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[22]~18 .shared_arith = "off";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\D_src2[22]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[22]~13 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[22]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[22]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[22]~13 .extended_lut = "off";
defparam \E_logic_result[22]~13 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[22]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~25 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[22]~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~25 .extended_lut = "off";
defparam \E_alu_result~25 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~25 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~25_combout ),
	.datac(!\Add24~109_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22] .extended_lut = "off";
defparam \E_alu_result[22] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[22] .shared_arith = "off";

dffeas \M_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[22]~q ),
	.prn(vcc));
defparam \M_alu_result[22] .is_wysiwyg = "true";
defparam \M_alu_result[22] .power_up = "low";

dffeas \A_inst_result[22] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(\M_alu_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[22]~q ),
	.prn(vcc));
defparam \A_inst_result[22] .is_wysiwyg = "true";
defparam \A_inst_result[22] .power_up = "low";

dffeas \A_inst_result[14] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.asdata(\M_alu_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[14]~q ),
	.prn(vcc));
defparam \A_inst_result[14] .is_wysiwyg = "true";
defparam \A_inst_result[14] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~24 (
	.dataa(!\A_inst_result[6]~q ),
	.datab(!\A_inst_result[22]~q ),
	.datac(!\A_inst_result[14]~q ),
	.datad(!\A_inst_result[30]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~24 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[6]~24 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[6]~10 (
	.dataa(!\M_rot_prestep2[6]~q ),
	.datab(!\M_rot_prestep2[30]~q ),
	.datac(!\M_rot_prestep2[22]~q ),
	.datad(!\M_rot_prestep2[14]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~10 .extended_lut = "off";
defparam \M_rot[6]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~10 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[6]~q ),
	.datae(!\M_rot[6]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~10 .extended_lut = "off";
defparam \A_shift_rot_result~10 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~10 .shared_arith = "off";

dffeas \A_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[6] .is_wysiwyg = "true";
defparam \A_shift_rot_result[6] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~25 (
	.dataa(!\A_slow_inst_result[6]~q ),
	.datab(!\A_wr_data_unfiltered[6]~24_combout ),
	.datac(!\A_mul_result[6]~q ),
	.datad(!\A_shift_rot_result[6]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~25 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[6]~25 .shared_arith = "off";

dffeas \W_wr_data[6] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[6]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[6]~q ),
	.prn(vcc));
defparam \W_wr_data[6] .is_wysiwyg = "true";
defparam \W_wr_data[6] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[6]~21 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\A_wr_data_unfiltered[6]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~21 .extended_lut = "off";
defparam \D_src2_reg[6]~21 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[6]~21 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[6]~22 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[6]~21_combout ),
	.datad(!\E_alu_result[6]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~22 .extended_lut = "off";
defparam \D_src2_reg[6]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[6]~22 .shared_arith = "off";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(\D_src2_reg[6]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~10 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~10 .extended_lut = "off";
defparam \E_alu_result~10 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6] (
	.dataa(!\Add24~21_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~10_combout ),
	.datae(!\E_extra_pc[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6] .extended_lut = "off";
defparam \E_alu_result[6] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[6] .shared_arith = "off";

dffeas \M_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[6]~q ),
	.prn(vcc));
defparam \M_alu_result[6] .is_wysiwyg = "true";
defparam \M_alu_result[6] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[6]~9 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\A_wr_data_unfiltered[6]~25_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[6]~9 .extended_lut = "off";
defparam \D_src1_reg[6]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[6]~9 .shared_arith = "off";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\D_src1_reg[6]~9_combout ),
	.asdata(\E_alu_result[6]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[6]~14 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_src1[4]~q ),
	.datad(!\E_src1[3]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[6]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[6]~14 .extended_lut = "off";
defparam \E_rot_step1[6]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[6]~14 .shared_arith = "off";

dffeas \M_rot_prestep2[10] (
	.clk(clk_clk),
	.d(\E_rot_step1[6]~14_combout ),
	.asdata(\E_rot_step1[10]~15_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[10]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[10] .is_wysiwyg = "true";
defparam \M_rot_prestep2[10] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~6 (
	.dataa(!\M_rot_prestep2[10]~q ),
	.datab(!\M_rot_prestep2[2]~q ),
	.datac(!\M_rot_prestep2[26]~q ),
	.datad(!\M_rot_prestep2[18]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~6 .extended_lut = "off";
defparam \M_rot[2]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~6 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[2]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~6 .extended_lut = "off";
defparam \A_shift_rot_result~6 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~6 .shared_arith = "off";

dffeas \A_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[10] .is_wysiwyg = "true";
defparam \A_shift_rot_result[10] .power_up = "low";

dffeas \A_inst_result[10] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(\M_alu_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[10]~q ),
	.prn(vcc));
defparam \A_inst_result[10] .is_wysiwyg = "true";
defparam \A_inst_result[10] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[10]~6 (
	.dataa(!\d_readdata_d1[10]~q ),
	.datab(!\d_readdata_d1[26]~q ),
	.datac(!\A_div_quot[10]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[10]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[10]~6 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[10]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[10]~6 .shared_arith = "off";

dffeas \A_slow_inst_result[10] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[10]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[10]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[10] .is_wysiwyg = "true";
defparam \A_slow_inst_result[10] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[10]~16 (
	.dataa(!\A_inst_result[10]~q ),
	.datab(!\A_inst_result[26]~q ),
	.datac(!\A_slow_inst_result[10]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[10]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[10]~16 .extended_lut = "off";
defparam \A_wr_data_unfiltered[10]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[10]~16 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[10]~17 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[10]~q ),
	.datad(!\A_shift_rot_result[10]~q ),
	.datae(!\A_wr_data_unfiltered[10]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[10]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[10]~17 .extended_lut = "off";
defparam \A_wr_data_unfiltered[10]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[10]~17 .shared_arith = "off";

dffeas \W_wr_data[10] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[10]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[10]~q ),
	.prn(vcc));
defparam \W_wr_data[10] .is_wysiwyg = "true";
defparam \W_wr_data[10] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[10]~16 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[10]~q ),
	.datae(!\A_shift_rot_result[10]~q ),
	.dataf(!\A_wr_data_unfiltered[10]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~16 .extended_lut = "off";
defparam \D_src2_reg[10]~16 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[10]~16 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~93 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[10]~q ),
	.dataf(!\D_src2_reg[10]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~93 .extended_lut = "off";
defparam \D_src2_reg[10]~93 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[10]~93 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[10]~2 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[10]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[10]~2 .extended_lut = "off";
defparam \E_logic_result[10]~2 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[10]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~6 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[10]~2_combout ),
	.datad(!\E_extra_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~6 .extended_lut = "off";
defparam \E_alu_result[10]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[10]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~119 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\D_src2_reg[10]~93_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[10]~6_combout ),
	.datag(!\Add24~13_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~119_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~119 .extended_lut = "on";
defparam \D_src2_reg[10]~119 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[10]~119 .shared_arith = "off";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(\D_src2_reg[10]~119_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[10] (
	.dataa(!\Add24~13_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[10]~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10] .extended_lut = "off";
defparam \E_alu_result[10] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[10] .shared_arith = "off";

dffeas \M_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[10]~q ),
	.prn(vcc));
defparam \M_alu_result[10] .is_wysiwyg = "true";
defparam \M_alu_result[10] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[10]~5 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\A_wr_data_unfiltered[10]~17_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\W_wr_data[10]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[10]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[10]~5 .extended_lut = "off";
defparam \D_src1_reg[10]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[10]~5 .shared_arith = "off";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\D_src1_reg[10]~5_combout ),
	.asdata(\E_alu_result[10]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[10]~15 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_src1[8]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[10]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[10]~15 .extended_lut = "off";
defparam \E_rot_step1[10]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[10]~15 .shared_arith = "off";

dffeas \M_rot_prestep2[14] (
	.clk(clk_clk),
	.d(\E_rot_step1[10]~15_combout ),
	.asdata(\E_rot_step1[14]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[14]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[14] .is_wysiwyg = "true";
defparam \M_rot_prestep2[14] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~13 (
	.dataa(!\M_rot_prestep2[14]~q ),
	.datab(!\M_rot_prestep2[6]~q ),
	.datac(!\M_rot_prestep2[30]~q ),
	.datad(!\M_rot_prestep2[22]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~13 .extended_lut = "off";
defparam \M_rot[6]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~13 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~13 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[6]~q ),
	.datae(!\M_rot[6]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~13 .extended_lut = "off";
defparam \A_shift_rot_result~13 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~13 .shared_arith = "off";

dffeas \A_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[14] .is_wysiwyg = "true";
defparam \A_shift_rot_result[14] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[14]~13 (
	.dataa(!\d_readdata_d1[14]~q ),
	.datab(!\d_readdata_d1[30]~q ),
	.datac(!\A_div_quot[14]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[14]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[14]~13 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[14]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[14]~13 .shared_arith = "off";

dffeas \A_slow_inst_result[14] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[14]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[14]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[14] .is_wysiwyg = "true";
defparam \A_slow_inst_result[14] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[14]~31 (
	.dataa(!\A_inst_result[14]~q ),
	.datab(!\A_inst_result[30]~q ),
	.datac(!\A_slow_inst_result[14]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[14]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[14]~31 .extended_lut = "off";
defparam \A_wr_data_unfiltered[14]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[14]~31 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[14]~32 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[14]~q ),
	.datad(!\A_shift_rot_result[14]~q ),
	.datae(!\A_wr_data_unfiltered[14]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[14]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[14]~32 .extended_lut = "off";
defparam \A_wr_data_unfiltered[14]~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[14]~32 .shared_arith = "off";

dffeas \W_wr_data[14] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[14]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[14]~q ),
	.prn(vcc));
defparam \W_wr_data[14] .is_wysiwyg = "true";
defparam \W_wr_data[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[14]~26 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[14]~q ),
	.datae(!\A_shift_rot_result[14]~q ),
	.dataf(!\A_wr_data_unfiltered[14]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~26 .extended_lut = "off";
defparam \D_src2_reg[14]~26 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[14]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[14]~97 (
	.dataa(!\M_alu_result[14]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[14]~q ),
	.dataf(!\D_src2_reg[14]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~97_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~97 .extended_lut = "off";
defparam \D_src2_reg[14]~97 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[14]~97 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[14]~7 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[14]~q ),
	.datad(!\E_src1[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[14]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[14]~7 .extended_lut = "off";
defparam \E_logic_result[14]~7 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[14]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14]~13 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[14]~7_combout ),
	.datad(!\E_extra_pc[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14]~13 .extended_lut = "off";
defparam \E_alu_result[14]~13 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[14]~13 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[14]~103 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\D_src2_reg[14]~97_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[14]~13_combout ),
	.datag(!\Add24~57_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~103_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~103 .extended_lut = "on";
defparam \D_src2_reg[14]~103 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[14]~103 .shared_arith = "off";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(\D_src2_reg[14]~103_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[14] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~57_sumout ),
	.datac(!\E_alu_result[14]~13_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14] .extended_lut = "off";
defparam \E_alu_result[14] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[14] .shared_arith = "off";

dffeas \M_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[14]~q ),
	.prn(vcc));
defparam \M_alu_result[14] .is_wysiwyg = "true";
defparam \M_alu_result[14] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[14]~12 (
	.dataa(!\M_alu_result[14]~q ),
	.datab(!\A_wr_data_unfiltered[14]~32_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\W_wr_data[14]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[14]~12 .extended_lut = "off";
defparam \D_src1_reg[14]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[14]~12 .shared_arith = "off";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\D_src1_reg[14]~12_combout ),
	.asdata(\E_alu_result[14]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[15]~30 (
	.dataa(!\E_src1[15]~q ),
	.datab(!\E_src1[14]~q ),
	.datac(!\E_src1[13]~q ),
	.datad(!\E_src1[12]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[15]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[15]~30 .extended_lut = "off";
defparam \E_rot_step1[15]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[15]~30 .shared_arith = "off";

dffeas \M_rot_prestep2[19] (
	.clk(clk_clk),
	.d(\E_rot_step1[15]~30_combout ),
	.asdata(\E_rot_step1[19]~31_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[19]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[19] .is_wysiwyg = "true";
defparam \M_rot_prestep2[19] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~22 (
	.dataa(!\M_rot_prestep2[19]~q ),
	.datab(!\M_rot_prestep2[11]~q ),
	.datac(!\M_rot_prestep2[3]~q ),
	.datad(!\M_rot_prestep2[27]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~22 .extended_lut = "off";
defparam \M_rot[3]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~22 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~22 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[3]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~22 .extended_lut = "off";
defparam \A_shift_rot_result~22 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~22 .shared_arith = "off";

dffeas \A_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[19] .is_wysiwyg = "true";
defparam \A_shift_rot_result[19] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[19]~22 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[19]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[19]~22 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[19]~22 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[19]~22 .shared_arith = "off";

dffeas \A_slow_inst_result[19] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[19]~22_combout ),
	.asdata(\A_div_quot[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[19]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[19] .is_wysiwyg = "true";
defparam \A_slow_inst_result[19] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[19]~49 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[19]~q ),
	.dataf(!\A_slow_inst_result[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[19]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[19]~49 .extended_lut = "off";
defparam \A_wr_data_unfiltered[19]~49 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[19]~49 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[19]~50 (
	.dataa(!\A_inst_result[19]~q ),
	.datab(!\A_ctrl_mul_lsw~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[19]~q ),
	.datae(!\A_wr_data_unfiltered[19]~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[19]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[19]~50 .extended_lut = "off";
defparam \A_wr_data_unfiltered[19]~50 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \A_wr_data_unfiltered[19]~50 .shared_arith = "off";

dffeas \W_wr_data[19] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[19]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[19]~q ),
	.prn(vcc));
defparam \W_wr_data[19] .is_wysiwyg = "true";
defparam \W_wr_data[19] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[19]~89 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\A_wr_data_unfiltered[19]~50_combout ),
	.dataf(!\M_alu_result[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~89 .extended_lut = "off";
defparam \D_src2_reg[19]~89 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[19]~89 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~90 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~23_combout ),
	.datac(!\Add24~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~90 .extended_lut = "off";
defparam \D_src2_reg[19]~90 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \D_src2_reg[19]~90 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~44 (
	.dataa(!\D_src2_reg[0]~31_combout ),
	.datab(!\D_src2_reg[29]~1_combout ),
	.datac(!\D_src2_reg[29]~2_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datae(!\D_src2_reg[19]~89_combout ),
	.dataf(!\D_src2_reg[19]~90_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~44 .extended_lut = "off";
defparam \D_src2_reg[19]~44 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \D_src2_reg[19]~44 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[19]~14 (
	.dataa(!\D_iw[9]~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\Equal300~0_combout ),
	.datae(!\D_src2_reg[19]~44_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~14 .extended_lut = "off";
defparam \D_src2[19]~14 .lut_mask = 64'h7FDFFFFF7FDFFFFF;
defparam \D_src2[19]~14 .shared_arith = "off";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\D_src2[19]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~23 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[19]~q ),
	.datae(!\E_src1[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~23 .extended_lut = "off";
defparam \E_alu_result~23 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~23 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~23_combout ),
	.datac(!\Add24~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19] .extended_lut = "off";
defparam \E_alu_result[19] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[19] .shared_arith = "off";

dffeas \M_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[19]~q ),
	.prn(vcc));
defparam \M_alu_result[19] .is_wysiwyg = "true";
defparam \M_alu_result[19] .power_up = "low";

dffeas \A_inst_result[19] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(\M_alu_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[19]~q ),
	.prn(vcc));
defparam \A_inst_result[19] .is_wysiwyg = "true";
defparam \A_inst_result[19] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[3]~35 (
	.dataa(!\A_inst_result[3]~q ),
	.datab(!\A_inst_result[19]~q ),
	.datac(!\A_inst_result[11]~q ),
	.datad(!\A_inst_result[27]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[3]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[3]~35 .extended_lut = "off";
defparam \A_wr_data_unfiltered[3]~35 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[3]~35 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[3]~15 (
	.dataa(!\M_rot_prestep2[3]~q ),
	.datab(!\M_rot_prestep2[27]~q ),
	.datac(!\M_rot_prestep2[19]~q ),
	.datad(!\M_rot_prestep2[11]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~15 .extended_lut = "off";
defparam \M_rot[3]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~15 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~15 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_mask[3]~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[3]~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~15 .extended_lut = "off";
defparam \A_shift_rot_result~15 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~15 .shared_arith = "off";

dffeas \A_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[3] .is_wysiwyg = "true";
defparam \A_shift_rot_result[3] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[3]~36 (
	.dataa(!\A_slow_inst_result[3]~q ),
	.datab(!\A_wr_data_unfiltered[3]~35_combout ),
	.datac(!\A_mul_result[3]~q ),
	.datad(!\A_shift_rot_result[3]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[3]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[3]~36 .extended_lut = "off";
defparam \A_wr_data_unfiltered[3]~36 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[3]~36 .shared_arith = "off";

dffeas \W_wr_data[3] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[3]~36_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[3]~q ),
	.prn(vcc));
defparam \W_wr_data[3] .is_wysiwyg = "true";
defparam \W_wr_data[3] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[3]~14 (
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\A_wr_data_unfiltered[3]~36_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\W_wr_data[3]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[3]~14 .extended_lut = "off";
defparam \D_src1_reg[3]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[3]~14 .shared_arith = "off";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\D_src1_reg[3]~14_combout ),
	.asdata(\E_alu_result[3]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~15 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~15 .extended_lut = "off";
defparam \E_alu_result~15 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~15 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3] (
	.dataa(!\Add24~29_sumout ),
	.datab(!\E_alu_result~15_combout ),
	.datac(!\E_ctrl_retaddr~q ),
	.datad(!\E_extra_pc[1]~q ),
	.datae(!\E_alu_result~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3] .extended_lut = "off";
defparam \E_alu_result[3] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \E_alu_result[3] .shared_arith = "off";

dffeas \M_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[3]~q ),
	.prn(vcc));
defparam \M_alu_result[3] .is_wysiwyg = "true";
defparam \M_alu_result[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[3]~28 (
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\W_wr_data[3]~q ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\A_wr_data_unfiltered[3]~36_combout ),
	.datae(!\D_src2_reg[29]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~28 .extended_lut = "off";
defparam \D_src2_reg[3]~28 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \D_src2_reg[3]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[3]~29 (
	.dataa(!\D_src2_reg[3]~28_combout ),
	.datab(!\D_src2_reg[29]~1_combout ),
	.datac(!\D_src2_reg[29]~2_combout ),
	.datad(!\E_alu_result[3]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~29 .extended_lut = "off";
defparam \D_src2_reg[3]~29 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[3]~29 .shared_arith = "off";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\D_iw[9]~q ),
	.asdata(\D_src2_reg[3]~29_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass2~0 .extended_lut = "off";
defparam \E_rot_pass2~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass2~0 .shared_arith = "off";

dffeas M_rot_pass2(
	.clk(clk_clk),
	.d(\E_rot_pass2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass2~q ),
	.prn(vcc));
defparam M_rot_pass2.is_wysiwyg = "true";
defparam M_rot_pass2.power_up = "low";

cyclonev_lcell_comb \M_rot[4]~27 (
	.dataa(!\M_rot_prestep2[20]~q ),
	.datab(!\M_rot_prestep2[12]~q ),
	.datac(!\M_rot_prestep2[4]~q ),
	.datad(!\M_rot_prestep2[28]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~27 .extended_lut = "off";
defparam \M_rot[4]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~27 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~27 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[4]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~27 .extended_lut = "off";
defparam \A_shift_rot_result~27 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~27 .shared_arith = "off";

dffeas \A_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[20] .is_wysiwyg = "true";
defparam \A_shift_rot_result[20] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[20]~27 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[20]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[20]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[20]~27 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[20]~27 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[20]~27 .shared_arith = "off";

dffeas \A_slow_inst_result[20] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[20]~27_combout ),
	.asdata(\A_div_quot[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[20]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[20] .is_wysiwyg = "true";
defparam \A_slow_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[20]~59 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[20]~q ),
	.dataf(!\A_slow_inst_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[20]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[20]~59 .extended_lut = "off";
defparam \A_wr_data_unfiltered[20]~59 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[20]~59 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[20]~60 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[20]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[20]~q ),
	.datae(!\A_wr_data_unfiltered[20]~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[20]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[20]~60 .extended_lut = "off";
defparam \A_wr_data_unfiltered[20]~60 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[20]~60 .shared_arith = "off";

dffeas \W_wr_data[20] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[20]~60_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[20]~q ),
	.prn(vcc));
defparam \W_wr_data[20] .is_wysiwyg = "true";
defparam \W_wr_data[20] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[20]~87 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\A_wr_data_unfiltered[20]~60_combout ),
	.dataf(!\M_alu_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~87 .extended_lut = "off";
defparam \D_src2_reg[20]~87 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[20]~87 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~88 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~27_combout ),
	.datac(!\Add24~117_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~88 .extended_lut = "off";
defparam \D_src2_reg[20]~88 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \D_src2_reg[20]~88 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~53 (
	.dataa(!\D_src2_reg[0]~31_combout ),
	.datab(!\D_src2_reg[29]~1_combout ),
	.datac(!\D_src2_reg[29]~2_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datae(!\D_src2_reg[20]~87_combout ),
	.dataf(!\D_src2_reg[20]~88_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~53 .extended_lut = "off";
defparam \D_src2_reg[20]~53 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \D_src2_reg[20]~53 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~21 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\Equal300~0_combout ),
	.datae(!\D_src2_reg[20]~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~21 .extended_lut = "off";
defparam \D_src2[20]~21 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \D_src2[20]~21 .shared_arith = "off";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\D_src2[20]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~27 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[20]~q ),
	.datae(!\E_src1[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~27 .extended_lut = "off";
defparam \E_alu_result~27 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~27 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~27_combout ),
	.datac(!\Add24~117_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20] .extended_lut = "off";
defparam \E_alu_result[20] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[20] .shared_arith = "off";

dffeas \M_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[20]~q ),
	.prn(vcc));
defparam \M_alu_result[20] .is_wysiwyg = "true";
defparam \M_alu_result[20] .power_up = "low";

dffeas \A_inst_result[20] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(\M_alu_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[20]~q ),
	.prn(vcc));
defparam \A_inst_result[20] .is_wysiwyg = "true";
defparam \A_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[4]~0 (
	.dataa(!\A_inst_result[4]~q ),
	.datab(!\A_inst_result[20]~q ),
	.datac(!\A_inst_result[12]~q ),
	.datad(!\A_inst_result[28]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[4]~0 .extended_lut = "off";
defparam \A_wr_data_unfiltered[4]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[4]~0 (
	.dataa(!\M_rot_prestep2[4]~q ),
	.datab(!\M_rot_prestep2[28]~q ),
	.datac(!\M_rot_prestep2[20]~q ),
	.datad(!\M_rot_prestep2[12]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~0 .extended_lut = "off";
defparam \M_rot[4]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~0 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[4]~q ),
	.datae(!\M_rot[4]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~0 .extended_lut = "off";
defparam \A_shift_rot_result~0 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~0 .shared_arith = "off";

dffeas \A_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[4] .is_wysiwyg = "true";
defparam \A_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[4]~3 (
	.dataa(!\A_slow_inst_result[4]~q ),
	.datab(!\A_wr_data_unfiltered[4]~0_combout ),
	.datac(!\A_mul_result[4]~q ),
	.datad(!\A_shift_rot_result[4]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[4]~3 .extended_lut = "off";
defparam \A_wr_data_unfiltered[4]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[4]~3 .shared_arith = "off";

dffeas \W_wr_data[4] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[4]~q ),
	.prn(vcc));
defparam \W_wr_data[4] .is_wysiwyg = "true";
defparam \W_wr_data[4] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[4]~5 (
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\A_wr_data_unfiltered[4]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~5 .extended_lut = "off";
defparam \D_src2_reg[4]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[4]~6 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[4]~5_combout ),
	.datad(!\E_alu_result[4]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~6 .extended_lut = "off";
defparam \D_src2_reg[4]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[4]~6 .shared_arith = "off";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\D_iw[10]~q ),
	.asdata(\D_src2_reg[4]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~1 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~1 .extended_lut = "off";
defparam \E_alu_result~1 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4] (
	.dataa(!\Add24~33_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~1_combout ),
	.datae(!\E_extra_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4] .extended_lut = "off";
defparam \E_alu_result[4] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[4] .shared_arith = "off";

dffeas \M_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[4]~q ),
	.prn(vcc));
defparam \M_alu_result[4] .is_wysiwyg = "true";
defparam \M_alu_result[4] .power_up = "low";

dffeas \A_mem_baddr[4] (
	.clk(clk_clk),
	.d(\M_alu_result[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[4]~q ),
	.prn(vcc));
defparam \A_mem_baddr[4] .is_wysiwyg = "true";
defparam \A_mem_baddr[4] .power_up = "low";

dffeas M_sel_data_master(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_sel_data_master~q ),
	.prn(vcc));
defparam M_sel_data_master.is_wysiwyg = "true";
defparam M_sel_data_master.power_up = "low";

cyclonev_lcell_comb \M_ctrl_st_nxt~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_st_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_st_nxt~0 .extended_lut = "off";
defparam \M_ctrl_st_nxt~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \M_ctrl_st_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_st_cache~0 (
	.dataa(!\E_iw[5]~q ),
	.datab(!\Add24~37_sumout ),
	.datac(!\M_ctrl_st_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_cache~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_cache~0 .extended_lut = "off";
defparam \E_st_cache~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \E_st_cache~0 .shared_arith = "off";

dffeas M_ctrl_st_non_bypass(
	.clk(clk_clk),
	.d(\E_st_cache~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st_non_bypass~q ),
	.prn(vcc));
defparam M_ctrl_st_non_bypass.is_wysiwyg = "true";
defparam M_ctrl_st_non_bypass.power_up = "low";

cyclonev_lcell_comb \M_dc_valid_st_cache_hit~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_sel_data_master~q ),
	.datac(!\M_ctrl_st_non_bypass~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_cache_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_cache_hit~0 .extended_lut = "off";
defparam \M_dc_valid_st_cache_hit~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_valid_st_cache_hit~0 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_valid_st_cache_hit~1 (
	.dataa(!\M_dc_valid_st_cache_hit~0_combout ),
	.datab(!\M_dc_hit~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_cache_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_cache_hit~1 .extended_lut = "off";
defparam \M_dc_valid_st_cache_hit~1 .lut_mask = 64'h7777777777777777;
defparam \M_dc_valid_st_cache_hit~1 .shared_arith = "off";

dffeas A_dc_valid_st_cache_hit(
	.clk(clk_clk),
	.d(\M_dc_valid_st_cache_hit~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_valid_st_cache_hit~q ),
	.prn(vcc));
defparam A_dc_valid_st_cache_hit.is_wysiwyg = "true";
defparam A_dc_valid_st_cache_hit.power_up = "low";

dffeas \A_mem_baddr[10] (
	.clk(clk_clk),
	.d(\M_alu_result[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[10]~q ),
	.prn(vcc));
defparam \A_mem_baddr[10] .is_wysiwyg = "true";
defparam \A_mem_baddr[10] .power_up = "low";

dffeas \A_mem_baddr[7] (
	.clk(clk_clk),
	.d(\M_alu_result[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[7]~q ),
	.prn(vcc));
defparam \A_mem_baddr[7] .is_wysiwyg = "true";
defparam \A_mem_baddr[7] .power_up = "low";

dffeas \A_mem_baddr[5] (
	.clk(clk_clk),
	.d(\M_alu_result[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[5]~q ),
	.prn(vcc));
defparam \A_mem_baddr[5] .is_wysiwyg = "true";
defparam \A_mem_baddr[5] .power_up = "low";

dffeas \A_mem_baddr[6] (
	.clk(clk_clk),
	.d(\M_alu_result[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[6]~q ),
	.prn(vcc));
defparam \A_mem_baddr[6] .is_wysiwyg = "true";
defparam \A_mem_baddr[6] .power_up = "low";

cyclonev_lcell_comb \Equal261~0 (
	.dataa(!\A_mem_baddr[5]~q ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\A_mem_baddr[6]~q ),
	.datad(!\M_alu_result[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal261~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal261~0 .extended_lut = "off";
defparam \Equal261~0 .lut_mask = 64'h6996699669966996;
defparam \Equal261~0 .shared_arith = "off";

dffeas \A_mem_baddr[9] (
	.clk(clk_clk),
	.d(\M_alu_result[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[9]~q ),
	.prn(vcc));
defparam \A_mem_baddr[9] .is_wysiwyg = "true";
defparam \A_mem_baddr[9] .power_up = "low";

dffeas \A_mem_baddr[8] (
	.clk(clk_clk),
	.d(\M_alu_result[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[8]~q ),
	.prn(vcc));
defparam \A_mem_baddr[8] .is_wysiwyg = "true";
defparam \A_mem_baddr[8] .power_up = "low";

cyclonev_lcell_comb \Equal261~1 (
	.dataa(!\A_mem_baddr[9]~q ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\A_mem_baddr[8]~q ),
	.datad(!\M_alu_result[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal261~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal261~1 .extended_lut = "off";
defparam \Equal261~1 .lut_mask = 64'h6996699669966996;
defparam \Equal261~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal261~2 (
	.dataa(!\A_mem_baddr[10]~q ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\A_mem_baddr[7]~q ),
	.datad(!\M_alu_result[7]~q ),
	.datae(!\Equal261~0_combout ),
	.dataf(!\Equal261~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal261~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal261~2 .extended_lut = "off";
defparam \Equal261~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \Equal261~2 .shared_arith = "off";

cyclonev_lcell_comb M_dc_dirty(
	.dataa(!\A_dc_valid_st_cache_hit~q ),
	.datab(!\Equal261~2_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_dirty~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_dirty.extended_lut = "off";
defparam M_dc_dirty.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam M_dc_dirty.shared_arith = "off";

dffeas A_dc_dirty(
	.clk(clk_clk),
	.d(\M_dc_dirty~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_dirty~q ),
	.prn(vcc));
defparam A_dc_dirty.is_wysiwyg = "true";
defparam A_dc_dirty.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_has_started_nxt~0 (
	.dataa(!\A_dc_xfer_rd_addr_has_started~q ),
	.datab(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_has_started_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .shared_arith = "off";

dffeas A_dc_xfer_rd_addr_has_started(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_has_started_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_has_started~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_has_started.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_has_started.power_up = "low";

cyclonev_lcell_comb \Equal191~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal191~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal191~0 .extended_lut = "off";
defparam \Equal191~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \Equal191~0 .shared_arith = "off";

dffeas M_ctrl_dc_index_wb_inv(
	.clk(clk_clk),
	.d(\Equal191~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_index_wb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_index_wb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_index_wb_inv.power_up = "low";

dffeas A_ctrl_dc_index_wb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_index_wb_inv~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_index_wb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_index_wb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_index_wb_inv.power_up = "low";

dffeas A_dc_hit(
	.clk(clk_clk),
	.d(\M_dc_hit~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_hit~q ),
	.prn(vcc));
defparam A_dc_hit.is_wysiwyg = "true";
defparam A_dc_hit.power_up = "low";

cyclonev_lcell_comb \E_ctrl_dc_addr_inv~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_dc_addr_inv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_dc_addr_inv~0 .extended_lut = "off";
defparam \E_ctrl_dc_addr_inv~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \E_ctrl_dc_addr_inv~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal179~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_ctrl_dc_addr_inv~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal179~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal179~0 .extended_lut = "off";
defparam \Equal179~0 .lut_mask = 64'h7777777777777777;
defparam \Equal179~0 .shared_arith = "off";

dffeas M_ctrl_dc_addr_wb_inv(
	.clk(clk_clk),
	.d(\Equal179~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_addr_wb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_addr_wb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_addr_wb_inv.power_up = "low";

dffeas A_ctrl_dc_addr_wb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_addr_wb_inv~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_addr_wb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_addr_wb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_addr_wb_inv.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_starting~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_ctrl_dc_index_wb_inv~q ),
	.datac(!\A_dc_hit~q ),
	.datad(!\A_ctrl_dc_addr_wb_inv~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_starting~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_starting~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \A_dc_xfer_rd_addr_starting~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_starting~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_dirty~q ),
	.datad(!\A_dc_xfer_rd_addr_has_started~q ),
	.datae(!\A_dc_xfer_rd_addr_starting~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_starting~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_starting~1 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_starting~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \A_dc_xfer_rd_addr_starting~1 .shared_arith = "off";

dffeas A_dc_xfer_rd_data_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_starting~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_starting~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_starting.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_starting.power_up = "low";

dffeas A_dc_xfer_wr_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_data_starting~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_starting~q ),
	.prn(vcc));
defparam A_dc_xfer_wr_starting.is_wysiwyg = "true";
defparam A_dc_xfer_wr_starting.power_up = "low";

dffeas A_dc_wb_rd_addr_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_starting~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_addr_starting~q ),
	.prn(vcc));
defparam A_dc_wb_rd_addr_starting.is_wysiwyg = "true";
defparam A_dc_wb_rd_addr_starting.power_up = "low";

dffeas A_dc_wb_rd_data_starting(
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_starting~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_data_starting~q ),
	.prn(vcc));
defparam A_dc_wb_rd_data_starting.is_wysiwyg = "true";
defparam A_dc_wb_rd_data_starting.power_up = "low";

cyclonev_lcell_comb \A_dc_wb_rd_data_first_nxt~0 (
	.dataa(!d_read1),
	.datab(!\A_dc_wb_rd_data_first~q ),
	.datac(!\A_dc_wb_rd_data_starting~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_data_first_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_data_first_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_rd_data_first_nxt~0 .lut_mask = 64'h4747474747474747;
defparam \A_dc_wb_rd_data_first_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_rd_data_first(
	.clk(clk_clk),
	.d(\A_dc_wb_rd_data_first_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_data_first~q ),
	.prn(vcc));
defparam A_dc_wb_rd_data_first.is_wysiwyg = "true";
defparam A_dc_wb_rd_data_first.power_up = "low";

cyclonev_lcell_comb A_dc_wb_wr_starting(
	.dataa(!d_read1),
	.datab(!\A_dc_wb_rd_data_first~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_starting~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_wr_starting.extended_lut = "off";
defparam A_dc_wb_wr_starting.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam A_dc_wb_wr_starting.shared_arith = "off";

cyclonev_lcell_comb \av_wr_data_transfer~0 (
	.dataa(!rst1),
	.datab(!d_write1),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_wr_data_transfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_wr_data_transfer~0 .extended_lut = "off";
defparam \av_wr_data_transfer~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \av_wr_data_transfer~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[0]~3 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\av_wr_data_transfer~0_combout ),
	.datac(!\A_dc_wr_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[0]~3 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \A_dc_wr_data_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_wr_active_nxt~0 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(!\A_dc_wr_data_cnt[3]~q ),
	.datad(!\av_wr_data_transfer~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_wr_active_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_wr_active_nxt~0 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \A_dc_wb_wr_active_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_wr_active(
	.clk(clk_clk),
	.d(\A_dc_wb_wr_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_wr_active~q ),
	.prn(vcc));
defparam A_dc_wb_wr_active.is_wysiwyg = "true";
defparam A_dc_wb_wr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt[0]~0 (
	.dataa(!rst1),
	.datab(!d_write1),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(!\A_dc_wb_wr_starting~combout ),
	.dataf(!\A_dc_wb_wr_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt[0]~0 .extended_lut = "off";
defparam \A_dc_wr_data_cnt[0]~0 .lut_mask = 64'hFFFFFFFFFFF7FFFF;
defparam \A_dc_wr_data_cnt[0]~0 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[0]~0_combout ),
	.q(\A_dc_wr_data_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[1]~2 (
	.dataa(!\av_wr_data_transfer~0_combout ),
	.datab(!\A_dc_wr_data_cnt[1]~q ),
	.datac(!\A_dc_wr_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_dc_wr_data_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[0]~0_combout ),
	.q(\A_dc_wr_data_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[2]~1 (
	.dataa(!\av_wr_data_transfer~0_combout ),
	.datab(!\A_dc_wr_data_cnt[2]~q ),
	.datac(!\A_dc_wr_data_cnt[1]~q ),
	.datad(!\A_dc_wr_data_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \A_dc_wr_data_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[0]~0_combout ),
	.q(\A_dc_wr_data_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[3]~0 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!\av_wr_data_transfer~0_combout ),
	.datad(!\A_dc_wr_data_cnt[2]~q ),
	.datae(!\A_dc_wr_data_cnt[1]~q ),
	.dataf(!\A_dc_wr_data_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[3]~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \A_dc_wr_data_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[0]~0_combout ),
	.q(\A_dc_wr_data_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[3] .power_up = "low";

cyclonev_lcell_comb \A_dc_wb_active_nxt~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!\av_wr_data_transfer~0_combout ),
	.datad(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_active_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_active_nxt~0 .lut_mask = 64'hD8FFD8FFD8FFD8FF;
defparam \A_dc_wb_active_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_active(
	.clk(clk_clk),
	.d(\A_dc_wb_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_active~q ),
	.prn(vcc));
defparam A_dc_wb_active.is_wysiwyg = "true";
defparam A_dc_wb_active.power_up = "low";

cyclonev_lcell_comb \A_dc_fill_has_started_nxt~0 (
	.dataa(!\A_dc_fill_has_started~q ),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_has_started_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_has_started_nxt~0 .extended_lut = "off";
defparam \A_dc_fill_has_started_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_dc_fill_has_started_nxt~0 .shared_arith = "off";

dffeas A_dc_fill_has_started(
	.clk(clk_clk),
	.d(\A_dc_fill_has_started_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_has_started~q ),
	.prn(vcc));
defparam A_dc_fill_has_started.is_wysiwyg = "true";
defparam A_dc_fill_has_started.power_up = "low";

cyclonev_lcell_comb \A_dc_fill_starting~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_fill_has_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_starting~0 .extended_lut = "off";
defparam \A_dc_fill_starting~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \A_dc_fill_starting~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[0]~1 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_data_cnt[0]~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_fill_has_started~q ),
	.datad(!\d_readdatavalid_d1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt[0]~1 .extended_lut = "off";
defparam \A_dc_rd_data_cnt[0]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \A_dc_rd_data_cnt[0]~1 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[1]~2 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(!\A_dc_fill_dp_offset[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[1]~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[2]~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(!\A_dc_fill_dp_offset[1]~q ),
	.datad(!\A_dc_fill_dp_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[2]~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \Equal263~0 (
	.dataa(!\A_mem_baddr[4]~q ),
	.datab(!\A_dc_fill_dp_offset[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal263~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal263~0 .extended_lut = "off";
defparam \Equal263~0 .lut_mask = 64'h6666666666666666;
defparam \Equal263~0 .shared_arith = "off";

dffeas \A_mem_baddr[3] (
	.clk(clk_clk),
	.d(\M_alu_result[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[3]~q ),
	.prn(vcc));
defparam \A_mem_baddr[3] .is_wysiwyg = "true";
defparam \A_mem_baddr[3] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[0]~3 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\d_readdatavalid_d1~q ),
	.datac(!\A_dc_rd_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[0]~3 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \A_dc_rd_data_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_data_cnt[0]~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_fill_has_started~q ),
	.datad(!\A_dc_fill_active~q ),
	.datae(!\d_readdatavalid_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt[0]~0 .extended_lut = "off";
defparam \A_dc_rd_data_cnt[0]~0 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \A_dc_rd_data_cnt[0]~0 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[1]~2 (
	.dataa(!\d_readdatavalid_d1~q ),
	.datab(!\A_dc_rd_data_cnt[1]~q ),
	.datac(!\A_dc_rd_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_dc_rd_data_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[2]~1 (
	.dataa(!\d_readdatavalid_d1~q ),
	.datab(!\A_dc_rd_data_cnt[2]~q ),
	.datac(!\A_dc_rd_data_cnt[1]~q ),
	.datad(!\A_dc_rd_data_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \A_dc_rd_data_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[3]~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_rd_data_cnt[3]~q ),
	.datac(!\d_readdatavalid_d1~q ),
	.datad(!\A_dc_rd_data_cnt[2]~q ),
	.datae(!\A_dc_rd_data_cnt[1]~q ),
	.dataf(!\A_dc_rd_data_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[3]~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \A_dc_rd_data_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[3] .power_up = "low";

cyclonev_lcell_comb A_ld_bypass_done(
	.dataa(!\A_dc_rd_data_cnt[3]~q ),
	.datab(!\d_readdatavalid_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_done~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_ld_bypass_done.extended_lut = "off";
defparam A_ld_bypass_done.lut_mask = 64'h7777777777777777;
defparam A_ld_bypass_done.shared_arith = "off";

cyclonev_lcell_comb \M_ctrl_ld_st_nxt~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_ld_st_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_ld_st_nxt~0 .extended_lut = "off";
defparam \M_ctrl_ld_st_nxt~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \M_ctrl_ld_st_nxt~0 .shared_arith = "off";

dffeas M_ctrl_ld_st(
	.clk(clk_clk),
	.d(\M_ctrl_ld_st_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\E_iw[0]~q ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st~q ),
	.prn(vcc));
defparam M_ctrl_ld_st.is_wysiwyg = "true";
defparam M_ctrl_ld_st.power_up = "low";

cyclonev_lcell_comb \M_valid_mem_d1~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_ld_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_valid_mem_d1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_valid_mem_d1~0 .extended_lut = "off";
defparam \M_valid_mem_d1~0 .lut_mask = 64'h7777777777777777;
defparam \M_valid_mem_d1~0 .shared_arith = "off";

dffeas M_valid_mem_d1(
	.clk(clk_clk),
	.d(\M_valid_mem_d1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_valid_mem_d1~q ),
	.prn(vcc));
defparam M_valid_mem_d1.is_wysiwyg = "true";
defparam M_valid_mem_d1.power_up = "low";

dffeas M_A_dc_line_match_d1(
	.clk(clk_clk),
	.d(\Equal261~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_A_dc_line_match_d1~q ),
	.prn(vcc));
defparam M_A_dc_line_match_d1.is_wysiwyg = "true";
defparam M_A_dc_line_match_d1.power_up = "low";

cyclonev_lcell_comb A_dc_fill_need_extra_stall_nxt(
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\M_alu_result[4]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\M_valid_mem_d1~q ),
	.datae(!\M_A_dc_line_match_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_need_extra_stall_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_fill_need_extra_stall_nxt.extended_lut = "off";
defparam A_dc_fill_need_extra_stall_nxt.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam A_dc_fill_need_extra_stall_nxt.shared_arith = "off";

dffeas A_dc_fill_need_extra_stall(
	.clk(clk_clk),
	.d(\A_dc_fill_need_extra_stall_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_need_extra_stall~q ),
	.prn(vcc));
defparam A_dc_fill_need_extra_stall.is_wysiwyg = "true";
defparam A_dc_fill_need_extra_stall.power_up = "low";

dffeas A_dc_rd_last_transfer_d1(
	.clk(clk_clk),
	.d(\A_ld_bypass_done~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_rd_last_transfer_d1~q ),
	.prn(vcc));
defparam A_dc_rd_last_transfer_d1.is_wysiwyg = "true";
defparam A_dc_rd_last_transfer_d1.power_up = "low";

cyclonev_lcell_comb \A_dc_fill_active_nxt~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\A_ld_bypass_done~combout ),
	.datad(!\A_dc_fill_need_extra_stall~q ),
	.datae(!\A_dc_rd_last_transfer_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_active_nxt~0 .extended_lut = "off";
defparam \A_dc_fill_active_nxt~0 .lut_mask = 64'hFFFFF7FDFFFFF7FD;
defparam \A_dc_fill_active_nxt~0 .shared_arith = "off";

dffeas A_dc_fill_active(
	.clk(clk_clk),
	.d(\A_dc_fill_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_active~q ),
	.prn(vcc));
defparam A_dc_fill_active.is_wysiwyg = "true";
defparam A_dc_fill_active.power_up = "low";

dffeas \A_mem_baddr[2] (
	.clk(clk_clk),
	.d(\M_alu_result[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[2]~q ),
	.prn(vcc));
defparam \A_mem_baddr[2] .is_wysiwyg = "true";
defparam \A_mem_baddr[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_wr_data~0 (
	.dataa(!\A_mem_baddr[3]~q ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\A_mem_baddr[2]~q ),
	.datad(!\A_dc_fill_dp_offset[0]~q ),
	.datae(!\A_dc_fill_dp_offset[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_wr_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_wr_data~0 .extended_lut = "off";
defparam \A_dc_fill_wr_data~0 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \A_dc_fill_wr_data~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_en~0 (
	.dataa(!\A_ctrl_div~q ),
	.datab(!\d_readdatavalid_d1~q ),
	.datac(!\A_ctrl_ld_bypass~q ),
	.datad(!\Equal263~0_combout ),
	.datae(!\A_dc_fill_wr_data~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_en~0 .extended_lut = "off";
defparam \A_slow_inst_result_en~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \A_slow_inst_result_en~0 .shared_arith = "off";

dffeas \A_slow_inst_result[2] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[2]~2_combout ),
	.asdata(\A_div_quot[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[2]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[2] .is_wysiwyg = "true";
defparam \A_slow_inst_result[2] .power_up = "low";

dffeas \A_inst_result[2] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\M_alu_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[2]~q ),
	.prn(vcc));
defparam \A_inst_result[2] .is_wysiwyg = "true";
defparam \A_inst_result[2] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[2]~6 (
	.dataa(!\A_inst_result[2]~q ),
	.datab(!\A_inst_result[18]~q ),
	.datac(!\A_inst_result[10]~q ),
	.datad(!\A_inst_result[26]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[2]~6 .extended_lut = "off";
defparam \A_wr_data_unfiltered[2]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[2]~2 (
	.dataa(!\M_rot_prestep2[2]~q ),
	.datab(!\M_rot_prestep2[26]~q ),
	.datac(!\M_rot_prestep2[18]~q ),
	.datad(!\M_rot_prestep2[10]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~2 .extended_lut = "off";
defparam \M_rot[2]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~2 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[2]~q ),
	.datae(!\M_rot[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~2 .extended_lut = "off";
defparam \A_shift_rot_result~2 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~2 .shared_arith = "off";

dffeas \A_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[2] .is_wysiwyg = "true";
defparam \A_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[2]~7 (
	.dataa(!\A_slow_inst_result[2]~q ),
	.datab(!\A_wr_data_unfiltered[2]~6_combout ),
	.datac(!\A_mul_result[2]~q ),
	.datad(!\A_shift_rot_result[2]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[2]~7 .extended_lut = "off";
defparam \A_wr_data_unfiltered[2]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[2]~7 .shared_arith = "off";

dffeas \W_wr_data[2] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[2]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[2]~q ),
	.prn(vcc));
defparam \W_wr_data[2] .is_wysiwyg = "true";
defparam \W_wr_data[2] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[2]~1 (
	.dataa(!\M_alu_result[2]~q ),
	.datab(!\A_wr_data_unfiltered[2]~7_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[2]~1 .extended_lut = "off";
defparam \D_src1_reg[2]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[2]~1 .shared_arith = "off";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\D_src1_reg[2]~1_combout ),
	.asdata(\E_alu_result[2]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~2 .extended_lut = "off";
defparam \E_alu_result~2 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2] (
	.dataa(!\Add24~25_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~2_combout ),
	.datae(!\E_extra_pc[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2] .extended_lut = "off";
defparam \E_alu_result[2] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[2] .shared_arith = "off";

dffeas \M_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[2]~q ),
	.prn(vcc));
defparam \M_alu_result[2] .is_wysiwyg = "true";
defparam \M_alu_result[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[2]~9 (
	.dataa(!\M_alu_result[2]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\A_wr_data_unfiltered[2]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~9 .extended_lut = "off";
defparam \D_src2_reg[2]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[2]~10 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[2]~9_combout ),
	.datad(!\E_alu_result[2]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~10 .extended_lut = "off";
defparam \D_src2_reg[2]~10 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[2]~10 .shared_arith = "off";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(\D_src2_reg[2]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[5]~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[5]~3 .extended_lut = "off";
defparam \E_rot_mask[5]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[5]~3 .shared_arith = "off";

dffeas \M_rot_mask[5] (
	.clk(clk_clk),
	.d(\E_rot_mask[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[5]~q ),
	.prn(vcc));
defparam \M_rot_mask[5] .is_wysiwyg = "true";
defparam \M_rot_mask[5] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~16 (
	.dataa(!\M_rot_prestep2[29]~q ),
	.datab(!\M_rot_prestep2[21]~q ),
	.datac(!\M_rot_prestep2[13]~q ),
	.datad(!\M_rot_prestep2[5]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~16 .extended_lut = "off";
defparam \M_rot[5]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~16 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~16 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[5]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~16 .extended_lut = "off";
defparam \A_shift_rot_result~16 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~16 .shared_arith = "off";

dffeas \A_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[29] .is_wysiwyg = "true";
defparam \A_shift_rot_result[29] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[29]~16 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[29]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[29]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[29]~16 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[29]~16 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[29]~16 .shared_arith = "off";

dffeas \A_slow_inst_result[29] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[29]~16_combout ),
	.asdata(\A_div_quot[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[29]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[29] .is_wysiwyg = "true";
defparam \A_slow_inst_result[29] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~37 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[29]~q ),
	.dataf(!\A_slow_inst_result[29]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~37 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~37 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[29]~37 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~38 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[29]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[29]~q ),
	.datae(!\A_wr_data_unfiltered[29]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~38 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~38 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[29]~38 .shared_arith = "off";

dffeas \W_wr_data[29] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[29]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[29]~q ),
	.prn(vcc));
defparam \W_wr_data[29] .is_wysiwyg = "true";
defparam \W_wr_data[29] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[29]~15 (
	.dataa(!\M_alu_result[29]~q ),
	.datab(!\A_wr_data_unfiltered[29]~38_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[29]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[29]~15 .extended_lut = "off";
defparam \D_src1_reg[29]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[29]~15 .shared_arith = "off";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\D_src1_reg[29]~15_combout ),
	.asdata(\E_alu_result[29]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[29]~32 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~17_combout ),
	.datad(!\Add24~81_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~32 .extended_lut = "off";
defparam \D_src2_reg[29]~32 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[29]~32 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~33 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\A_wr_data_unfiltered[29]~38_combout ),
	.dataf(!\M_alu_result[29]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~33 .extended_lut = "off";
defparam \D_src2_reg[29]~33 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[29]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[29]~2 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\Equal300~0_combout ),
	.datac(!\D_iw[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~2 .extended_lut = "off";
defparam \D_src2[29]~2 .lut_mask = 64'h4747474747474747;
defparam \D_src2[29]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[29]~3 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[29]~32_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datae(!\D_src2_reg[29]~33_combout ),
	.dataf(!\D_src2[29]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~3 .extended_lut = "off";
defparam \D_src2[29]~3 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[29]~3 .shared_arith = "off";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\D_src2[29]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[29]~9 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[29]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[29]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[29]~9 .extended_lut = "off";
defparam \E_logic_result[29]~9 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[29]~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~0 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[26]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_src2[25]~q ),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~0 .extended_lut = "off";
defparam \Equal305~0 .lut_mask = 64'h6996966996696996;
defparam \Equal305~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~1 (
	.dataa(!\E_src2[0]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[19]~q ),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~1 .extended_lut = "off";
defparam \Equal305~1 .lut_mask = 64'h6996966996696996;
defparam \Equal305~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~2 (
	.dataa(!\E_logic_result[29]~9_combout ),
	.datab(!\E_logic_result[28]~10_combout ),
	.datac(!\E_logic_result[27]~11_combout ),
	.datad(!\E_logic_result[30]~12_combout ),
	.datae(!\Equal305~0_combout ),
	.dataf(!\Equal305~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~2 .extended_lut = "off";
defparam \Equal305~2 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal305~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~3 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src2[7]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~3 .extended_lut = "off";
defparam \Equal305~3 .lut_mask = 64'h6996966996696996;
defparam \Equal305~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~4 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src2[9]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~4 .extended_lut = "off";
defparam \Equal305~4 .lut_mask = 64'h6996966996696996;
defparam \Equal305~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~5 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[11]~q ),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~5 .extended_lut = "off";
defparam \Equal305~5 .lut_mask = 64'h6996966996696996;
defparam \Equal305~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~6 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[13]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(!\E_src2[12]~q ),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~6 .extended_lut = "off";
defparam \Equal305~6 .lut_mask = 64'h6996966996696996;
defparam \Equal305~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~7 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[16]~q ),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~7 .extended_lut = "off";
defparam \Equal305~7 .lut_mask = 64'h6996966996696996;
defparam \Equal305~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~8 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[15]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(!\E_src2[14]~q ),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~8 .extended_lut = "off";
defparam \Equal305~8 .lut_mask = 64'h6996966996696996;
defparam \Equal305~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~9 (
	.dataa(!\Equal305~3_combout ),
	.datab(!\Equal305~4_combout ),
	.datac(!\Equal305~5_combout ),
	.datad(!\Equal305~6_combout ),
	.datae(!\Equal305~7_combout ),
	.dataf(!\Equal305~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~9 .extended_lut = "off";
defparam \Equal305~9 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal305~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~10 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[17]~q ),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~10 .extended_lut = "off";
defparam \Equal305~10 .lut_mask = 64'h6996966996696996;
defparam \Equal305~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~11 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[20]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(!\E_src2[18]~q ),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~11 .extended_lut = "off";
defparam \Equal305~11 .lut_mask = 64'h6996966996696996;
defparam \Equal305~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~12 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[24]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(!\E_src2[23]~q ),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~12 .extended_lut = "off";
defparam \Equal305~12 .lut_mask = 64'h6996966996696996;
defparam \Equal305~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~13 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src2[5]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~13 .extended_lut = "off";
defparam \Equal305~13 .lut_mask = 64'h6996966996696996;
defparam \Equal305~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~14 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[31]~q ),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~14 .extended_lut = "off";
defparam \Equal305~14 .lut_mask = 64'h6996966996696996;
defparam \Equal305~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal305~15 (
	.dataa(!\E_logic_result[22]~13_combout ),
	.datab(!\E_logic_result[21]~14_combout ),
	.datac(!\Equal305~11_combout ),
	.datad(!\Equal305~12_combout ),
	.datae(!\Equal305~13_combout ),
	.dataf(!\Equal305~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal305~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal305~15 .extended_lut = "off";
defparam \Equal305~15 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal305~15 .shared_arith = "off";

dffeas \E_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_compare_op[1]~q ),
	.prn(vcc));
defparam \E_compare_op[1] .is_wysiwyg = "true";
defparam \E_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \E_br_result~0 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal305~2_combout ),
	.datac(!\Equal305~9_combout ),
	.datad(!\Equal305~10_combout ),
	.datae(!\Equal305~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~0 .extended_lut = "off";
defparam \E_br_result~0 .lut_mask = 64'hFFFFFFFF7DD7D77D;
defparam \E_br_result~0 .shared_arith = "off";

cyclonev_lcell_comb \E_br_result~1 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal305~2_combout ),
	.datac(!\Equal305~9_combout ),
	.datad(!\Equal305~10_combout ),
	.datae(!\Equal305~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~1 .extended_lut = "off";
defparam \E_br_result~1 .lut_mask = 64'hBEEBEBBEFFFFFFFF;
defparam \E_br_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[0]~15 (
	.dataa(!\E_src2[0]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[0]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[0]~15 .extended_lut = "off";
defparam \E_logic_result[0]~15 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[0]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0]~16 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_logic_result[0]~15_combout ),
	.datad(!\Add24~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0]~16 .extended_lut = "off";
defparam \E_alu_result[0]~16 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \E_alu_result[0]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0] (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\Add24~65_sumout ),
	.datac(!\E_br_result~0_combout ),
	.datad(!\E_br_result~1_combout ),
	.datae(!\E_alu_result[0]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0] .extended_lut = "off";
defparam \E_alu_result[0] .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \E_alu_result[0] .shared_arith = "off";

dffeas \M_alu_result[0] (
	.clk(clk_clk),
	.d(\E_alu_result[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[0]~q ),
	.prn(vcc));
defparam \M_alu_result[0] .is_wysiwyg = "true";
defparam \M_alu_result[0] .power_up = "low";

cyclonev_lcell_comb \M_ld_align_sh8~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\M_ctrl_ld8~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_sh8~0 .extended_lut = "off";
defparam \M_ld_align_sh8~0 .lut_mask = 64'h7777777777777777;
defparam \M_ld_align_sh8~0 .shared_arith = "off";

dffeas A_ld_align_sh8(
	.clk(clk_clk),
	.d(\M_ld_align_sh8~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_sh8~q ),
	.prn(vcc));
defparam A_ld_align_sh8.is_wysiwyg = "true";
defparam A_ld_align_sh8.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[1]~23 (
	.dataa(!\d_readdata_d1[1]~q ),
	.datab(!\d_readdata_d1[17]~q ),
	.datac(!\d_readdata_d1[9]~q ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[1]~23 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[1]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[1]~23 .shared_arith = "off";

dffeas \A_slow_inst_result[1] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[1]~23_combout ),
	.asdata(\A_div_quot[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[1]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[1] .is_wysiwyg = "true";
defparam \A_slow_inst_result[1] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[1]~1 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\M_ctrl_mem~q ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[1]~1 .extended_lut = "off";
defparam \M_inst_result[1]~1 .lut_mask = 64'h4747474747474747;
defparam \M_inst_result[1]~1 .shared_arith = "off";

dffeas A_ienable_reg_irq1(
	.clk(clk_clk),
	.d(\M_alu_result[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ienable_reg_irq0~0_combout ),
	.q(\A_ienable_reg_irq1~q ),
	.prn(vcc));
defparam A_ienable_reg_irq1.is_wysiwyg = "true";
defparam A_ienable_reg_irq1.power_up = "low";

cyclonev_lcell_comb A_ipending_reg_irq1_nxt(
	.dataa(!\A_ienable_reg_irq1~q ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_oci|the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_ienable[1]~q ),
	.datac(!irq_mask),
	.datad(!edge_capture),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ipending_reg_irq1_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_ipending_reg_irq1_nxt.extended_lut = "off";
defparam A_ipending_reg_irq1_nxt.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam A_ipending_reg_irq1_nxt.shared_arith = "off";

dffeas A_ipending_reg_irq1(
	.clk(clk_clk),
	.d(\A_ipending_reg_irq1_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_ipending_reg_irq1~q ),
	.prn(vcc));
defparam A_ipending_reg_irq1.is_wysiwyg = "true";
defparam A_ipending_reg_irq1.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[1]~2 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\A_ipending_reg_irq1~q ),
	.datad(!\D_iw[7]~q ),
	.datae(!\A_ienable_reg_irq1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[1]~2 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[1]~2 .lut_mask = 64'h9F6FFFFF9F6FFFFF;
defparam \D_control_reg_rddata_muxed[1]~2 .shared_arith = "off";

dffeas \E_control_reg_rddata[1] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_control_reg_rddata[1]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[1] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[1] .power_up = "low";

dffeas \M_control_reg_rddata[1] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_control_reg_rddata[1]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[1] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[1] .power_up = "low";

dffeas \A_inst_result[1] (
	.clk(clk_clk),
	.d(\M_inst_result[1]~1_combout ),
	.asdata(\M_control_reg_rddata[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_ctrl_rdctl_inst~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[1]~q ),
	.prn(vcc));
defparam \A_inst_result[1] .is_wysiwyg = "true";
defparam \A_inst_result[1] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[1]~51 (
	.dataa(!\A_inst_result[1]~q ),
	.datab(!\A_inst_result[17]~q ),
	.datac(!\A_inst_result[9]~q ),
	.datad(!\A_inst_result[25]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[1]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[1]~51 .extended_lut = "off";
defparam \A_wr_data_unfiltered[1]~51 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[1]~51 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[1]~23 (
	.dataa(!\M_rot_prestep2[1]~q ),
	.datab(!\M_rot_prestep2[25]~q ),
	.datac(!\M_rot_prestep2[17]~q ),
	.datad(!\M_rot_prestep2[9]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~23 .extended_lut = "off";
defparam \M_rot[1]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~23 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~23 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[1]~q ),
	.datae(!\M_rot[1]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~23 .extended_lut = "off";
defparam \A_shift_rot_result~23 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~23 .shared_arith = "off";

dffeas \A_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[1] .is_wysiwyg = "true";
defparam \A_shift_rot_result[1] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[1]~52 (
	.dataa(!\A_slow_inst_result[1]~q ),
	.datab(!\A_wr_data_unfiltered[1]~51_combout ),
	.datac(!\A_mul_result[1]~q ),
	.datad(!\A_shift_rot_result[1]~q ),
	.datae(!\A_wr_data_unfiltered[6]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[6]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[1]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[1]~52 .extended_lut = "off";
defparam \A_wr_data_unfiltered[1]~52 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[1]~52 .shared_arith = "off";

dffeas \W_wr_data[1] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[1]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[1]~q ),
	.prn(vcc));
defparam \W_wr_data[1] .is_wysiwyg = "true";
defparam \W_wr_data[1] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[1]~45 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\W_wr_data[1]~q ),
	.datad(!\A_wr_data_unfiltered[1]~52_combout ),
	.datae(!\M_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~45 .extended_lut = "off";
defparam \D_src2_reg[1]~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~45 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[1]~46 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[1]~45_combout ),
	.datad(!\E_alu_result[1]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~46 .extended_lut = "off";
defparam \D_src2_reg[1]~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~46 .shared_arith = "off";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(\D_src2_reg[1]~46_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[1]~16 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[1]~16 .extended_lut = "off";
defparam \E_logic_result[1]~16 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[1]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[1] (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add24~69_sumout ),
	.datad(!\E_logic_result[1]~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[1] .extended_lut = "off";
defparam \E_alu_result[1] .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \E_alu_result[1] .shared_arith = "off";

dffeas \M_alu_result[1] (
	.clk(clk_clk),
	.d(\E_alu_result[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[1]~q ),
	.prn(vcc));
defparam \M_alu_result[1] .is_wysiwyg = "true";
defparam \M_alu_result[1] .power_up = "low";

cyclonev_lcell_comb \M_data_ram_ld_align_sign_bit_16_hi~0 (
	.dataa(!\Add24~73_sumout ),
	.datab(!\Equal185~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_ram_ld_align_sign_bit_16_hi~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .extended_lut = "off";
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .lut_mask = 64'h7777777777777777;
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .shared_arith = "off";

dffeas M_data_ram_ld_align_sign_bit_16_hi(
	.clk(clk_clk),
	.d(\M_data_ram_ld_align_sign_bit_16_hi~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_data_ram_ld_align_sign_bit_16_hi~q ),
	.prn(vcc));
defparam M_data_ram_ld_align_sign_bit_16_hi.is_wysiwyg = "true";
defparam M_data_ram_ld_align_sign_bit_16_hi.power_up = "low";

cyclonev_lcell_comb \M_data_ram_ld_align_sign_bit~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\Qsys_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\M_alu_result[1]~q ),
	.dataf(!\M_data_ram_ld_align_sign_bit_16_hi~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_ram_ld_align_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_data_ram_ld_align_sign_bit~0 .extended_lut = "off";
defparam \M_data_ram_ld_align_sign_bit~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_data_ram_ld_align_sign_bit~0 .shared_arith = "off";

dffeas A_data_ram_ld_align_sign_bit(
	.clk(clk_clk),
	.d(\M_data_ram_ld_align_sign_bit~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_data_ram_ld_align_sign_bit~q ),
	.prn(vcc));
defparam A_data_ram_ld_align_sign_bit.is_wysiwyg = "true";
defparam A_data_ram_ld_align_sign_bit.power_up = "low";

cyclonev_lcell_comb \M_rot[0]~11 (
	.dataa(!\M_rot_prestep2[16]~q ),
	.datab(!\M_rot_prestep2[8]~q ),
	.datac(!\M_rot_prestep2[0]~q ),
	.datad(!\M_rot_prestep2[24]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~11 .extended_lut = "off";
defparam \M_rot[0]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~11 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~11 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[0]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~11 .extended_lut = "off";
defparam \A_shift_rot_result~11 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~11 .shared_arith = "off";

dffeas \A_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[16] .is_wysiwyg = "true";
defparam \A_shift_rot_result[16] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[16]~11 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[16]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[16]~11 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[16]~11 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[16]~11 .shared_arith = "off";

dffeas \A_slow_inst_result[16] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[16]~11_combout ),
	.asdata(\A_div_quot[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[16]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[16] .is_wysiwyg = "true";
defparam \A_slow_inst_result[16] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[16]~27 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[16]~q ),
	.dataf(!\A_slow_inst_result[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[16]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[16]~27 .extended_lut = "off";
defparam \A_wr_data_unfiltered[16]~27 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[16]~27 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[16]~28 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[16]~q ),
	.datac(!\A_mul_result[16]~q ),
	.datad(!\A_wr_data_unfiltered[22]~26_combout ),
	.datae(!\A_wr_data_unfiltered[16]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[16]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[16]~28 .extended_lut = "off";
defparam \A_wr_data_unfiltered[16]~28 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \A_wr_data_unfiltered[16]~28 .shared_arith = "off";

dffeas \W_wr_data[16] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[16]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[16]~q ),
	.prn(vcc));
defparam \W_wr_data[16] .is_wysiwyg = "true";
defparam \W_wr_data[16] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[16]~23 (
	.dataa(!\M_alu_result[16]~q ),
	.datab(!\D_src2_reg[29]~3_combout ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\W_wr_data[16]~q ),
	.datae(!\A_wr_data_unfiltered[16]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~23 .extended_lut = "off";
defparam \D_src2_reg[16]~23 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[16]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[16]~5 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[16]~q ),
	.datad(!\E_src1[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[16]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[16]~5 .extended_lut = "off";
defparam \E_logic_result[16]~5 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[16]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[16]~11 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[16]~5_combout ),
	.datad(!\E_extra_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16]~11 .extended_lut = "off";
defparam \E_alu_result[16]~11 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[16]~11 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[16]~24 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~49_sumout ),
	.datac(!\D_src2_reg[29]~2_combout ),
	.datad(!\E_alu_result[16]~11_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~24 .extended_lut = "off";
defparam \D_src2_reg[16]~24 .lut_mask = 64'hFFFFDFD5FFFFDFD5;
defparam \D_src2_reg[16]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~0 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\Equal300~0_combout ),
	.datac(!\D_iw[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~0 .extended_lut = "off";
defparam \D_src2[16]~0 .lut_mask = 64'h4747474747474747;
defparam \D_src2[16]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~1 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_ctrl_src2_choose_imm~q ),
	.datad(!\D_src2_reg[16]~23_combout ),
	.datae(!\D_src2_reg[16]~24_combout ),
	.dataf(!\D_src2[16]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~1 .extended_lut = "off";
defparam \D_src2[16]~1 .lut_mask = 64'hFFFFDEFFFFFFFFFF;
defparam \D_src2[16]~1 .shared_arith = "off";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\D_src2[16]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[18]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[16] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~49_sumout ),
	.datac(!\E_alu_result[16]~11_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16] .extended_lut = "off";
defparam \E_alu_result[16] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[16] .shared_arith = "off";

dffeas \M_alu_result[16] (
	.clk(clk_clk),
	.d(\E_alu_result[16]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[16]~q ),
	.prn(vcc));
defparam \M_alu_result[16] .is_wysiwyg = "true";
defparam \M_alu_result[16] .power_up = "low";

cyclonev_lcell_comb \M_dc_hit~0 (
	.dataa(!\M_alu_result[12]~q ),
	.datab(!\M_alu_result[11]~q ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[6] ),
	.datad(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_hit~0 .extended_lut = "off";
defparam \M_dc_hit~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \M_dc_hit~0 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_hit~1 (
	.dataa(!\M_alu_result[14]~q ),
	.datab(!\M_alu_result[13]~q ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_hit~1 .extended_lut = "off";
defparam \M_dc_hit~1 .lut_mask = 64'h6996699669966996;
defparam \M_dc_hit~1 .shared_arith = "off";

cyclonev_lcell_comb M_dc_hit(
	.dataa(!\M_alu_result[16]~q ),
	.datab(!\M_alu_result[15]~q ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datae(!\M_dc_hit~0_combout ),
	.dataf(!\M_dc_hit~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_hit~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_hit.extended_lut = "off";
defparam M_dc_hit.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam M_dc_hit.shared_arith = "off";

cyclonev_lcell_comb \M_dc_valid_st_bypass_hit~0 (
	.dataa(!\M_ctrl_st_bypass~q ),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_dc_hit~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_bypass_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_bypass_hit~0 .extended_lut = "off";
defparam \M_dc_valid_st_bypass_hit~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_valid_st_bypass_hit~0 .shared_arith = "off";

dffeas A_dc_valid_st_bypass_hit(
	.clk(clk_clk),
	.d(\M_dc_valid_st_bypass_hit~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_valid_st_bypass_hit~q ),
	.prn(vcc));
defparam A_dc_valid_st_bypass_hit.is_wysiwyg = "true";
defparam A_dc_valid_st_bypass_hit.power_up = "low";

cyclonev_lcell_comb A_st_bypass_transfer_done(
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!rst1),
	.datad(!d_write1),
	.datae(!suppress_change_dest_id),
	.dataf(!WideOr01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_transfer_done~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_st_bypass_transfer_done.extended_lut = "off";
defparam A_st_bypass_transfer_done.lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam A_st_bypass_transfer_done.shared_arith = "off";

dffeas A_st_bypass_transfer_done_d1(
	.clk(clk_clk),
	.d(\A_st_bypass_transfer_done~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_st_bypass_transfer_done_d1~q ),
	.prn(vcc));
defparam A_st_bypass_transfer_done_d1.is_wysiwyg = "true";
defparam A_st_bypass_transfer_done_d1.power_up = "low";

dffeas A_ctrl_st_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_st_bypass~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_st_bypass~q ),
	.prn(vcc));
defparam A_ctrl_st_bypass.is_wysiwyg = "true";
defparam A_ctrl_st_bypass.power_up = "low";

cyclonev_lcell_comb \E_ctrl_dc_nowb_inv~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_dc_nowb_inv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_dc_nowb_inv~0 .extended_lut = "off";
defparam \E_ctrl_dc_nowb_inv~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \E_ctrl_dc_nowb_inv~0 .shared_arith = "off";

dffeas M_ctrl_dc_nowb_inv(
	.clk(clk_clk),
	.d(\E_ctrl_dc_nowb_inv~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_nowb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_nowb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_nowb_inv.power_up = "low";

dffeas A_ctrl_dc_nowb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_nowb_inv~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_nowb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_nowb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_nowb_inv.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[0]~1 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[1]~0 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_active_nxt~0 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_done~q ),
	.datac(!\A_dc_xfer_rd_addr_active~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_active_nxt~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_active_nxt~0 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \A_dc_xfer_rd_addr_active_nxt~0 .shared_arith = "off";

dffeas A_dc_xfer_rd_addr_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_active~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_active.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[2]~2 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[2] .power_up = "low";

cyclonev_lcell_comb A_dc_xfer_rd_addr_done_nxt(
	.dataa(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(!\A_dc_xfer_rd_addr_active~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_done_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_xfer_rd_addr_done_nxt.extended_lut = "off";
defparam A_dc_xfer_rd_addr_done_nxt.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam A_dc_xfer_rd_addr_done_nxt.shared_arith = "off";

dffeas A_dc_xfer_rd_addr_done(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_done_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_done~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_done.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_done.power_up = "low";

cyclonev_lcell_comb \A_dc_dcache_management_done_nxt~0 (
	.dataa(!\A_dc_dirty~q ),
	.datab(!\A_ctrl_dc_index_wb_inv~q ),
	.datac(!\A_dc_hit~q ),
	.datad(!\A_ctrl_dc_addr_wb_inv~q ),
	.datae(!\A_ctrl_dc_nowb_inv~q ),
	.dataf(!\A_dc_xfer_rd_addr_done~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_dcache_management_done_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_dcache_management_done_nxt~0 .extended_lut = "off";
defparam \A_dc_dcache_management_done_nxt~0 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \A_dc_dcache_management_done_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_dcache_management_done_nxt(
	.dataa(!\A_valid~q ),
	.datab(!\A_stall~combout ),
	.datac(!\A_dc_dcache_management_done_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_dcache_management_done_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_dcache_management_done_nxt.extended_lut = "off";
defparam A_dc_dcache_management_done_nxt.lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam A_dc_dcache_management_done_nxt.shared_arith = "off";

dffeas A_dc_dcache_management_done(
	.clk(clk_clk),
	.d(\A_dc_dcache_management_done_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_dcache_management_done~q ),
	.prn(vcc));
defparam A_dc_dcache_management_done.is_wysiwyg = "true";
defparam A_dc_dcache_management_done.power_up = "low";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~0 (
	.dataa(!\E_valid~1_combout ),
	.datab(!\M_ctrl_mem_nxt~0_combout ),
	.datac(!\M_dc_valid_st_cache_hit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~1 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\Add24~1_sumout ),
	.datad(!\Add24~5_sumout ),
	.datae(!\M_dc_potential_hazard_after_st_unfiltered~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~2 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\Add24~17_sumout ),
	.datad(!\Add24~21_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .lut_mask = 64'h6996699669966996;
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~3 (
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\M_alu_result[4]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\Add24~25_sumout ),
	.datae(!\Add24~29_sumout ),
	.dataf(!\Add24~33_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .lut_mask = 64'h6996966996696996;
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~4 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\Add24~9_sumout ),
	.datad(!\Add24~13_sumout ),
	.datae(!\M_dc_potential_hazard_after_st_unfiltered~2_combout ),
	.dataf(!\M_dc_potential_hazard_after_st_unfiltered~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~5 (
	.dataa(!\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.datab(!\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .lut_mask = 64'h7777777777777777;
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .shared_arith = "off";

dffeas A_dc_potential_hazard_after_st(
	.clk(clk_clk),
	.d(\M_dc_potential_hazard_after_st_unfiltered~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_potential_hazard_after_st~q ),
	.prn(vcc));
defparam A_dc_potential_hazard_after_st.is_wysiwyg = "true";
defparam A_dc_potential_hazard_after_st.power_up = "low";

cyclonev_lcell_comb \A_mem_stall_nxt~1 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_ld_bypass_done~combout ),
	.datac(!\A_ctrl_ld_bypass~q ),
	.datad(!\A_dc_fill_need_extra_stall~q ),
	.datae(!\A_dc_rd_last_transfer_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~1 .extended_lut = "off";
defparam \A_mem_stall_nxt~1 .lut_mask = 64'h5F3FFFFF5F3FFFFF;
defparam \A_mem_stall_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~2 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_dc_dcache_management_done~q ),
	.datac(!\A_dc_valid_st_cache_hit~q ),
	.datad(!\A_dc_potential_hazard_after_st~q ),
	.datae(!\A_mem_stall_nxt~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~2 .extended_lut = "off";
defparam \A_mem_stall_nxt~2 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \A_mem_stall_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~3 (
	.dataa(!\A_dc_valid_st_bypass_hit~q ),
	.datab(!\A_st_bypass_transfer_done_d1~q ),
	.datac(!\A_ctrl_st_bypass~q ),
	.datad(!\A_st_bypass_transfer_done~combout ),
	.datae(!\A_mem_stall_nxt~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~3 .extended_lut = "off";
defparam \A_mem_stall_nxt~3 .lut_mask = 64'hFFD8FFFFFFD8FFFF;
defparam \A_mem_stall_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~4 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_stall~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~4 .extended_lut = "off";
defparam \A_mem_stall_nxt~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \A_mem_stall_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~5 (
	.dataa(!\A_mem_stall_nxt~0_combout ),
	.datab(!\A_mem_stall_nxt~3_combout ),
	.datac(!\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.datad(!\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.datae(!\M_dc_want_fill~combout ),
	.dataf(!\A_mem_stall_nxt~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~5 .extended_lut = "off";
defparam \A_mem_stall_nxt~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \A_mem_stall_nxt~5 .shared_arith = "off";

dffeas A_mem_stall(
	.clk(clk_clk),
	.d(\A_mem_stall_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mem_stall~q ),
	.prn(vcc));
defparam A_mem_stall.is_wysiwyg = "true";
defparam A_mem_stall.power_up = "low";

cyclonev_lcell_comb \always138~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_ctrl_div~q ),
	.datac(!\A_div_done~q ),
	.datad(!\A_mem_stall~q ),
	.datae(!\A_mul_stall~q ),
	.dataf(!\M_valid_from_E~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always138~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always138~0 .extended_lut = "off";
defparam \always138~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \always138~0 .shared_arith = "off";

cyclonev_lcell_comb \A_mul_cnt_nxt[0]~2 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[0]~2 .extended_lut = "off";
defparam \A_mul_cnt_nxt[0]~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \A_mul_cnt_nxt[0]~2 .shared_arith = "off";

dffeas \A_mul_cnt[0] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[0]~q ),
	.prn(vcc));
defparam \A_mul_cnt[0] .is_wysiwyg = "true";
defparam \A_mul_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_mul_cnt_nxt[1]~1 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[1]~q ),
	.datac(!\A_mul_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[1]~1 .extended_lut = "off";
defparam \A_mul_cnt_nxt[1]~1 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_mul_cnt_nxt[1]~1 .shared_arith = "off";

dffeas \A_mul_cnt[1] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[1]~q ),
	.prn(vcc));
defparam \A_mul_cnt[1] .is_wysiwyg = "true";
defparam \A_mul_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_mul_cnt_nxt[2]~0 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[2]~q ),
	.datac(!\A_mul_cnt[1]~q ),
	.datad(!\A_mul_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[2]~0 .extended_lut = "off";
defparam \A_mul_cnt_nxt[2]~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_mul_cnt_nxt[2]~0 .shared_arith = "off";

dffeas \A_mul_cnt[2] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[2]~q ),
	.prn(vcc));
defparam \A_mul_cnt[2] .is_wysiwyg = "true";
defparam \A_mul_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_mul_stall_nxt~0 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\always138~0_combout ),
	.datac(!\M_ctrl_mul_lsw~q ),
	.datad(!\A_mul_cnt[2]~q ),
	.datae(!\A_mul_cnt[1]~q ),
	.dataf(!\A_mul_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_stall_nxt~0 .extended_lut = "off";
defparam \A_mul_stall_nxt~0 .lut_mask = 64'hBFFFFFFF1FFFFFFF;
defparam \A_mul_stall_nxt~0 .shared_arith = "off";

dffeas A_mul_stall(
	.clk(clk_clk),
	.d(\A_mul_stall_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall~q ),
	.prn(vcc));
defparam A_mul_stall.is_wysiwyg = "true";
defparam A_mul_stall.power_up = "low";

dffeas A_mul_stall_d1(
	.clk(clk_clk),
	.d(\A_mul_stall~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d1~q ),
	.prn(vcc));
defparam A_mul_stall_d1.is_wysiwyg = "true";
defparam A_mul_stall_d1.power_up = "low";

dffeas A_mul_stall_d2(
	.clk(clk_clk),
	.d(\A_mul_stall_d1~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d2~q ),
	.prn(vcc));
defparam A_mul_stall_d2.is_wysiwyg = "true";
defparam A_mul_stall_d2.power_up = "low";

dffeas A_mul_stall_d3(
	.clk(clk_clk),
	.d(\A_mul_stall_d2~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d3~q ),
	.prn(vcc));
defparam A_mul_stall_d3.is_wysiwyg = "true";
defparam A_mul_stall_d3.power_up = "low";

dffeas \A_mul_result[0] (
	.clk(clk_clk),
	.d(\Add26~5_sumout ),
	.asdata(\A_mul_partial_prod[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[0]~q ),
	.prn(vcc));
defparam \A_mul_result[0] .is_wysiwyg = "true";
defparam \A_mul_result[0] .power_up = "low";

cyclonev_lcell_comb \Add26~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[1]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[1]~q ),
	.datag(gnd),
	.cin(\Add26~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~93_sumout ),
	.cout(\Add26~94 ),
	.shareout());
defparam \Add26~93 .extended_lut = "off";
defparam \Add26~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~93 .shared_arith = "off";

dffeas \A_mul_result[1] (
	.clk(clk_clk),
	.d(\Add26~93_sumout ),
	.asdata(\A_mul_partial_prod[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[1]~q ),
	.prn(vcc));
defparam \A_mul_result[1] .is_wysiwyg = "true";
defparam \A_mul_result[1] .power_up = "low";

cyclonev_lcell_comb \Add26~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[2]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[2]~q ),
	.datag(gnd),
	.cin(\Add26~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~9_sumout ),
	.cout(\Add26~10 ),
	.shareout());
defparam \Add26~9 .extended_lut = "off";
defparam \Add26~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~9 .shared_arith = "off";

dffeas \A_mul_result[2] (
	.clk(clk_clk),
	.d(\Add26~9_sumout ),
	.asdata(\A_mul_partial_prod[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[2]~q ),
	.prn(vcc));
defparam \A_mul_result[2] .is_wysiwyg = "true";
defparam \A_mul_result[2] .power_up = "low";

cyclonev_lcell_comb \Add26~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[3]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[3]~q ),
	.datag(gnd),
	.cin(\Add26~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~61_sumout ),
	.cout(\Add26~62 ),
	.shareout());
defparam \Add26~61 .extended_lut = "off";
defparam \Add26~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~61 .shared_arith = "off";

dffeas \A_mul_result[3] (
	.clk(clk_clk),
	.d(\Add26~61_sumout ),
	.asdata(\A_mul_partial_prod[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[3]~q ),
	.prn(vcc));
defparam \A_mul_result[3] .is_wysiwyg = "true";
defparam \A_mul_result[3] .power_up = "low";

cyclonev_lcell_comb \Add26~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[4]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[4]~q ),
	.datag(gnd),
	.cin(\Add26~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~1_sumout ),
	.cout(\Add26~2 ),
	.shareout());
defparam \Add26~1 .extended_lut = "off";
defparam \Add26~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~1 .shared_arith = "off";

dffeas \A_mul_result[4] (
	.clk(clk_clk),
	.d(\Add26~1_sumout ),
	.asdata(\A_mul_partial_prod[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[4]~q ),
	.prn(vcc));
defparam \A_mul_result[4] .is_wysiwyg = "true";
defparam \A_mul_result[4] .power_up = "low";

cyclonev_lcell_comb \Add26~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[5]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[5]~q ),
	.datag(gnd),
	.cin(\Add26~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~13_sumout ),
	.cout(\Add26~14 ),
	.shareout());
defparam \Add26~13 .extended_lut = "off";
defparam \Add26~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~13 .shared_arith = "off";

dffeas \A_mul_result[5] (
	.clk(clk_clk),
	.d(\Add26~13_sumout ),
	.asdata(\A_mul_partial_prod[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[5]~q ),
	.prn(vcc));
defparam \A_mul_result[5] .is_wysiwyg = "true";
defparam \A_mul_result[5] .power_up = "low";

cyclonev_lcell_comb \Add26~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[6]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[6]~q ),
	.datag(gnd),
	.cin(\Add26~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~41_sumout ),
	.cout(\Add26~42 ),
	.shareout());
defparam \Add26~41 .extended_lut = "off";
defparam \Add26~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~41 .shared_arith = "off";

dffeas \A_mul_result[6] (
	.clk(clk_clk),
	.d(\Add26~41_sumout ),
	.asdata(\A_mul_partial_prod[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[6]~q ),
	.prn(vcc));
defparam \A_mul_result[6] .is_wysiwyg = "true";
defparam \A_mul_result[6] .power_up = "low";

cyclonev_lcell_comb \Add26~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[7]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[7]~q ),
	.datag(gnd),
	.cin(\Add26~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~37_sumout ),
	.cout(\Add26~38 ),
	.shareout());
defparam \Add26~37 .extended_lut = "off";
defparam \Add26~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~37 .shared_arith = "off";

dffeas \A_mul_result[7] (
	.clk(clk_clk),
	.d(\Add26~37_sumout ),
	.asdata(\A_mul_partial_prod[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[7]~q ),
	.prn(vcc));
defparam \A_mul_result[7] .is_wysiwyg = "true";
defparam \A_mul_result[7] .power_up = "low";

cyclonev_lcell_comb \Add26~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[8]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[8]~q ),
	.datag(gnd),
	.cin(\Add26~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~33_sumout ),
	.cout(\Add26~34 ),
	.shareout());
defparam \Add26~33 .extended_lut = "off";
defparam \Add26~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~33 .shared_arith = "off";

dffeas \A_mul_result[8] (
	.clk(clk_clk),
	.d(\Add26~33_sumout ),
	.asdata(\A_mul_partial_prod[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[8]~q ),
	.prn(vcc));
defparam \A_mul_result[8] .is_wysiwyg = "true";
defparam \A_mul_result[8] .power_up = "low";

cyclonev_lcell_comb \Add26~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[9]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[9]~q ),
	.datag(gnd),
	.cin(\Add26~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~29_sumout ),
	.cout(\Add26~30 ),
	.shareout());
defparam \Add26~29 .extended_lut = "off";
defparam \Add26~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~29 .shared_arith = "off";

dffeas \A_mul_result[9] (
	.clk(clk_clk),
	.d(\Add26~29_sumout ),
	.asdata(\A_mul_partial_prod[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[9]~q ),
	.prn(vcc));
defparam \A_mul_result[9] .is_wysiwyg = "true";
defparam \A_mul_result[9] .power_up = "low";

cyclonev_lcell_comb \Add26~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[10]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[10]~q ),
	.datag(gnd),
	.cin(\Add26~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~25_sumout ),
	.cout(\Add26~26 ),
	.shareout());
defparam \Add26~25 .extended_lut = "off";
defparam \Add26~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~25 .shared_arith = "off";

dffeas \A_mul_result[10] (
	.clk(clk_clk),
	.d(\Add26~25_sumout ),
	.asdata(\A_mul_partial_prod[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[10]~q ),
	.prn(vcc));
defparam \A_mul_result[10] .is_wysiwyg = "true";
defparam \A_mul_result[10] .power_up = "low";

cyclonev_lcell_comb \Add26~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[11]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[11]~q ),
	.datag(gnd),
	.cin(\Add26~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~21_sumout ),
	.cout(\Add26~22 ),
	.shareout());
defparam \Add26~21 .extended_lut = "off";
defparam \Add26~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~21 .shared_arith = "off";

dffeas \A_mul_result[11] (
	.clk(clk_clk),
	.d(\Add26~21_sumout ),
	.asdata(\A_mul_partial_prod[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[11]~q ),
	.prn(vcc));
defparam \A_mul_result[11] .is_wysiwyg = "true";
defparam \A_mul_result[11] .power_up = "low";

cyclonev_lcell_comb \Add26~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[12]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[12]~q ),
	.datag(gnd),
	.cin(\Add26~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~17_sumout ),
	.cout(\Add26~18 ),
	.shareout());
defparam \Add26~17 .extended_lut = "off";
defparam \Add26~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~17 .shared_arith = "off";

dffeas \A_mul_result[12] (
	.clk(clk_clk),
	.d(\Add26~17_sumout ),
	.asdata(\A_mul_partial_prod[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[12]~q ),
	.prn(vcc));
defparam \A_mul_result[12] .is_wysiwyg = "true";
defparam \A_mul_result[12] .power_up = "low";

cyclonev_lcell_comb \Add26~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[13]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[13]~q ),
	.datag(gnd),
	.cin(\Add26~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~57_sumout ),
	.cout(\Add26~58 ),
	.shareout());
defparam \Add26~57 .extended_lut = "off";
defparam \Add26~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~57 .shared_arith = "off";

dffeas \A_mul_result[13] (
	.clk(clk_clk),
	.d(\Add26~57_sumout ),
	.asdata(\A_mul_partial_prod[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[13]~q ),
	.prn(vcc));
defparam \A_mul_result[13] .is_wysiwyg = "true";
defparam \A_mul_result[13] .power_up = "low";

cyclonev_lcell_comb \Add26~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[14]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[14]~q ),
	.datag(gnd),
	.cin(\Add26~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~53_sumout ),
	.cout(\Add26~54 ),
	.shareout());
defparam \Add26~53 .extended_lut = "off";
defparam \Add26~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~53 .shared_arith = "off";

dffeas \A_mul_result[14] (
	.clk(clk_clk),
	.d(\Add26~53_sumout ),
	.asdata(\A_mul_partial_prod[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[14]~q ),
	.prn(vcc));
defparam \A_mul_result[14] .is_wysiwyg = "true";
defparam \A_mul_result[14] .power_up = "low";

dffeas \A_mul_result[15] (
	.clk(clk_clk),
	.d(\Add26~49_sumout ),
	.asdata(\A_mul_partial_prod[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[15]~q ),
	.prn(vcc));
defparam \A_mul_result[15] .is_wysiwyg = "true";
defparam \A_mul_result[15] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~12 (
	.dataa(!\M_rot_prestep2[15]~q ),
	.datab(!\M_rot_prestep2[7]~q ),
	.datac(!\M_rot_prestep2[31]~q ),
	.datad(!\M_rot_prestep2[23]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~12 .extended_lut = "off";
defparam \M_rot[7]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~12 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~12 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[7]~q ),
	.datae(!\M_rot[7]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~12 .extended_lut = "off";
defparam \A_shift_rot_result~12 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~12 .shared_arith = "off";

dffeas \A_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[15] .is_wysiwyg = "true";
defparam \A_shift_rot_result[15] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[15]~12 (
	.dataa(!\d_readdata_d1[15]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\A_div_quot[15]~q ),
	.datad(!\A_slow_ld_data_fill_bit~0_combout ),
	.datae(!\A_slow_inst_result[15]~0_combout ),
	.dataf(!\A_slow_inst_result[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[15]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[15]~12 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[15]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[15]~12 .shared_arith = "off";

dffeas \A_slow_inst_result[15] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[15]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[15]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[15] .is_wysiwyg = "true";
defparam \A_slow_inst_result[15] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~29 (
	.dataa(!\A_inst_result[15]~q ),
	.datab(!\A_inst_result[31]~q ),
	.datac(!\A_slow_inst_result[15]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[8]~10_combout ),
	.dataf(!\A_wr_data_unfiltered[8]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~29 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[15]~29 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~30 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[15]~q ),
	.datad(!\A_shift_rot_result[15]~q ),
	.datae(!\A_wr_data_unfiltered[15]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~30 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[15]~30 .shared_arith = "off";

dffeas \W_wr_data[15] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[15]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[15]~q ),
	.prn(vcc));
defparam \W_wr_data[15] .is_wysiwyg = "true";
defparam \W_wr_data[15] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[15]~25 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[29]~4_combout ),
	.datad(!\A_mul_result[15]~q ),
	.datae(!\A_shift_rot_result[15]~q ),
	.dataf(!\A_wr_data_unfiltered[15]~29_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~25 .extended_lut = "off";
defparam \D_src2_reg[15]~25 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[15]~25 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[15]~96 (
	.dataa(!\M_alu_result[15]~q ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[29]~3_combout ),
	.datad(!\D_src2_reg[3]~13_combout ),
	.datae(!\W_wr_data[15]~q ),
	.dataf(!\D_src2_reg[15]~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~96 .extended_lut = "off";
defparam \D_src2_reg[15]~96 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[15]~96 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[15]~6 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[15]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[15]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[15]~6 .extended_lut = "off";
defparam \E_logic_result[15]~6 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[15]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15]~12 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[15]~6_combout ),
	.datad(!\E_extra_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15]~12 .extended_lut = "off";
defparam \E_alu_result[15]~12 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[15]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[15]~107 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\D_src2_reg[15]~96_combout ),
	.datae(!\D_src2_reg[29]~2_combout ),
	.dataf(!\E_alu_result[15]~12_combout ),
	.datag(!\Add24~53_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~107_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~107 .extended_lut = "on";
defparam \D_src2_reg[15]~107 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[15]~107 .shared_arith = "off";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_src2_reg[15]~107_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[15] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~53_sumout ),
	.datac(!\E_alu_result[15]~12_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15] .extended_lut = "off";
defparam \E_alu_result[15] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[15] .shared_arith = "off";

dffeas \M_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[15]~q ),
	.prn(vcc));
defparam \M_alu_result[15] .is_wysiwyg = "true";
defparam \M_alu_result[15] .power_up = "low";

cyclonev_lcell_comb \M_dc_want_fill~0 (
	.dataa(!\M_alu_result[16]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_want_fill~0 .extended_lut = "off";
defparam \M_dc_want_fill~0 .lut_mask = 64'h6666666666666666;
defparam \M_dc_want_fill~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ld_st_cache~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\Add24~37_sumout ),
	.datad(!\M_ctrl_ld_st_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_cache~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_cache~0 .extended_lut = "off";
defparam \E_ld_st_cache~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \E_ld_st_cache~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_non_bypass(
	.clk(clk_clk),
	.d(\E_ld_st_cache~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_non_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_non_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_st_non_bypass.power_up = "low";

cyclonev_lcell_comb \M_dc_want_fill~1 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_ld_st_non_bypass~q ),
	.datac(!\M_sel_data_master~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_want_fill~1 .extended_lut = "off";
defparam \M_dc_want_fill~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_want_fill~1 .shared_arith = "off";

cyclonev_lcell_comb M_dc_want_fill(
	.dataa(!\M_alu_result[15]~q ),
	.datab(!\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\M_dc_hit~0_combout ),
	.datad(!\M_dc_hit~1_combout ),
	.datae(!\M_dc_want_fill~0_combout ),
	.dataf(!\M_dc_want_fill~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_want_fill.extended_lut = "off";
defparam M_dc_want_fill.lut_mask = 64'hFFF6FFFFFFFFFFFF;
defparam M_dc_want_fill.shared_arith = "off";

dffeas A_dc_want_fill(
	.clk(clk_clk),
	.d(\M_dc_want_fill~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_want_fill~q ),
	.prn(vcc));
defparam A_dc_want_fill.is_wysiwyg = "true";
defparam A_dc_want_fill.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_sel_nxt~0 (
	.dataa(!\A_ctrl_div~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_ctrl_ld_bypass~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_sel_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_sel_nxt~0 .extended_lut = "off";
defparam \A_slow_inst_sel_nxt~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_slow_inst_sel_nxt~0 .shared_arith = "off";

dffeas A_slow_inst_sel(
	.clk(clk_clk),
	.d(\A_slow_inst_sel_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_slow_inst_sel~q ),
	.prn(vcc));
defparam A_slow_inst_sel.is_wysiwyg = "true";
defparam A_slow_inst_sel.power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~26 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_ld_align_byte2_byte3_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~26 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~26 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \A_wr_data_unfiltered[22]~26 .shared_arith = "off";

dffeas \A_mul_partial_prod[31] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_mult_cell|Add0~61_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[31]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[31] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[31] .power_up = "low";

cyclonev_lcell_comb \Add26~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[31]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[31]~q ),
	.datag(gnd),
	.cin(\Add26~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add26~125_sumout ),
	.cout(),
	.shareout());
defparam \Add26~125 .extended_lut = "off";
defparam \Add26~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add26~125 .shared_arith = "off";

dffeas \A_mul_result[31] (
	.clk(clk_clk),
	.d(\Add26~125_sumout ),
	.asdata(\A_mul_partial_prod[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[31]~q ),
	.prn(vcc));
defparam \A_mul_result[31] .is_wysiwyg = "true";
defparam \A_mul_result[31] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~31 (
	.dataa(!\M_rot_prestep2[31]~q ),
	.datab(!\M_rot_prestep2[23]~q ),
	.datac(!\M_rot_prestep2[15]~q ),
	.datad(!\M_rot_prestep2[7]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~31 .extended_lut = "off";
defparam \M_rot[7]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~31 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~31 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[7]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~31 .extended_lut = "off";
defparam \A_shift_rot_result~31 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~31 .shared_arith = "off";

dffeas \A_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[31] .is_wysiwyg = "true";
defparam \A_shift_rot_result[31] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[31]~31 (
	.dataa(!\A_ld_align_byte2_byte3_fill~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[31]~31 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[31]~31 .lut_mask = 64'h2727272727272727;
defparam \A_slow_inst_result_nxt[31]~31 .shared_arith = "off";

cyclonev_lcell_comb \Add14~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_quot[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~125_sumout ),
	.cout(),
	.shareout());
defparam \Add14~125 .extended_lut = "off";
defparam \Add14~125 .lut_mask = 64'h00000000000000FF;
defparam \Add14~125 .shared_arith = "off";

dffeas \A_div_quot[31] (
	.clk(clk_clk),
	.d(\Add14~125_sumout ),
	.asdata(\M_div_negate_result~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_quot_en~combout ),
	.q(\A_div_quot[31]~q ),
	.prn(vcc));
defparam \A_div_quot[31] .is_wysiwyg = "true";
defparam \A_div_quot[31] .power_up = "low";

dffeas \A_slow_inst_result[31] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[31]~31_combout ),
	.asdata(\A_div_quot[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_div~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[31]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[31] .is_wysiwyg = "true";
defparam \A_slow_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[31]~67 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_data_ram_ld_align_sign_bit~q ),
	.datad(!\A_ctrl_ld_signed~q ),
	.datae(!\A_shift_rot_result[31]~q ),
	.dataf(!\A_slow_inst_result[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[31]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[31]~67 .extended_lut = "off";
defparam \A_wr_data_unfiltered[31]~67 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[31]~67 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[31]~68 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[31]~q ),
	.datac(!\A_wr_data_unfiltered[22]~26_combout ),
	.datad(!\A_mul_result[31]~q ),
	.datae(!\A_wr_data_unfiltered[31]~67_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[31]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[31]~68 .extended_lut = "off";
defparam \A_wr_data_unfiltered[31]~68 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[31]~68 .shared_arith = "off";

dffeas \W_wr_data[31] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[31]~68_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[31]~q ),
	.prn(vcc));
defparam \W_wr_data[31] .is_wysiwyg = "true";
defparam \W_wr_data[31] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[31]~31 (
	.dataa(!\M_alu_result[31]~q ),
	.datab(!\A_wr_data_unfiltered[31]~68_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\E_src1[3]~0_combout ),
	.dataf(!\E_src1[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[31]~31 .extended_lut = "off";
defparam \D_src1_reg[31]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[31]~31 .shared_arith = "off";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\D_src1_reg[31]~31_combout ),
	.asdata(\E_alu_result[31]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal298~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

cyclonev_lcell_comb \Add24~37 (
	.dataa(!\E_ctrl_alu_signed_comparison~q ),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(\Add24~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~37_sumout ),
	.cout(\Add24~38 ),
	.shareout());
defparam \Add24~37 .extended_lut = "off";
defparam \Add24~37 .lut_mask = 64'h000055AA00009966;
defparam \Add24~37 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~60 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~37_sumout ),
	.datac(!\D_src2_reg[0]~31_combout ),
	.datad(!\E_alu_result~31_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~60 .extended_lut = "off";
defparam \D_src2_reg[31]~60 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[31]~60 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~61 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\D_src2_reg[3]~13_combout ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\A_wr_data_unfiltered[31]~68_combout ),
	.dataf(!\M_alu_result[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~61 .extended_lut = "off";
defparam \D_src2_reg[31]~61 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[31]~61 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~28 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~28 .extended_lut = "off";
defparam \D_src2[31]~28 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_src2[31]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~29 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~30_combout ),
	.datac(!\D_src2_reg[31]~60_combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\D_src2_reg[31]~61_combout ),
	.dataf(!\D_src2[31]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~29 .extended_lut = "off";
defparam \D_src2[31]~29 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[31]~29 .shared_arith = "off";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\D_src2[31]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclonev_lcell_comb \Add24~65 (
	.dataa(gnd),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~65_sumout ),
	.cout(),
	.shareout());
defparam \Add24~65 .extended_lut = "off";
defparam \Add24~65 .lut_mask = 64'h0000000000003333;
defparam \Add24~65 .shared_arith = "off";

cyclonev_lcell_comb \E_br_result~2 (
	.dataa(!\Add24~65_sumout ),
	.datab(!\E_br_result~0_combout ),
	.datac(!\E_br_result~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~2 .extended_lut = "off";
defparam \E_br_result~2 .lut_mask = 64'h2727272727272727;
defparam \E_br_result~2 .shared_arith = "off";

dffeas E_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_br_cond~q ),
	.prn(vcc));
defparam E_ctrl_br_cond.is_wysiwyg = "true";
defparam E_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~0 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~0 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_flush_pipe_always~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~1 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\D_ctrl_flush_pipe_always~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~1 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~1 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_flush_pipe_always~1 .shared_arith = "off";

dffeas E_ctrl_flush_pipe_always(
	.clk(clk_clk),
	.d(\D_ctrl_flush_pipe_always~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_flush_pipe_always~q ),
	.prn(vcc));
defparam E_ctrl_flush_pipe_always.is_wysiwyg = "true";
defparam E_ctrl_flush_pipe_always.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_nxt~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_bht_data[1]~q ),
	.datad(!\E_br_result~2_combout ),
	.datae(!\E_ctrl_br_cond~q ),
	.dataf(!\E_ctrl_flush_pipe_always~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_nxt~0 .extended_lut = "off";
defparam \M_pipe_flush_nxt~0 .lut_mask = 64'hFFFFFFFFFFFFEFFE;
defparam \M_pipe_flush_nxt~0 .shared_arith = "off";

dffeas M_pipe_flush(
	.clk(clk_clk),
	.d(\M_pipe_flush_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush~q ),
	.prn(vcc));
defparam M_pipe_flush.is_wysiwyg = "true";
defparam M_pipe_flush.power_up = "low";

dffeas E_wr_dst_reg_from_D(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_wr_dst_reg_from_D~q ),
	.prn(vcc));
defparam E_wr_dst_reg_from_D.is_wysiwyg = "true";
defparam E_wr_dst_reg_from_D.power_up = "low";

cyclonev_lcell_comb \E_wr_dst_reg~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_wr_dst_reg_from_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wr_dst_reg~0 .extended_lut = "off";
defparam \E_wr_dst_reg~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~0 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\E_dst_regnum[0]~q ),
	.datad(!\E_dst_regnum[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~1 (
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(!\E_dst_regnum[3]~q ),
	.datad(!\E_dst_regnum[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_b_cmp_F(
	.dataa(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\E_dst_regnum[2]~q ),
	.datac(!\E_wr_dst_reg~0_combout ),
	.datad(!\E_regnum_b_cmp_F~0_combout ),
	.datae(!\E_regnum_b_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_b_cmp_F.extended_lut = "off";
defparam E_regnum_b_cmp_F.lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam E_regnum_b_cmp_F.shared_arith = "off";

dffeas M_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_b_cmp_F~combout ),
	.asdata(\E_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\M_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_b_cmp_D.is_wysiwyg = "true";
defparam M_regnum_b_cmp_D.power_up = "low";

cyclonev_lcell_comb \D_src2_reg[29]~0 (
	.dataa(!\M_regnum_b_cmp_D~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\W_regnum_b_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~0 .extended_lut = "off";
defparam \D_src2_reg[29]~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_src2_reg[29]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~1 .extended_lut = "off";
defparam \D_src2_reg[29]~1 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \D_src2_reg[29]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~7 (
	.dataa(!\D_src2_reg[29]~3_combout ),
	.datab(!\D_src2_reg[29]~4_combout ),
	.datac(!\W_wr_data[0]~q ),
	.datad(!\A_wr_data_unfiltered[0]~5_combout ),
	.datae(!\M_alu_result[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~7 .extended_lut = "off";
defparam \D_src2_reg[0]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[0]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~8 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\E_alu_result[0]~combout ),
	.datad(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\D_src2_reg[0]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~8 .extended_lut = "off";
defparam \D_src2_reg[0]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[0]~8 .shared_arith = "off";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(\D_src2_reg[0]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[0]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

cyclonev_lcell_comb \Add9~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~17_sumout ),
	.cout(\Add9~18 ),
	.shareout());
defparam \Add9~17 .extended_lut = "off";
defparam \Add9~17 .lut_mask = 64'h000000000000FF00;
defparam \Add9~17 .shared_arith = "off";

dffeas \M_div_src2[0] (
	.clk(clk_clk),
	.d(\Add9~17_sumout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[0]~q ),
	.prn(vcc));
defparam \M_div_src2[0] .is_wysiwyg = "true";
defparam \M_div_src2[0] .power_up = "low";

cyclonev_lcell_comb \A_div_den[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_div_den[0]~q ),
	.datac(!\Add11~1_sumout ),
	.datad(!\A_div_discover_quotient_bits~0_combout ),
	.datae(!\M_div_src2[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_den[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_den[0]~0 .extended_lut = "off";
defparam \A_div_den[0]~0 .lut_mask = 64'hBF1FFFFFBF1FFFFF;
defparam \A_div_den[0]~0 .shared_arith = "off";

dffeas \A_div_den[0] (
	.clk(clk_clk),
	.d(\A_div_den[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_den[0]~q ),
	.prn(vcc));
defparam \A_div_den[0] .is_wysiwyg = "true";
defparam \A_div_den[0] .power_up = "low";

cyclonev_lcell_comb \Add9~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~21_sumout ),
	.cout(\Add9~22 ),
	.shareout());
defparam \Add9~21 .extended_lut = "off";
defparam \Add9~21 .lut_mask = 64'h000000000000FF00;
defparam \Add9~21 .shared_arith = "off";

dffeas \M_div_src2[1] (
	.clk(clk_clk),
	.d(\Add9~21_sumout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[1]~q ),
	.prn(vcc));
defparam \M_div_src2[1] .is_wysiwyg = "true";
defparam \M_div_src2[1] .power_up = "low";

cyclonev_lcell_comb A_div_den_en(
	.dataa(!\A_stall~combout ),
	.datab(!\Add11~1_sumout ),
	.datac(!\A_div_discover_quotient_bits~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_den_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_div_den_en.extended_lut = "off";
defparam A_div_den_en.lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam A_div_den_en.shared_arith = "off";

dffeas \A_div_den[1] (
	.clk(clk_clk),
	.d(\A_div_den[0]~q ),
	.asdata(\M_div_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[1]~q ),
	.prn(vcc));
defparam \A_div_den[1] .is_wysiwyg = "true";
defparam \A_div_den[1] .power_up = "low";

cyclonev_lcell_comb \Add9~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~25_sumout ),
	.cout(\Add9~26 ),
	.shareout());
defparam \Add9~25 .extended_lut = "off";
defparam \Add9~25 .lut_mask = 64'h000000000000FF00;
defparam \Add9~25 .shared_arith = "off";

dffeas \M_div_src2[2] (
	.clk(clk_clk),
	.d(\Add9~25_sumout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[2]~q ),
	.prn(vcc));
defparam \M_div_src2[2] .is_wysiwyg = "true";
defparam \M_div_src2[2] .power_up = "low";

dffeas \A_div_den[2] (
	.clk(clk_clk),
	.d(\A_div_den[1]~q ),
	.asdata(\M_div_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[2]~q ),
	.prn(vcc));
defparam \A_div_den[2] .is_wysiwyg = "true";
defparam \A_div_den[2] .power_up = "low";

cyclonev_lcell_comb \Add9~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~29_sumout ),
	.cout(\Add9~30 ),
	.shareout());
defparam \Add9~29 .extended_lut = "off";
defparam \Add9~29 .lut_mask = 64'h000000000000FF00;
defparam \Add9~29 .shared_arith = "off";

dffeas \M_div_src2[3] (
	.clk(clk_clk),
	.d(\Add9~29_sumout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[3]~q ),
	.prn(vcc));
defparam \M_div_src2[3] .is_wysiwyg = "true";
defparam \M_div_src2[3] .power_up = "low";

dffeas \A_div_den[3] (
	.clk(clk_clk),
	.d(\A_div_den[2]~q ),
	.asdata(\M_div_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[3]~q ),
	.prn(vcc));
defparam \A_div_den[3] .is_wysiwyg = "true";
defparam \A_div_den[3] .power_up = "low";

cyclonev_lcell_comb \Add9~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~33_sumout ),
	.cout(\Add9~34 ),
	.shareout());
defparam \Add9~33 .extended_lut = "off";
defparam \Add9~33 .lut_mask = 64'h000000000000FF00;
defparam \Add9~33 .shared_arith = "off";

dffeas \M_div_src2[4] (
	.clk(clk_clk),
	.d(\Add9~33_sumout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[4]~q ),
	.prn(vcc));
defparam \M_div_src2[4] .is_wysiwyg = "true";
defparam \M_div_src2[4] .power_up = "low";

dffeas \A_div_den[4] (
	.clk(clk_clk),
	.d(\A_div_den[3]~q ),
	.asdata(\M_div_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[4]~q ),
	.prn(vcc));
defparam \A_div_den[4] .is_wysiwyg = "true";
defparam \A_div_den[4] .power_up = "low";

cyclonev_lcell_comb \Add9~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~37_sumout ),
	.cout(\Add9~38 ),
	.shareout());
defparam \Add9~37 .extended_lut = "off";
defparam \Add9~37 .lut_mask = 64'h000000000000FF00;
defparam \Add9~37 .shared_arith = "off";

dffeas \M_div_src2[5] (
	.clk(clk_clk),
	.d(\Add9~37_sumout ),
	.asdata(\E_src2[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[5]~q ),
	.prn(vcc));
defparam \M_div_src2[5] .is_wysiwyg = "true";
defparam \M_div_src2[5] .power_up = "low";

dffeas \A_div_den[5] (
	.clk(clk_clk),
	.d(\A_div_den[4]~q ),
	.asdata(\M_div_src2[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[5]~q ),
	.prn(vcc));
defparam \A_div_den[5] .is_wysiwyg = "true";
defparam \A_div_den[5] .power_up = "low";

cyclonev_lcell_comb \Add9~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~41_sumout ),
	.cout(\Add9~42 ),
	.shareout());
defparam \Add9~41 .extended_lut = "off";
defparam \Add9~41 .lut_mask = 64'h000000000000FF00;
defparam \Add9~41 .shared_arith = "off";

dffeas \M_div_src2[6] (
	.clk(clk_clk),
	.d(\Add9~41_sumout ),
	.asdata(\E_src2[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[6]~q ),
	.prn(vcc));
defparam \M_div_src2[6] .is_wysiwyg = "true";
defparam \M_div_src2[6] .power_up = "low";

dffeas \A_div_den[6] (
	.clk(clk_clk),
	.d(\A_div_den[5]~q ),
	.asdata(\M_div_src2[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[6]~q ),
	.prn(vcc));
defparam \A_div_den[6] .is_wysiwyg = "true";
defparam \A_div_den[6] .power_up = "low";

cyclonev_lcell_comb \Add9~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~45_sumout ),
	.cout(\Add9~46 ),
	.shareout());
defparam \Add9~45 .extended_lut = "off";
defparam \Add9~45 .lut_mask = 64'h000000000000FF00;
defparam \Add9~45 .shared_arith = "off";

dffeas \M_div_src2[7] (
	.clk(clk_clk),
	.d(\Add9~45_sumout ),
	.asdata(\E_src2[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[7]~q ),
	.prn(vcc));
defparam \M_div_src2[7] .is_wysiwyg = "true";
defparam \M_div_src2[7] .power_up = "low";

dffeas \A_div_den[7] (
	.clk(clk_clk),
	.d(\A_div_den[6]~q ),
	.asdata(\M_div_src2[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[7]~q ),
	.prn(vcc));
defparam \A_div_den[7] .is_wysiwyg = "true";
defparam \A_div_den[7] .power_up = "low";

cyclonev_lcell_comb \Add9~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~49_sumout ),
	.cout(\Add9~50 ),
	.shareout());
defparam \Add9~49 .extended_lut = "off";
defparam \Add9~49 .lut_mask = 64'h000000000000FF00;
defparam \Add9~49 .shared_arith = "off";

dffeas \M_div_src2[8] (
	.clk(clk_clk),
	.d(\Add9~49_sumout ),
	.asdata(\E_src2[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[8]~q ),
	.prn(vcc));
defparam \M_div_src2[8] .is_wysiwyg = "true";
defparam \M_div_src2[8] .power_up = "low";

dffeas \A_div_den[8] (
	.clk(clk_clk),
	.d(\A_div_den[7]~q ),
	.asdata(\M_div_src2[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[8]~q ),
	.prn(vcc));
defparam \A_div_den[8] .is_wysiwyg = "true";
defparam \A_div_den[8] .power_up = "low";

cyclonev_lcell_comb \Add9~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~53_sumout ),
	.cout(\Add9~54 ),
	.shareout());
defparam \Add9~53 .extended_lut = "off";
defparam \Add9~53 .lut_mask = 64'h000000000000FF00;
defparam \Add9~53 .shared_arith = "off";

dffeas \M_div_src2[9] (
	.clk(clk_clk),
	.d(\Add9~53_sumout ),
	.asdata(\E_src2[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[9]~q ),
	.prn(vcc));
defparam \M_div_src2[9] .is_wysiwyg = "true";
defparam \M_div_src2[9] .power_up = "low";

dffeas \A_div_den[9] (
	.clk(clk_clk),
	.d(\A_div_den[8]~q ),
	.asdata(\M_div_src2[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[9]~q ),
	.prn(vcc));
defparam \A_div_den[9] .is_wysiwyg = "true";
defparam \A_div_den[9] .power_up = "low";

cyclonev_lcell_comb \Add9~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~57_sumout ),
	.cout(\Add9~58 ),
	.shareout());
defparam \Add9~57 .extended_lut = "off";
defparam \Add9~57 .lut_mask = 64'h000000000000FF00;
defparam \Add9~57 .shared_arith = "off";

dffeas \M_div_src2[10] (
	.clk(clk_clk),
	.d(\Add9~57_sumout ),
	.asdata(\E_src2[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[10]~q ),
	.prn(vcc));
defparam \M_div_src2[10] .is_wysiwyg = "true";
defparam \M_div_src2[10] .power_up = "low";

dffeas \A_div_den[10] (
	.clk(clk_clk),
	.d(\A_div_den[9]~q ),
	.asdata(\M_div_src2[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[10]~q ),
	.prn(vcc));
defparam \A_div_den[10] .is_wysiwyg = "true";
defparam \A_div_den[10] .power_up = "low";

cyclonev_lcell_comb \Add9~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~61_sumout ),
	.cout(\Add9~62 ),
	.shareout());
defparam \Add9~61 .extended_lut = "off";
defparam \Add9~61 .lut_mask = 64'h000000000000FF00;
defparam \Add9~61 .shared_arith = "off";

dffeas \M_div_src2[11] (
	.clk(clk_clk),
	.d(\Add9~61_sumout ),
	.asdata(\E_src2[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[11]~q ),
	.prn(vcc));
defparam \M_div_src2[11] .is_wysiwyg = "true";
defparam \M_div_src2[11] .power_up = "low";

dffeas \A_div_den[11] (
	.clk(clk_clk),
	.d(\A_div_den[10]~q ),
	.asdata(\M_div_src2[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[11]~q ),
	.prn(vcc));
defparam \A_div_den[11] .is_wysiwyg = "true";
defparam \A_div_den[11] .power_up = "low";

cyclonev_lcell_comb \Add9~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~65_sumout ),
	.cout(\Add9~66 ),
	.shareout());
defparam \Add9~65 .extended_lut = "off";
defparam \Add9~65 .lut_mask = 64'h000000000000FF00;
defparam \Add9~65 .shared_arith = "off";

dffeas \M_div_src2[12] (
	.clk(clk_clk),
	.d(\Add9~65_sumout ),
	.asdata(\E_src2[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[12]~q ),
	.prn(vcc));
defparam \M_div_src2[12] .is_wysiwyg = "true";
defparam \M_div_src2[12] .power_up = "low";

dffeas \A_div_den[12] (
	.clk(clk_clk),
	.d(\A_div_den[11]~q ),
	.asdata(\M_div_src2[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[12]~q ),
	.prn(vcc));
defparam \A_div_den[12] .is_wysiwyg = "true";
defparam \A_div_den[12] .power_up = "low";

cyclonev_lcell_comb \Add9~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~69_sumout ),
	.cout(\Add9~70 ),
	.shareout());
defparam \Add9~69 .extended_lut = "off";
defparam \Add9~69 .lut_mask = 64'h000000000000FF00;
defparam \Add9~69 .shared_arith = "off";

dffeas \M_div_src2[13] (
	.clk(clk_clk),
	.d(\Add9~69_sumout ),
	.asdata(\E_src2[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[13]~q ),
	.prn(vcc));
defparam \M_div_src2[13] .is_wysiwyg = "true";
defparam \M_div_src2[13] .power_up = "low";

dffeas \A_div_den[13] (
	.clk(clk_clk),
	.d(\A_div_den[12]~q ),
	.asdata(\M_div_src2[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[13]~q ),
	.prn(vcc));
defparam \A_div_den[13] .is_wysiwyg = "true";
defparam \A_div_den[13] .power_up = "low";

cyclonev_lcell_comb \Add9~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~73_sumout ),
	.cout(\Add9~74 ),
	.shareout());
defparam \Add9~73 .extended_lut = "off";
defparam \Add9~73 .lut_mask = 64'h000000000000FF00;
defparam \Add9~73 .shared_arith = "off";

dffeas \M_div_src2[14] (
	.clk(clk_clk),
	.d(\Add9~73_sumout ),
	.asdata(\E_src2[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[14]~q ),
	.prn(vcc));
defparam \M_div_src2[14] .is_wysiwyg = "true";
defparam \M_div_src2[14] .power_up = "low";

dffeas \A_div_den[14] (
	.clk(clk_clk),
	.d(\A_div_den[13]~q ),
	.asdata(\M_div_src2[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[14]~q ),
	.prn(vcc));
defparam \A_div_den[14] .is_wysiwyg = "true";
defparam \A_div_den[14] .power_up = "low";

cyclonev_lcell_comb \Add9~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~77_sumout ),
	.cout(\Add9~78 ),
	.shareout());
defparam \Add9~77 .extended_lut = "off";
defparam \Add9~77 .lut_mask = 64'h000000000000FF00;
defparam \Add9~77 .shared_arith = "off";

dffeas \M_div_src2[15] (
	.clk(clk_clk),
	.d(\Add9~77_sumout ),
	.asdata(\E_src2[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[15]~q ),
	.prn(vcc));
defparam \M_div_src2[15] .is_wysiwyg = "true";
defparam \M_div_src2[15] .power_up = "low";

dffeas \A_div_den[15] (
	.clk(clk_clk),
	.d(\A_div_den[14]~q ),
	.asdata(\M_div_src2[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[15]~q ),
	.prn(vcc));
defparam \A_div_den[15] .is_wysiwyg = "true";
defparam \A_div_den[15] .power_up = "low";

cyclonev_lcell_comb \Add9~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~85_sumout ),
	.cout(\Add9~86 ),
	.shareout());
defparam \Add9~85 .extended_lut = "off";
defparam \Add9~85 .lut_mask = 64'h000000000000FF00;
defparam \Add9~85 .shared_arith = "off";

dffeas \M_div_src2[16] (
	.clk(clk_clk),
	.d(\Add9~85_sumout ),
	.asdata(\E_src2[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[16]~q ),
	.prn(vcc));
defparam \M_div_src2[16] .is_wysiwyg = "true";
defparam \M_div_src2[16] .power_up = "low";

dffeas \A_div_den[16] (
	.clk(clk_clk),
	.d(\A_div_den[15]~q ),
	.asdata(\M_div_src2[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[16]~q ),
	.prn(vcc));
defparam \A_div_den[16] .is_wysiwyg = "true";
defparam \A_div_den[16] .power_up = "low";

cyclonev_lcell_comb \Add9~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~89_sumout ),
	.cout(\Add9~90 ),
	.shareout());
defparam \Add9~89 .extended_lut = "off";
defparam \Add9~89 .lut_mask = 64'h000000000000FF00;
defparam \Add9~89 .shared_arith = "off";

dffeas \M_div_src2[17] (
	.clk(clk_clk),
	.d(\Add9~89_sumout ),
	.asdata(\E_src2[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[17]~q ),
	.prn(vcc));
defparam \M_div_src2[17] .is_wysiwyg = "true";
defparam \M_div_src2[17] .power_up = "low";

dffeas \A_div_den[17] (
	.clk(clk_clk),
	.d(\A_div_den[16]~q ),
	.asdata(\M_div_src2[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[17]~q ),
	.prn(vcc));
defparam \A_div_den[17] .is_wysiwyg = "true";
defparam \A_div_den[17] .power_up = "low";

cyclonev_lcell_comb \Add9~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~93_sumout ),
	.cout(\Add9~94 ),
	.shareout());
defparam \Add9~93 .extended_lut = "off";
defparam \Add9~93 .lut_mask = 64'h000000000000FF00;
defparam \Add9~93 .shared_arith = "off";

dffeas \M_div_src2[18] (
	.clk(clk_clk),
	.d(\Add9~93_sumout ),
	.asdata(\E_src2[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[18]~q ),
	.prn(vcc));
defparam \M_div_src2[18] .is_wysiwyg = "true";
defparam \M_div_src2[18] .power_up = "low";

dffeas \A_div_den[18] (
	.clk(clk_clk),
	.d(\A_div_den[17]~q ),
	.asdata(\M_div_src2[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[18]~q ),
	.prn(vcc));
defparam \A_div_den[18] .is_wysiwyg = "true";
defparam \A_div_den[18] .power_up = "low";

cyclonev_lcell_comb \Add9~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~97_sumout ),
	.cout(\Add9~98 ),
	.shareout());
defparam \Add9~97 .extended_lut = "off";
defparam \Add9~97 .lut_mask = 64'h000000000000FF00;
defparam \Add9~97 .shared_arith = "off";

dffeas \M_div_src2[19] (
	.clk(clk_clk),
	.d(\Add9~97_sumout ),
	.asdata(\E_src2[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[19]~q ),
	.prn(vcc));
defparam \M_div_src2[19] .is_wysiwyg = "true";
defparam \M_div_src2[19] .power_up = "low";

dffeas \A_div_den[19] (
	.clk(clk_clk),
	.d(\A_div_den[18]~q ),
	.asdata(\M_div_src2[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[19]~q ),
	.prn(vcc));
defparam \A_div_den[19] .is_wysiwyg = "true";
defparam \A_div_den[19] .power_up = "low";

cyclonev_lcell_comb \Add9~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~101_sumout ),
	.cout(\Add9~102 ),
	.shareout());
defparam \Add9~101 .extended_lut = "off";
defparam \Add9~101 .lut_mask = 64'h000000000000FF00;
defparam \Add9~101 .shared_arith = "off";

dffeas \M_div_src2[20] (
	.clk(clk_clk),
	.d(\Add9~101_sumout ),
	.asdata(\E_src2[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[20]~q ),
	.prn(vcc));
defparam \M_div_src2[20] .is_wysiwyg = "true";
defparam \M_div_src2[20] .power_up = "low";

dffeas \A_div_den[20] (
	.clk(clk_clk),
	.d(\A_div_den[19]~q ),
	.asdata(\M_div_src2[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[20]~q ),
	.prn(vcc));
defparam \A_div_den[20] .is_wysiwyg = "true";
defparam \A_div_den[20] .power_up = "low";

cyclonev_lcell_comb \Add9~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~105_sumout ),
	.cout(\Add9~106 ),
	.shareout());
defparam \Add9~105 .extended_lut = "off";
defparam \Add9~105 .lut_mask = 64'h000000000000FF00;
defparam \Add9~105 .shared_arith = "off";

dffeas \M_div_src2[21] (
	.clk(clk_clk),
	.d(\Add9~105_sumout ),
	.asdata(\E_src2[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[21]~q ),
	.prn(vcc));
defparam \M_div_src2[21] .is_wysiwyg = "true";
defparam \M_div_src2[21] .power_up = "low";

dffeas \A_div_den[21] (
	.clk(clk_clk),
	.d(\A_div_den[20]~q ),
	.asdata(\M_div_src2[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[21]~q ),
	.prn(vcc));
defparam \A_div_den[21] .is_wysiwyg = "true";
defparam \A_div_den[21] .power_up = "low";

cyclonev_lcell_comb \Add9~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~109_sumout ),
	.cout(\Add9~110 ),
	.shareout());
defparam \Add9~109 .extended_lut = "off";
defparam \Add9~109 .lut_mask = 64'h000000000000FF00;
defparam \Add9~109 .shared_arith = "off";

dffeas \M_div_src2[22] (
	.clk(clk_clk),
	.d(\Add9~109_sumout ),
	.asdata(\E_src2[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[22]~q ),
	.prn(vcc));
defparam \M_div_src2[22] .is_wysiwyg = "true";
defparam \M_div_src2[22] .power_up = "low";

dffeas \A_div_den[22] (
	.clk(clk_clk),
	.d(\A_div_den[21]~q ),
	.asdata(\M_div_src2[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[22]~q ),
	.prn(vcc));
defparam \A_div_den[22] .is_wysiwyg = "true";
defparam \A_div_den[22] .power_up = "low";

cyclonev_lcell_comb \Add9~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~113_sumout ),
	.cout(\Add9~114 ),
	.shareout());
defparam \Add9~113 .extended_lut = "off";
defparam \Add9~113 .lut_mask = 64'h000000000000FF00;
defparam \Add9~113 .shared_arith = "off";

dffeas \M_div_src2[23] (
	.clk(clk_clk),
	.d(\Add9~113_sumout ),
	.asdata(\E_src2[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[23]~q ),
	.prn(vcc));
defparam \M_div_src2[23] .is_wysiwyg = "true";
defparam \M_div_src2[23] .power_up = "low";

dffeas \A_div_den[23] (
	.clk(clk_clk),
	.d(\A_div_den[22]~q ),
	.asdata(\M_div_src2[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[23]~q ),
	.prn(vcc));
defparam \A_div_den[23] .is_wysiwyg = "true";
defparam \A_div_den[23] .power_up = "low";

cyclonev_lcell_comb \Add9~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~117_sumout ),
	.cout(\Add9~118 ),
	.shareout());
defparam \Add9~117 .extended_lut = "off";
defparam \Add9~117 .lut_mask = 64'h000000000000FF00;
defparam \Add9~117 .shared_arith = "off";

dffeas \M_div_src2[24] (
	.clk(clk_clk),
	.d(\Add9~117_sumout ),
	.asdata(\E_src2[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[24]~q ),
	.prn(vcc));
defparam \M_div_src2[24] .is_wysiwyg = "true";
defparam \M_div_src2[24] .power_up = "low";

dffeas \A_div_den[24] (
	.clk(clk_clk),
	.d(\A_div_den[23]~q ),
	.asdata(\M_div_src2[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[24]~q ),
	.prn(vcc));
defparam \A_div_den[24] .is_wysiwyg = "true";
defparam \A_div_den[24] .power_up = "low";

cyclonev_lcell_comb \Add9~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~121_sumout ),
	.cout(\Add9~122 ),
	.shareout());
defparam \Add9~121 .extended_lut = "off";
defparam \Add9~121 .lut_mask = 64'h000000000000FF00;
defparam \Add9~121 .shared_arith = "off";

dffeas \M_div_src2[25] (
	.clk(clk_clk),
	.d(\Add9~121_sumout ),
	.asdata(\E_src2[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[25]~q ),
	.prn(vcc));
defparam \M_div_src2[25] .is_wysiwyg = "true";
defparam \M_div_src2[25] .power_up = "low";

dffeas \A_div_den[25] (
	.clk(clk_clk),
	.d(\A_div_den[24]~q ),
	.asdata(\M_div_src2[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[25]~q ),
	.prn(vcc));
defparam \A_div_den[25] .is_wysiwyg = "true";
defparam \A_div_den[25] .power_up = "low";

cyclonev_lcell_comb \Add9~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~125_sumout ),
	.cout(\Add9~126 ),
	.shareout());
defparam \Add9~125 .extended_lut = "off";
defparam \Add9~125 .lut_mask = 64'h000000000000FF00;
defparam \Add9~125 .shared_arith = "off";

dffeas \M_div_src2[26] (
	.clk(clk_clk),
	.d(\Add9~125_sumout ),
	.asdata(\E_src2[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[26]~q ),
	.prn(vcc));
defparam \M_div_src2[26] .is_wysiwyg = "true";
defparam \M_div_src2[26] .power_up = "low";

dffeas \A_div_den[26] (
	.clk(clk_clk),
	.d(\A_div_den[25]~q ),
	.asdata(\M_div_src2[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[26]~q ),
	.prn(vcc));
defparam \A_div_den[26] .is_wysiwyg = "true";
defparam \A_div_den[26] .power_up = "low";

cyclonev_lcell_comb \Add9~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~81_sumout ),
	.cout(\Add9~82 ),
	.shareout());
defparam \Add9~81 .extended_lut = "off";
defparam \Add9~81 .lut_mask = 64'h000000000000FF00;
defparam \Add9~81 .shared_arith = "off";

dffeas \M_div_src2[27] (
	.clk(clk_clk),
	.d(\Add9~81_sumout ),
	.asdata(\E_src2[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[27]~q ),
	.prn(vcc));
defparam \M_div_src2[27] .is_wysiwyg = "true";
defparam \M_div_src2[27] .power_up = "low";

dffeas \A_div_den[27] (
	.clk(clk_clk),
	.d(\A_div_den[26]~q ),
	.asdata(\M_div_src2[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[27]~q ),
	.prn(vcc));
defparam \A_div_den[27] .is_wysiwyg = "true";
defparam \A_div_den[27] .power_up = "low";

cyclonev_lcell_comb \Add9~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~13_sumout ),
	.cout(\Add9~14 ),
	.shareout());
defparam \Add9~13 .extended_lut = "off";
defparam \Add9~13 .lut_mask = 64'h000000000000FF00;
defparam \Add9~13 .shared_arith = "off";

dffeas \M_div_src2[28] (
	.clk(clk_clk),
	.d(\Add9~13_sumout ),
	.asdata(\E_src2[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[28]~q ),
	.prn(vcc));
defparam \M_div_src2[28] .is_wysiwyg = "true";
defparam \M_div_src2[28] .power_up = "low";

dffeas \A_div_den[28] (
	.clk(clk_clk),
	.d(\A_div_den[27]~q ),
	.asdata(\M_div_src2[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[28]~q ),
	.prn(vcc));
defparam \A_div_den[28] .is_wysiwyg = "true";
defparam \A_div_den[28] .power_up = "low";

cyclonev_lcell_comb \Add9~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~9_sumout ),
	.cout(\Add9~10 ),
	.shareout());
defparam \Add9~9 .extended_lut = "off";
defparam \Add9~9 .lut_mask = 64'h000000000000FF00;
defparam \Add9~9 .shared_arith = "off";

dffeas \M_div_src2[29] (
	.clk(clk_clk),
	.d(\Add9~9_sumout ),
	.asdata(\E_src2[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[29]~q ),
	.prn(vcc));
defparam \M_div_src2[29] .is_wysiwyg = "true";
defparam \M_div_src2[29] .power_up = "low";

dffeas \A_div_den[29] (
	.clk(clk_clk),
	.d(\A_div_den[28]~q ),
	.asdata(\M_div_src2[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[29]~q ),
	.prn(vcc));
defparam \A_div_den[29] .is_wysiwyg = "true";
defparam \A_div_den[29] .power_up = "low";

cyclonev_lcell_comb \Add9~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~5_sumout ),
	.cout(\Add9~6 ),
	.shareout());
defparam \Add9~5 .extended_lut = "off";
defparam \Add9~5 .lut_mask = 64'h000000000000FF00;
defparam \Add9~5 .shared_arith = "off";

dffeas \M_div_src2[30] (
	.clk(clk_clk),
	.d(\Add9~5_sumout ),
	.asdata(\E_src2[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[30]~q ),
	.prn(vcc));
defparam \M_div_src2[30] .is_wysiwyg = "true";
defparam \M_div_src2[30] .power_up = "low";

dffeas \A_div_den[30] (
	.clk(clk_clk),
	.d(\A_div_den[29]~q ),
	.asdata(\M_div_src2[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[30]~q ),
	.prn(vcc));
defparam \A_div_den[30] .is_wysiwyg = "true";
defparam \A_div_den[30] .power_up = "low";

cyclonev_lcell_comb \Add9~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~1_sumout ),
	.cout(),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h000000000000FF00;
defparam \Add9~1 .shared_arith = "off";

dffeas \M_div_src2[31] (
	.clk(clk_clk),
	.d(\Add9~1_sumout ),
	.asdata(\E_src2[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src2~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src2[31]~q ),
	.prn(vcc));
defparam \M_div_src2[31] .is_wysiwyg = "true";
defparam \M_div_src2[31] .power_up = "low";

dffeas \A_div_den[31] (
	.clk(clk_clk),
	.d(\A_div_den[30]~q ),
	.asdata(\M_div_src2[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_den_en~combout ),
	.q(\A_div_den[31]~q ),
	.prn(vcc));
defparam \A_div_den[31] .is_wysiwyg = "true";
defparam \A_div_den[31] .power_up = "low";

cyclonev_lcell_comb \Add8~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~9_sumout ),
	.cout(\Add8~10 ),
	.shareout());
defparam \Add8~9 .extended_lut = "off";
defparam \Add8~9 .lut_mask = 64'h000000000000FF00;
defparam \Add8~9 .shared_arith = "off";

dffeas \M_div_src1[0] (
	.clk(clk_clk),
	.d(\Add8~9_sumout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[0]~q ),
	.prn(vcc));
defparam \M_div_src1[0] .is_wysiwyg = "true";
defparam \M_div_src1[0] .power_up = "low";

cyclonev_lcell_comb \A_div_rem[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_div_rem[0]~q ),
	.datac(!\Add11~1_sumout ),
	.datad(!\A_div_discover_quotient_bits~0_combout ),
	.datae(!\M_div_src1[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_rem[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_rem[0]~0 .extended_lut = "off";
defparam \A_div_rem[0]~0 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \A_div_rem[0]~0 .shared_arith = "off";

dffeas \A_div_rem[0] (
	.clk(clk_clk),
	.d(\A_div_rem[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_rem[0]~q ),
	.prn(vcc));
defparam \A_div_rem[0] .is_wysiwyg = "true";
defparam \A_div_rem[0] .power_up = "low";

cyclonev_lcell_comb \Add11~134 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add11~134_cout ),
	.shareout());
defparam \Add11~134 .extended_lut = "off";
defparam \Add11~134 .lut_mask = 64'h0000000000005555;
defparam \Add11~134 .shared_arith = "off";

cyclonev_lcell_comb \Add11~129 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[0]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[0]~q ),
	.datag(gnd),
	.cin(\Add11~134_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~129_sumout ),
	.cout(\Add11~130 ),
	.shareout());
defparam \Add11~129 .extended_lut = "off";
defparam \Add11~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~129 .shared_arith = "off";

cyclonev_lcell_comb \Add8~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~13_sumout ),
	.cout(\Add8~14 ),
	.shareout());
defparam \Add8~13 .extended_lut = "off";
defparam \Add8~13 .lut_mask = 64'h000000000000FF00;
defparam \Add8~13 .shared_arith = "off";

dffeas \M_div_src1[1] (
	.clk(clk_clk),
	.d(\Add8~13_sumout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[1]~q ),
	.prn(vcc));
defparam \M_div_src1[1] .is_wysiwyg = "true";
defparam \M_div_src1[1] .power_up = "low";

cyclonev_lcell_comb A_div_rem_en(
	.dataa(!\A_stall~combout ),
	.datab(!\Add11~1_sumout ),
	.datac(!\A_div_discover_quotient_bits~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_rem_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_div_rem_en.extended_lut = "off";
defparam A_div_rem_en.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam A_div_rem_en.shared_arith = "off";

dffeas \A_div_rem[1] (
	.clk(clk_clk),
	.d(\Add11~129_sumout ),
	.asdata(\M_div_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[1]~q ),
	.prn(vcc));
defparam \A_div_rem[1] .is_wysiwyg = "true";
defparam \A_div_rem[1] .power_up = "low";

cyclonev_lcell_comb \Add11~125 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[1]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[1]~q ),
	.datag(gnd),
	.cin(\Add11~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~125_sumout ),
	.cout(\Add11~126 ),
	.shareout());
defparam \Add11~125 .extended_lut = "off";
defparam \Add11~125 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~125 .shared_arith = "off";

cyclonev_lcell_comb \Add8~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~17_sumout ),
	.cout(\Add8~18 ),
	.shareout());
defparam \Add8~17 .extended_lut = "off";
defparam \Add8~17 .lut_mask = 64'h000000000000FF00;
defparam \Add8~17 .shared_arith = "off";

dffeas \M_div_src1[2] (
	.clk(clk_clk),
	.d(\Add8~17_sumout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[2]~q ),
	.prn(vcc));
defparam \M_div_src1[2] .is_wysiwyg = "true";
defparam \M_div_src1[2] .power_up = "low";

dffeas \A_div_rem[2] (
	.clk(clk_clk),
	.d(\Add11~125_sumout ),
	.asdata(\M_div_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[2]~q ),
	.prn(vcc));
defparam \A_div_rem[2] .is_wysiwyg = "true";
defparam \A_div_rem[2] .power_up = "low";

cyclonev_lcell_comb \Add11~121 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[2]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[2]~q ),
	.datag(gnd),
	.cin(\Add11~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~121_sumout ),
	.cout(\Add11~122 ),
	.shareout());
defparam \Add11~121 .extended_lut = "off";
defparam \Add11~121 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~121 .shared_arith = "off";

cyclonev_lcell_comb \Add8~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~21_sumout ),
	.cout(\Add8~22 ),
	.shareout());
defparam \Add8~21 .extended_lut = "off";
defparam \Add8~21 .lut_mask = 64'h000000000000FF00;
defparam \Add8~21 .shared_arith = "off";

dffeas \M_div_src1[3] (
	.clk(clk_clk),
	.d(\Add8~21_sumout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[3]~q ),
	.prn(vcc));
defparam \M_div_src1[3] .is_wysiwyg = "true";
defparam \M_div_src1[3] .power_up = "low";

dffeas \A_div_rem[3] (
	.clk(clk_clk),
	.d(\Add11~121_sumout ),
	.asdata(\M_div_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[3]~q ),
	.prn(vcc));
defparam \A_div_rem[3] .is_wysiwyg = "true";
defparam \A_div_rem[3] .power_up = "low";

cyclonev_lcell_comb \Add11~117 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[3]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[3]~q ),
	.datag(gnd),
	.cin(\Add11~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~117_sumout ),
	.cout(\Add11~118 ),
	.shareout());
defparam \Add11~117 .extended_lut = "off";
defparam \Add11~117 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~117 .shared_arith = "off";

cyclonev_lcell_comb \Add8~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~25_sumout ),
	.cout(\Add8~26 ),
	.shareout());
defparam \Add8~25 .extended_lut = "off";
defparam \Add8~25 .lut_mask = 64'h000000000000FF00;
defparam \Add8~25 .shared_arith = "off";

dffeas \M_div_src1[4] (
	.clk(clk_clk),
	.d(\Add8~25_sumout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[4]~q ),
	.prn(vcc));
defparam \M_div_src1[4] .is_wysiwyg = "true";
defparam \M_div_src1[4] .power_up = "low";

dffeas \A_div_rem[4] (
	.clk(clk_clk),
	.d(\Add11~117_sumout ),
	.asdata(\M_div_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[4]~q ),
	.prn(vcc));
defparam \A_div_rem[4] .is_wysiwyg = "true";
defparam \A_div_rem[4] .power_up = "low";

cyclonev_lcell_comb \Add11~113 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[4]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[4]~q ),
	.datag(gnd),
	.cin(\Add11~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~113_sumout ),
	.cout(\Add11~114 ),
	.shareout());
defparam \Add11~113 .extended_lut = "off";
defparam \Add11~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~113 .shared_arith = "off";

cyclonev_lcell_comb \Add8~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~29_sumout ),
	.cout(\Add8~30 ),
	.shareout());
defparam \Add8~29 .extended_lut = "off";
defparam \Add8~29 .lut_mask = 64'h000000000000FF00;
defparam \Add8~29 .shared_arith = "off";

dffeas \M_div_src1[5] (
	.clk(clk_clk),
	.d(\Add8~29_sumout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[5]~q ),
	.prn(vcc));
defparam \M_div_src1[5] .is_wysiwyg = "true";
defparam \M_div_src1[5] .power_up = "low";

dffeas \A_div_rem[5] (
	.clk(clk_clk),
	.d(\Add11~113_sumout ),
	.asdata(\M_div_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[5]~q ),
	.prn(vcc));
defparam \A_div_rem[5] .is_wysiwyg = "true";
defparam \A_div_rem[5] .power_up = "low";

cyclonev_lcell_comb \Add11~109 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[5]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[5]~q ),
	.datag(gnd),
	.cin(\Add11~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~109_sumout ),
	.cout(\Add11~110 ),
	.shareout());
defparam \Add11~109 .extended_lut = "off";
defparam \Add11~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~109 .shared_arith = "off";

cyclonev_lcell_comb \Add8~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~33_sumout ),
	.cout(\Add8~34 ),
	.shareout());
defparam \Add8~33 .extended_lut = "off";
defparam \Add8~33 .lut_mask = 64'h000000000000FF00;
defparam \Add8~33 .shared_arith = "off";

dffeas \M_div_src1[6] (
	.clk(clk_clk),
	.d(\Add8~33_sumout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[6]~q ),
	.prn(vcc));
defparam \M_div_src1[6] .is_wysiwyg = "true";
defparam \M_div_src1[6] .power_up = "low";

dffeas \A_div_rem[6] (
	.clk(clk_clk),
	.d(\Add11~109_sumout ),
	.asdata(\M_div_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[6]~q ),
	.prn(vcc));
defparam \A_div_rem[6] .is_wysiwyg = "true";
defparam \A_div_rem[6] .power_up = "low";

cyclonev_lcell_comb \Add11~105 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[6]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[6]~q ),
	.datag(gnd),
	.cin(\Add11~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~105_sumout ),
	.cout(\Add11~106 ),
	.shareout());
defparam \Add11~105 .extended_lut = "off";
defparam \Add11~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~105 .shared_arith = "off";

cyclonev_lcell_comb \Add8~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~37_sumout ),
	.cout(\Add8~38 ),
	.shareout());
defparam \Add8~37 .extended_lut = "off";
defparam \Add8~37 .lut_mask = 64'h000000000000FF00;
defparam \Add8~37 .shared_arith = "off";

dffeas \M_div_src1[7] (
	.clk(clk_clk),
	.d(\Add8~37_sumout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[7]~q ),
	.prn(vcc));
defparam \M_div_src1[7] .is_wysiwyg = "true";
defparam \M_div_src1[7] .power_up = "low";

dffeas \A_div_rem[7] (
	.clk(clk_clk),
	.d(\Add11~105_sumout ),
	.asdata(\M_div_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[7]~q ),
	.prn(vcc));
defparam \A_div_rem[7] .is_wysiwyg = "true";
defparam \A_div_rem[7] .power_up = "low";

cyclonev_lcell_comb \Add11~101 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[7]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[7]~q ),
	.datag(gnd),
	.cin(\Add11~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~101_sumout ),
	.cout(\Add11~102 ),
	.shareout());
defparam \Add11~101 .extended_lut = "off";
defparam \Add11~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~101 .shared_arith = "off";

cyclonev_lcell_comb \Add8~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~41_sumout ),
	.cout(\Add8~42 ),
	.shareout());
defparam \Add8~41 .extended_lut = "off";
defparam \Add8~41 .lut_mask = 64'h000000000000FF00;
defparam \Add8~41 .shared_arith = "off";

dffeas \M_div_src1[8] (
	.clk(clk_clk),
	.d(\Add8~41_sumout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[8]~q ),
	.prn(vcc));
defparam \M_div_src1[8] .is_wysiwyg = "true";
defparam \M_div_src1[8] .power_up = "low";

dffeas \A_div_rem[8] (
	.clk(clk_clk),
	.d(\Add11~101_sumout ),
	.asdata(\M_div_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[8]~q ),
	.prn(vcc));
defparam \A_div_rem[8] .is_wysiwyg = "true";
defparam \A_div_rem[8] .power_up = "low";

cyclonev_lcell_comb \Add11~97 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[8]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[8]~q ),
	.datag(gnd),
	.cin(\Add11~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~97_sumout ),
	.cout(\Add11~98 ),
	.shareout());
defparam \Add11~97 .extended_lut = "off";
defparam \Add11~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~97 .shared_arith = "off";

cyclonev_lcell_comb \Add8~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~45_sumout ),
	.cout(\Add8~46 ),
	.shareout());
defparam \Add8~45 .extended_lut = "off";
defparam \Add8~45 .lut_mask = 64'h000000000000FF00;
defparam \Add8~45 .shared_arith = "off";

dffeas \M_div_src1[9] (
	.clk(clk_clk),
	.d(\Add8~45_sumout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[9]~q ),
	.prn(vcc));
defparam \M_div_src1[9] .is_wysiwyg = "true";
defparam \M_div_src1[9] .power_up = "low";

dffeas \A_div_rem[9] (
	.clk(clk_clk),
	.d(\Add11~97_sumout ),
	.asdata(\M_div_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[9]~q ),
	.prn(vcc));
defparam \A_div_rem[9] .is_wysiwyg = "true";
defparam \A_div_rem[9] .power_up = "low";

cyclonev_lcell_comb \Add11~93 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[9]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[9]~q ),
	.datag(gnd),
	.cin(\Add11~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~93_sumout ),
	.cout(\Add11~94 ),
	.shareout());
defparam \Add11~93 .extended_lut = "off";
defparam \Add11~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~93 .shared_arith = "off";

cyclonev_lcell_comb \Add8~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~49_sumout ),
	.cout(\Add8~50 ),
	.shareout());
defparam \Add8~49 .extended_lut = "off";
defparam \Add8~49 .lut_mask = 64'h000000000000FF00;
defparam \Add8~49 .shared_arith = "off";

dffeas \M_div_src1[10] (
	.clk(clk_clk),
	.d(\Add8~49_sumout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[10]~q ),
	.prn(vcc));
defparam \M_div_src1[10] .is_wysiwyg = "true";
defparam \M_div_src1[10] .power_up = "low";

dffeas \A_div_rem[10] (
	.clk(clk_clk),
	.d(\Add11~93_sumout ),
	.asdata(\M_div_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[10]~q ),
	.prn(vcc));
defparam \A_div_rem[10] .is_wysiwyg = "true";
defparam \A_div_rem[10] .power_up = "low";

cyclonev_lcell_comb \Add11~89 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[10]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[10]~q ),
	.datag(gnd),
	.cin(\Add11~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~89_sumout ),
	.cout(\Add11~90 ),
	.shareout());
defparam \Add11~89 .extended_lut = "off";
defparam \Add11~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~89 .shared_arith = "off";

cyclonev_lcell_comb \Add8~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~53_sumout ),
	.cout(\Add8~54 ),
	.shareout());
defparam \Add8~53 .extended_lut = "off";
defparam \Add8~53 .lut_mask = 64'h000000000000FF00;
defparam \Add8~53 .shared_arith = "off";

dffeas \M_div_src1[11] (
	.clk(clk_clk),
	.d(\Add8~53_sumout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[11]~q ),
	.prn(vcc));
defparam \M_div_src1[11] .is_wysiwyg = "true";
defparam \M_div_src1[11] .power_up = "low";

dffeas \A_div_rem[11] (
	.clk(clk_clk),
	.d(\Add11~89_sumout ),
	.asdata(\M_div_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[11]~q ),
	.prn(vcc));
defparam \A_div_rem[11] .is_wysiwyg = "true";
defparam \A_div_rem[11] .power_up = "low";

cyclonev_lcell_comb \Add11~85 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[11]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[11]~q ),
	.datag(gnd),
	.cin(\Add11~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~85_sumout ),
	.cout(\Add11~86 ),
	.shareout());
defparam \Add11~85 .extended_lut = "off";
defparam \Add11~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~85 .shared_arith = "off";

cyclonev_lcell_comb \Add8~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~57_sumout ),
	.cout(\Add8~58 ),
	.shareout());
defparam \Add8~57 .extended_lut = "off";
defparam \Add8~57 .lut_mask = 64'h000000000000FF00;
defparam \Add8~57 .shared_arith = "off";

dffeas \M_div_src1[12] (
	.clk(clk_clk),
	.d(\Add8~57_sumout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[12]~q ),
	.prn(vcc));
defparam \M_div_src1[12] .is_wysiwyg = "true";
defparam \M_div_src1[12] .power_up = "low";

dffeas \A_div_rem[12] (
	.clk(clk_clk),
	.d(\Add11~85_sumout ),
	.asdata(\M_div_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[12]~q ),
	.prn(vcc));
defparam \A_div_rem[12] .is_wysiwyg = "true";
defparam \A_div_rem[12] .power_up = "low";

cyclonev_lcell_comb \Add11~81 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[12]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[12]~q ),
	.datag(gnd),
	.cin(\Add11~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~81_sumout ),
	.cout(\Add11~82 ),
	.shareout());
defparam \Add11~81 .extended_lut = "off";
defparam \Add11~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~81 .shared_arith = "off";

cyclonev_lcell_comb \Add8~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~61_sumout ),
	.cout(\Add8~62 ),
	.shareout());
defparam \Add8~61 .extended_lut = "off";
defparam \Add8~61 .lut_mask = 64'h000000000000FF00;
defparam \Add8~61 .shared_arith = "off";

dffeas \M_div_src1[13] (
	.clk(clk_clk),
	.d(\Add8~61_sumout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[13]~q ),
	.prn(vcc));
defparam \M_div_src1[13] .is_wysiwyg = "true";
defparam \M_div_src1[13] .power_up = "low";

dffeas \A_div_rem[13] (
	.clk(clk_clk),
	.d(\Add11~81_sumout ),
	.asdata(\M_div_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[13]~q ),
	.prn(vcc));
defparam \A_div_rem[13] .is_wysiwyg = "true";
defparam \A_div_rem[13] .power_up = "low";

cyclonev_lcell_comb \Add11~77 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[13]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[13]~q ),
	.datag(gnd),
	.cin(\Add11~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~77_sumout ),
	.cout(\Add11~78 ),
	.shareout());
defparam \Add11~77 .extended_lut = "off";
defparam \Add11~77 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~77 .shared_arith = "off";

cyclonev_lcell_comb \Add8~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~65_sumout ),
	.cout(\Add8~66 ),
	.shareout());
defparam \Add8~65 .extended_lut = "off";
defparam \Add8~65 .lut_mask = 64'h000000000000FF00;
defparam \Add8~65 .shared_arith = "off";

dffeas \M_div_src1[14] (
	.clk(clk_clk),
	.d(\Add8~65_sumout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[14]~q ),
	.prn(vcc));
defparam \M_div_src1[14] .is_wysiwyg = "true";
defparam \M_div_src1[14] .power_up = "low";

dffeas \A_div_rem[14] (
	.clk(clk_clk),
	.d(\Add11~77_sumout ),
	.asdata(\M_div_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[14]~q ),
	.prn(vcc));
defparam \A_div_rem[14] .is_wysiwyg = "true";
defparam \A_div_rem[14] .power_up = "low";

cyclonev_lcell_comb \Add11~73 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[14]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[14]~q ),
	.datag(gnd),
	.cin(\Add11~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~73_sumout ),
	.cout(\Add11~74 ),
	.shareout());
defparam \Add11~73 .extended_lut = "off";
defparam \Add11~73 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~73 .shared_arith = "off";

cyclonev_lcell_comb \Add8~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~69_sumout ),
	.cout(\Add8~70 ),
	.shareout());
defparam \Add8~69 .extended_lut = "off";
defparam \Add8~69 .lut_mask = 64'h000000000000FF00;
defparam \Add8~69 .shared_arith = "off";

dffeas \M_div_src1[15] (
	.clk(clk_clk),
	.d(\Add8~69_sumout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[15]~q ),
	.prn(vcc));
defparam \M_div_src1[15] .is_wysiwyg = "true";
defparam \M_div_src1[15] .power_up = "low";

dffeas \A_div_rem[15] (
	.clk(clk_clk),
	.d(\Add11~73_sumout ),
	.asdata(\M_div_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[15]~q ),
	.prn(vcc));
defparam \A_div_rem[15] .is_wysiwyg = "true";
defparam \A_div_rem[15] .power_up = "low";

cyclonev_lcell_comb \Add11~69 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[15]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[15]~q ),
	.datag(gnd),
	.cin(\Add11~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~69_sumout ),
	.cout(\Add11~70 ),
	.shareout());
defparam \Add11~69 .extended_lut = "off";
defparam \Add11~69 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~69 .shared_arith = "off";

cyclonev_lcell_comb \Add8~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~77_sumout ),
	.cout(\Add8~78 ),
	.shareout());
defparam \Add8~77 .extended_lut = "off";
defparam \Add8~77 .lut_mask = 64'h000000000000FF00;
defparam \Add8~77 .shared_arith = "off";

dffeas \M_div_src1[16] (
	.clk(clk_clk),
	.d(\Add8~77_sumout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[16]~q ),
	.prn(vcc));
defparam \M_div_src1[16] .is_wysiwyg = "true";
defparam \M_div_src1[16] .power_up = "low";

dffeas \A_div_rem[16] (
	.clk(clk_clk),
	.d(\Add11~69_sumout ),
	.asdata(\M_div_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[16]~q ),
	.prn(vcc));
defparam \A_div_rem[16] .is_wysiwyg = "true";
defparam \A_div_rem[16] .power_up = "low";

cyclonev_lcell_comb \Add11~65 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[16]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[16]~q ),
	.datag(gnd),
	.cin(\Add11~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~65_sumout ),
	.cout(\Add11~66 ),
	.shareout());
defparam \Add11~65 .extended_lut = "off";
defparam \Add11~65 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~65 .shared_arith = "off";

cyclonev_lcell_comb \Add8~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~81_sumout ),
	.cout(\Add8~82 ),
	.shareout());
defparam \Add8~81 .extended_lut = "off";
defparam \Add8~81 .lut_mask = 64'h000000000000FF00;
defparam \Add8~81 .shared_arith = "off";

dffeas \M_div_src1[17] (
	.clk(clk_clk),
	.d(\Add8~81_sumout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[17]~q ),
	.prn(vcc));
defparam \M_div_src1[17] .is_wysiwyg = "true";
defparam \M_div_src1[17] .power_up = "low";

dffeas \A_div_rem[17] (
	.clk(clk_clk),
	.d(\Add11~65_sumout ),
	.asdata(\M_div_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[17]~q ),
	.prn(vcc));
defparam \A_div_rem[17] .is_wysiwyg = "true";
defparam \A_div_rem[17] .power_up = "low";

cyclonev_lcell_comb \Add11~61 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[17]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[17]~q ),
	.datag(gnd),
	.cin(\Add11~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~61_sumout ),
	.cout(\Add11~62 ),
	.shareout());
defparam \Add11~61 .extended_lut = "off";
defparam \Add11~61 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~61 .shared_arith = "off";

cyclonev_lcell_comb \Add8~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~85_sumout ),
	.cout(\Add8~86 ),
	.shareout());
defparam \Add8~85 .extended_lut = "off";
defparam \Add8~85 .lut_mask = 64'h000000000000FF00;
defparam \Add8~85 .shared_arith = "off";

dffeas \M_div_src1[18] (
	.clk(clk_clk),
	.d(\Add8~85_sumout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[18]~q ),
	.prn(vcc));
defparam \M_div_src1[18] .is_wysiwyg = "true";
defparam \M_div_src1[18] .power_up = "low";

dffeas \A_div_rem[18] (
	.clk(clk_clk),
	.d(\Add11~61_sumout ),
	.asdata(\M_div_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[18]~q ),
	.prn(vcc));
defparam \A_div_rem[18] .is_wysiwyg = "true";
defparam \A_div_rem[18] .power_up = "low";

cyclonev_lcell_comb \Add11~57 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[18]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[18]~q ),
	.datag(gnd),
	.cin(\Add11~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~57_sumout ),
	.cout(\Add11~58 ),
	.shareout());
defparam \Add11~57 .extended_lut = "off";
defparam \Add11~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~57 .shared_arith = "off";

cyclonev_lcell_comb \Add8~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~89_sumout ),
	.cout(\Add8~90 ),
	.shareout());
defparam \Add8~89 .extended_lut = "off";
defparam \Add8~89 .lut_mask = 64'h000000000000FF00;
defparam \Add8~89 .shared_arith = "off";

dffeas \M_div_src1[19] (
	.clk(clk_clk),
	.d(\Add8~89_sumout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[19]~q ),
	.prn(vcc));
defparam \M_div_src1[19] .is_wysiwyg = "true";
defparam \M_div_src1[19] .power_up = "low";

dffeas \A_div_rem[19] (
	.clk(clk_clk),
	.d(\Add11~57_sumout ),
	.asdata(\M_div_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[19]~q ),
	.prn(vcc));
defparam \A_div_rem[19] .is_wysiwyg = "true";
defparam \A_div_rem[19] .power_up = "low";

cyclonev_lcell_comb \Add11~53 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[19]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[19]~q ),
	.datag(gnd),
	.cin(\Add11~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~53_sumout ),
	.cout(\Add11~54 ),
	.shareout());
defparam \Add11~53 .extended_lut = "off";
defparam \Add11~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~53 .shared_arith = "off";

cyclonev_lcell_comb \Add8~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~93_sumout ),
	.cout(\Add8~94 ),
	.shareout());
defparam \Add8~93 .extended_lut = "off";
defparam \Add8~93 .lut_mask = 64'h000000000000FF00;
defparam \Add8~93 .shared_arith = "off";

dffeas \M_div_src1[20] (
	.clk(clk_clk),
	.d(\Add8~93_sumout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[20]~q ),
	.prn(vcc));
defparam \M_div_src1[20] .is_wysiwyg = "true";
defparam \M_div_src1[20] .power_up = "low";

dffeas \A_div_rem[20] (
	.clk(clk_clk),
	.d(\Add11~53_sumout ),
	.asdata(\M_div_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[20]~q ),
	.prn(vcc));
defparam \A_div_rem[20] .is_wysiwyg = "true";
defparam \A_div_rem[20] .power_up = "low";

cyclonev_lcell_comb \Add11~49 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[20]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[20]~q ),
	.datag(gnd),
	.cin(\Add11~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~49_sumout ),
	.cout(\Add11~50 ),
	.shareout());
defparam \Add11~49 .extended_lut = "off";
defparam \Add11~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~49 .shared_arith = "off";

cyclonev_lcell_comb \Add8~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~97_sumout ),
	.cout(\Add8~98 ),
	.shareout());
defparam \Add8~97 .extended_lut = "off";
defparam \Add8~97 .lut_mask = 64'h000000000000FF00;
defparam \Add8~97 .shared_arith = "off";

dffeas \M_div_src1[21] (
	.clk(clk_clk),
	.d(\Add8~97_sumout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[21]~q ),
	.prn(vcc));
defparam \M_div_src1[21] .is_wysiwyg = "true";
defparam \M_div_src1[21] .power_up = "low";

dffeas \A_div_rem[21] (
	.clk(clk_clk),
	.d(\Add11~49_sumout ),
	.asdata(\M_div_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[21]~q ),
	.prn(vcc));
defparam \A_div_rem[21] .is_wysiwyg = "true";
defparam \A_div_rem[21] .power_up = "low";

cyclonev_lcell_comb \Add11~45 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[21]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[21]~q ),
	.datag(gnd),
	.cin(\Add11~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~45_sumout ),
	.cout(\Add11~46 ),
	.shareout());
defparam \Add11~45 .extended_lut = "off";
defparam \Add11~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~45 .shared_arith = "off";

cyclonev_lcell_comb \Add8~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~101_sumout ),
	.cout(\Add8~102 ),
	.shareout());
defparam \Add8~101 .extended_lut = "off";
defparam \Add8~101 .lut_mask = 64'h000000000000FF00;
defparam \Add8~101 .shared_arith = "off";

dffeas \M_div_src1[22] (
	.clk(clk_clk),
	.d(\Add8~101_sumout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[22]~q ),
	.prn(vcc));
defparam \M_div_src1[22] .is_wysiwyg = "true";
defparam \M_div_src1[22] .power_up = "low";

dffeas \A_div_rem[22] (
	.clk(clk_clk),
	.d(\Add11~45_sumout ),
	.asdata(\M_div_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[22]~q ),
	.prn(vcc));
defparam \A_div_rem[22] .is_wysiwyg = "true";
defparam \A_div_rem[22] .power_up = "low";

cyclonev_lcell_comb \Add11~41 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[22]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[22]~q ),
	.datag(gnd),
	.cin(\Add11~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~41_sumout ),
	.cout(\Add11~42 ),
	.shareout());
defparam \Add11~41 .extended_lut = "off";
defparam \Add11~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~41 .shared_arith = "off";

cyclonev_lcell_comb \Add8~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~105_sumout ),
	.cout(\Add8~106 ),
	.shareout());
defparam \Add8~105 .extended_lut = "off";
defparam \Add8~105 .lut_mask = 64'h000000000000FF00;
defparam \Add8~105 .shared_arith = "off";

dffeas \M_div_src1[23] (
	.clk(clk_clk),
	.d(\Add8~105_sumout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[23]~q ),
	.prn(vcc));
defparam \M_div_src1[23] .is_wysiwyg = "true";
defparam \M_div_src1[23] .power_up = "low";

dffeas \A_div_rem[23] (
	.clk(clk_clk),
	.d(\Add11~41_sumout ),
	.asdata(\M_div_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[23]~q ),
	.prn(vcc));
defparam \A_div_rem[23] .is_wysiwyg = "true";
defparam \A_div_rem[23] .power_up = "low";

cyclonev_lcell_comb \Add11~37 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[23]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[23]~q ),
	.datag(gnd),
	.cin(\Add11~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~37_sumout ),
	.cout(\Add11~38 ),
	.shareout());
defparam \Add11~37 .extended_lut = "off";
defparam \Add11~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~37 .shared_arith = "off";

cyclonev_lcell_comb \Add8~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~109_sumout ),
	.cout(\Add8~110 ),
	.shareout());
defparam \Add8~109 .extended_lut = "off";
defparam \Add8~109 .lut_mask = 64'h000000000000FF00;
defparam \Add8~109 .shared_arith = "off";

dffeas \M_div_src1[24] (
	.clk(clk_clk),
	.d(\Add8~109_sumout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[24]~q ),
	.prn(vcc));
defparam \M_div_src1[24] .is_wysiwyg = "true";
defparam \M_div_src1[24] .power_up = "low";

dffeas \A_div_rem[24] (
	.clk(clk_clk),
	.d(\Add11~37_sumout ),
	.asdata(\M_div_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[24]~q ),
	.prn(vcc));
defparam \A_div_rem[24] .is_wysiwyg = "true";
defparam \A_div_rem[24] .power_up = "low";

cyclonev_lcell_comb \Add11~33 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[24]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[24]~q ),
	.datag(gnd),
	.cin(\Add11~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~33_sumout ),
	.cout(\Add11~34 ),
	.shareout());
defparam \Add11~33 .extended_lut = "off";
defparam \Add11~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~33 .shared_arith = "off";

cyclonev_lcell_comb \Add8~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~113_sumout ),
	.cout(\Add8~114 ),
	.shareout());
defparam \Add8~113 .extended_lut = "off";
defparam \Add8~113 .lut_mask = 64'h000000000000FF00;
defparam \Add8~113 .shared_arith = "off";

dffeas \M_div_src1[25] (
	.clk(clk_clk),
	.d(\Add8~113_sumout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[25]~q ),
	.prn(vcc));
defparam \M_div_src1[25] .is_wysiwyg = "true";
defparam \M_div_src1[25] .power_up = "low";

dffeas \A_div_rem[25] (
	.clk(clk_clk),
	.d(\Add11~33_sumout ),
	.asdata(\M_div_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[25]~q ),
	.prn(vcc));
defparam \A_div_rem[25] .is_wysiwyg = "true";
defparam \A_div_rem[25] .power_up = "low";

cyclonev_lcell_comb \Add11~29 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[25]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[25]~q ),
	.datag(gnd),
	.cin(\Add11~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~29_sumout ),
	.cout(\Add11~30 ),
	.shareout());
defparam \Add11~29 .extended_lut = "off";
defparam \Add11~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~29 .shared_arith = "off";

cyclonev_lcell_comb \Add8~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~117_sumout ),
	.cout(\Add8~118 ),
	.shareout());
defparam \Add8~117 .extended_lut = "off";
defparam \Add8~117 .lut_mask = 64'h000000000000FF00;
defparam \Add8~117 .shared_arith = "off";

dffeas \M_div_src1[26] (
	.clk(clk_clk),
	.d(\Add8~117_sumout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[26]~q ),
	.prn(vcc));
defparam \M_div_src1[26] .is_wysiwyg = "true";
defparam \M_div_src1[26] .power_up = "low";

dffeas \A_div_rem[26] (
	.clk(clk_clk),
	.d(\Add11~29_sumout ),
	.asdata(\M_div_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[26]~q ),
	.prn(vcc));
defparam \A_div_rem[26] .is_wysiwyg = "true";
defparam \A_div_rem[26] .power_up = "low";

cyclonev_lcell_comb \Add11~25 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[26]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[26]~q ),
	.datag(gnd),
	.cin(\Add11~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~25_sumout ),
	.cout(\Add11~26 ),
	.shareout());
defparam \Add11~25 .extended_lut = "off";
defparam \Add11~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~25 .shared_arith = "off";

cyclonev_lcell_comb \Add8~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~121_sumout ),
	.cout(\Add8~122 ),
	.shareout());
defparam \Add8~121 .extended_lut = "off";
defparam \Add8~121 .lut_mask = 64'h000000000000FF00;
defparam \Add8~121 .shared_arith = "off";

dffeas \M_div_src1[27] (
	.clk(clk_clk),
	.d(\Add8~121_sumout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[27]~q ),
	.prn(vcc));
defparam \M_div_src1[27] .is_wysiwyg = "true";
defparam \M_div_src1[27] .power_up = "low";

dffeas \A_div_rem[27] (
	.clk(clk_clk),
	.d(\Add11~25_sumout ),
	.asdata(\M_div_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[27]~q ),
	.prn(vcc));
defparam \A_div_rem[27] .is_wysiwyg = "true";
defparam \A_div_rem[27] .power_up = "low";

cyclonev_lcell_comb \Add11~21 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[27]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[27]~q ),
	.datag(gnd),
	.cin(\Add11~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~21_sumout ),
	.cout(\Add11~22 ),
	.shareout());
defparam \Add11~21 .extended_lut = "off";
defparam \Add11~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~21 .shared_arith = "off";

cyclonev_lcell_comb \Add8~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~125_sumout ),
	.cout(\Add8~126 ),
	.shareout());
defparam \Add8~125 .extended_lut = "off";
defparam \Add8~125 .lut_mask = 64'h000000000000FF00;
defparam \Add8~125 .shared_arith = "off";

dffeas \M_div_src1[28] (
	.clk(clk_clk),
	.d(\Add8~125_sumout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[28]~q ),
	.prn(vcc));
defparam \M_div_src1[28] .is_wysiwyg = "true";
defparam \M_div_src1[28] .power_up = "low";

dffeas \A_div_rem[28] (
	.clk(clk_clk),
	.d(\Add11~21_sumout ),
	.asdata(\M_div_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[28]~q ),
	.prn(vcc));
defparam \A_div_rem[28] .is_wysiwyg = "true";
defparam \A_div_rem[28] .power_up = "low";

cyclonev_lcell_comb \Add11~17 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[28]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[28]~q ),
	.datag(gnd),
	.cin(\Add11~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~17_sumout ),
	.cout(\Add11~18 ),
	.shareout());
defparam \Add11~17 .extended_lut = "off";
defparam \Add11~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~17 .shared_arith = "off";

cyclonev_lcell_comb \Add8~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~73_sumout ),
	.cout(\Add8~74 ),
	.shareout());
defparam \Add8~73 .extended_lut = "off";
defparam \Add8~73 .lut_mask = 64'h000000000000FF00;
defparam \Add8~73 .shared_arith = "off";

dffeas \M_div_src1[29] (
	.clk(clk_clk),
	.d(\Add8~73_sumout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[29]~q ),
	.prn(vcc));
defparam \M_div_src1[29] .is_wysiwyg = "true";
defparam \M_div_src1[29] .power_up = "low";

dffeas \A_div_rem[29] (
	.clk(clk_clk),
	.d(\Add11~17_sumout ),
	.asdata(\M_div_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[29]~q ),
	.prn(vcc));
defparam \A_div_rem[29] .is_wysiwyg = "true";
defparam \A_div_rem[29] .power_up = "low";

cyclonev_lcell_comb \Add11~13 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[29]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[29]~q ),
	.datag(gnd),
	.cin(\Add11~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~13_sumout ),
	.cout(\Add11~14 ),
	.shareout());
defparam \Add11~13 .extended_lut = "off";
defparam \Add11~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~13 .shared_arith = "off";

cyclonev_lcell_comb \Add8~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~5_sumout ),
	.cout(\Add8~6 ),
	.shareout());
defparam \Add8~5 .extended_lut = "off";
defparam \Add8~5 .lut_mask = 64'h000000000000FF00;
defparam \Add8~5 .shared_arith = "off";

dffeas \M_div_src1[30] (
	.clk(clk_clk),
	.d(\Add8~5_sumout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[30]~q ),
	.prn(vcc));
defparam \M_div_src1[30] .is_wysiwyg = "true";
defparam \M_div_src1[30] .power_up = "low";

dffeas \A_div_rem[30] (
	.clk(clk_clk),
	.d(\Add11~13_sumout ),
	.asdata(\M_div_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[30]~q ),
	.prn(vcc));
defparam \A_div_rem[30] .is_wysiwyg = "true";
defparam \A_div_rem[30] .power_up = "low";

cyclonev_lcell_comb \Add11~9 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[30]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[30]~q ),
	.datag(gnd),
	.cin(\Add11~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~9_sumout ),
	.cout(\Add11~10 ),
	.shareout());
defparam \Add11~9 .extended_lut = "off";
defparam \Add11~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~9 .shared_arith = "off";

cyclonev_lcell_comb \Add8~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src1[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~1_sumout ),
	.cout(),
	.shareout());
defparam \Add8~1 .extended_lut = "off";
defparam \Add8~1 .lut_mask = 64'h000000000000FF00;
defparam \Add8~1 .shared_arith = "off";

dffeas \M_div_src1[31] (
	.clk(clk_clk),
	.d(\Add8~1_sumout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_div_negate_src1~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_div_src1[31]~q ),
	.prn(vcc));
defparam \M_div_src1[31] .is_wysiwyg = "true";
defparam \M_div_src1[31] .power_up = "low";

dffeas \A_div_rem[31] (
	.clk(clk_clk),
	.d(\Add11~9_sumout ),
	.asdata(\M_div_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_stall~combout ),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[31]~q ),
	.prn(vcc));
defparam \A_div_rem[31] .is_wysiwyg = "true";
defparam \A_div_rem[31] .power_up = "low";

cyclonev_lcell_comb \Add11~5 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_den[31]~q ),
	.datae(gnd),
	.dataf(!\A_div_rem[31]~q ),
	.datag(gnd),
	.cin(\Add11~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~5_sumout ),
	.cout(\Add11~6 ),
	.shareout());
defparam \Add11~5 .extended_lut = "off";
defparam \Add11~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~5 .shared_arith = "off";

dffeas \A_div_rem[32] (
	.clk(clk_clk),
	.d(\Add11~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(\A_div_rem_en~combout ),
	.q(\A_div_rem[32]~q ),
	.prn(vcc));
defparam \A_div_rem[32] .is_wysiwyg = "true";
defparam \A_div_rem[32] .power_up = "low";

cyclonev_lcell_comb \Add11~1 (
	.dataa(!\A_div_do_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_rem[32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~1_sumout ),
	.cout(),
	.shareout());
defparam \Add11~1 .extended_lut = "off";
defparam \Add11~1 .lut_mask = 64'h0000AAAA000000FF;
defparam \Add11~1 .shared_arith = "off";

cyclonev_lcell_comb A_div_discover_quotient_bits(
	.dataa(!\Add11~1_sumout ),
	.datab(!\A_div_discover_quotient_bits~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_discover_quotient_bits~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_div_discover_quotient_bits.extended_lut = "off";
defparam A_div_discover_quotient_bits.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam A_div_discover_quotient_bits.shared_arith = "off";

cyclonev_lcell_comb \Add13~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~9_sumout ),
	.cout(\Add13~10 ),
	.shareout());
defparam \Add13~9 .extended_lut = "off";
defparam \Add13~9 .lut_mask = 64'h00000000000000FF;
defparam \Add13~9 .shared_arith = "off";

cyclonev_lcell_comb \A_div_norm_cnt_nxt[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\Add13~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_norm_cnt_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_norm_cnt_nxt[0]~0 .extended_lut = "off";
defparam \A_div_norm_cnt_nxt[0]~0 .lut_mask = 64'h7777777777777777;
defparam \A_div_norm_cnt_nxt[0]~0 .shared_arith = "off";

dffeas \A_div_norm_cnt[0] (
	.clk(clk_clk),
	.d(\A_div_norm_cnt_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[0]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[0] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add13~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[1]~q ),
	.datae(gnd),
	.dataf(!\A_div_discover_quotient_bits~combout ),
	.datag(gnd),
	.cin(\Add13~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~17_sumout ),
	.cout(\Add13~18 ),
	.shareout());
defparam \Add13~17 .extended_lut = "off";
defparam \Add13~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add13~17 .shared_arith = "off";

dffeas \A_div_norm_cnt[1] (
	.clk(clk_clk),
	.d(\Add13~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[1]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[1] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add13~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[2]~q ),
	.datae(gnd),
	.dataf(!\A_div_discover_quotient_bits~combout ),
	.datag(gnd),
	.cin(\Add13~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~21_sumout ),
	.cout(\Add13~22 ),
	.shareout());
defparam \Add13~21 .extended_lut = "off";
defparam \Add13~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add13~21 .shared_arith = "off";

dffeas \A_div_norm_cnt[2] (
	.clk(clk_clk),
	.d(\Add13~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[2]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[2] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add13~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[3]~q ),
	.datae(gnd),
	.dataf(!\A_div_discover_quotient_bits~combout ),
	.datag(gnd),
	.cin(\Add13~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~5_sumout ),
	.cout(\Add13~6 ),
	.shareout());
defparam \Add13~5 .extended_lut = "off";
defparam \Add13~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add13~5 .shared_arith = "off";

dffeas \A_div_norm_cnt[3] (
	.clk(clk_clk),
	.d(\Add13~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[3]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[3] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Add13~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[4]~q ),
	.datae(gnd),
	.dataf(!\A_div_discover_quotient_bits~combout ),
	.datag(gnd),
	.cin(\Add13~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~13_sumout ),
	.cout(\Add13~14 ),
	.shareout());
defparam \Add13~13 .extended_lut = "off";
defparam \Add13~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add13~13 .shared_arith = "off";

dffeas \A_div_norm_cnt[4] (
	.clk(clk_clk),
	.d(\Add13~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[4]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[4] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Add13~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_div_norm_cnt[5]~q ),
	.datae(gnd),
	.dataf(!\A_div_discover_quotient_bits~combout ),
	.datag(gnd),
	.cin(\Add13~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~1_sumout ),
	.cout(),
	.shareout());
defparam \Add13~1 .extended_lut = "off";
defparam \Add13~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add13~1 .shared_arith = "off";

dffeas \A_div_norm_cnt[5] (
	.clk(clk_clk),
	.d(\Add13~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_norm_cnt[5]~q ),
	.prn(vcc));
defparam \A_div_norm_cnt[5] .is_wysiwyg = "true";
defparam \A_div_norm_cnt[5] .power_up = "low";

cyclonev_lcell_comb \A_div_last_quotient_bit_nxt~0 (
	.dataa(!\A_div_norm_cnt[0]~q ),
	.datab(!\A_div_norm_cnt[4]~q ),
	.datac(!\A_div_norm_cnt[1]~q ),
	.datad(!\A_div_norm_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_last_quotient_bit_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_div_last_quotient_bit_nxt~0 .extended_lut = "off";
defparam \A_div_last_quotient_bit_nxt~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \A_div_last_quotient_bit_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb A_div_last_quotient_bit_nxt(
	.dataa(!\A_div_norm_cnt[5]~q ),
	.datab(!\Add11~1_sumout ),
	.datac(!\A_div_norm_cnt[3]~q ),
	.datad(!\A_div_discover_quotient_bits~0_combout ),
	.datae(!\A_div_last_quotient_bit_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_div_last_quotient_bit_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_div_last_quotient_bit_nxt.extended_lut = "off";
defparam A_div_last_quotient_bit_nxt.lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam A_div_last_quotient_bit_nxt.shared_arith = "off";

dffeas A_div_last_quotient_bit(
	.clk(clk_clk),
	.d(\A_div_last_quotient_bit_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_last_quotient_bit~q ),
	.prn(vcc));
defparam A_div_last_quotient_bit.is_wysiwyg = "true";
defparam A_div_last_quotient_bit.power_up = "low";

dffeas A_div_quot_ready(
	.clk(clk_clk),
	.d(\A_div_last_quotient_bit~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_quot_ready~q ),
	.prn(vcc));
defparam A_div_quot_ready.is_wysiwyg = "true";
defparam A_div_quot_ready.power_up = "low";

dffeas A_div_done(
	.clk(clk_clk),
	.d(\A_div_quot_ready~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_div_done~q ),
	.prn(vcc));
defparam A_div_done.is_wysiwyg = "true";
defparam A_div_done.power_up = "low";

cyclonev_lcell_comb A_stall(
	.dataa(!\A_valid~q ),
	.datab(!\A_ctrl_div~q ),
	.datac(!\A_div_done~q ),
	.datad(!\A_mem_stall~q ),
	.datae(!\A_mul_stall~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_stall.extended_lut = "off";
defparam A_stall.lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam A_stall.shared_arith = "off";

dffeas M_ctrl_late_result(
	.clk(clk_clk),
	.d(\E_ctrl_late_result~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_late_result~q ),
	.prn(vcc));
defparam M_ctrl_late_result.is_wysiwyg = "true";
defparam M_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \D_data_depend~1 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\D_ctrl_b_is_dst~q ),
	.datac(!\M_ctrl_late_result~q ),
	.datad(!\M_regnum_b_cmp_D~q ),
	.datae(!\M_regnum_a_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~1 .extended_lut = "off";
defparam \D_data_depend~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_data_depend~1 .shared_arith = "off";

cyclonev_lcell_comb \D_dep_stall~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_issue~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dep_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dep_stall~0 .extended_lut = "off";
defparam \D_dep_stall~0 .lut_mask = 64'h7777777777777777;
defparam \D_dep_stall~0 .shared_arith = "off";

cyclonev_lcell_comb F_stall(
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_stall.extended_lut = "off";
defparam F_stall.lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam F_stall.shared_arith = "off";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_break~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_ctrl_logic~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~0 .extended_lut = "off";
defparam \D_ctrl_break~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_ctrl_break~0 .shared_arith = "off";

dffeas E_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_break~q ),
	.prn(vcc));
defparam E_ctrl_break.is_wysiwyg = "true";
defparam E_ctrl_break.power_up = "low";

dffeas M_ctrl_break(
	.clk(clk_clk),
	.d(\E_ctrl_break~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_break~q ),
	.prn(vcc));
defparam M_ctrl_break.is_wysiwyg = "true";
defparam M_ctrl_break.power_up = "low";

dffeas \M_iw[14] (
	.clk(clk_clk),
	.d(\E_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[14]~q ),
	.prn(vcc));
defparam \M_iw[14] .is_wysiwyg = "true";
defparam \M_iw[14] .power_up = "low";

dffeas \M_iw[11] (
	.clk(clk_clk),
	.d(\E_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[11]~q ),
	.prn(vcc));
defparam \M_iw[11] .is_wysiwyg = "true";
defparam \M_iw[11] .power_up = "low";

dffeas \M_iw[5] (
	.clk(clk_clk),
	.d(\E_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[5]~q ),
	.prn(vcc));
defparam \M_iw[5] .is_wysiwyg = "true";
defparam \M_iw[5] .power_up = "low";

dffeas \M_iw[0] (
	.clk(clk_clk),
	.d(\E_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[0]~q ),
	.prn(vcc));
defparam \M_iw[0] .is_wysiwyg = "true";
defparam \M_iw[0] .power_up = "low";

dffeas \M_iw[16] (
	.clk(clk_clk),
	.d(\E_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[16]~q ),
	.prn(vcc));
defparam \M_iw[16] .is_wysiwyg = "true";
defparam \M_iw[16] .power_up = "low";

dffeas \M_iw[15] (
	.clk(clk_clk),
	.d(\E_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[15]~q ),
	.prn(vcc));
defparam \M_iw[15] .is_wysiwyg = "true";
defparam \M_iw[15] .power_up = "low";

dffeas \M_iw[13] (
	.clk(clk_clk),
	.d(\E_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[13]~q ),
	.prn(vcc));
defparam \M_iw[13] .is_wysiwyg = "true";
defparam \M_iw[13] .power_up = "low";

dffeas \M_iw[12] (
	.clk(clk_clk),
	.d(\E_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[12]~q ),
	.prn(vcc));
defparam \M_iw[12] .is_wysiwyg = "true";
defparam \M_iw[12] .power_up = "low";

cyclonev_lcell_comb \M_op_eret~0 (
	.dataa(!\M_iw[16]~q ),
	.datab(!\M_iw[15]~q ),
	.datac(!\M_iw[13]~q ),
	.datad(!\M_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~0 .extended_lut = "off";
defparam \M_op_eret~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \M_op_eret~0 .shared_arith = "off";

dffeas \M_iw[4] (
	.clk(clk_clk),
	.d(\E_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[4]~q ),
	.prn(vcc));
defparam \M_iw[4] .is_wysiwyg = "true";
defparam \M_iw[4] .power_up = "low";

dffeas \M_iw[3] (
	.clk(clk_clk),
	.d(\E_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[3]~q ),
	.prn(vcc));
defparam \M_iw[3] .is_wysiwyg = "true";
defparam \M_iw[3] .power_up = "low";

dffeas \M_iw[2] (
	.clk(clk_clk),
	.d(\E_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[2]~q ),
	.prn(vcc));
defparam \M_iw[2] .is_wysiwyg = "true";
defparam \M_iw[2] .power_up = "low";

dffeas \M_iw[1] (
	.clk(clk_clk),
	.d(\E_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[1]~q ),
	.prn(vcc));
defparam \M_iw[1] .is_wysiwyg = "true";
defparam \M_iw[1] .power_up = "low";

cyclonev_lcell_comb \M_op_eret~1 (
	.dataa(!\M_iw[4]~q ),
	.datab(!\M_iw[3]~q ),
	.datac(!\M_iw[2]~q ),
	.datad(!\M_iw[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~1 .extended_lut = "off";
defparam \M_op_eret~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \M_op_eret~1 .shared_arith = "off";

cyclonev_lcell_comb \M_op_eret~2 (
	.dataa(!\M_iw[11]~q ),
	.datab(!\M_iw[5]~q ),
	.datac(!\M_iw[0]~q ),
	.datad(!\M_op_eret~0_combout ),
	.datae(!\M_op_eret~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~2 .extended_lut = "off";
defparam \M_op_eret~2 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \M_op_eret~2 .shared_arith = "off";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\A_status_reg_pie~q ),
	.datac(!\M_iw[6]~q ),
	.datad(!\M_iw[7]~q ),
	.datae(!\M_iw[8]~q ),
	.dataf(!\M_ctrl_wrctl_inst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~0 .lut_mask = 64'h7FF7F77FF77F7FF7;
defparam \A_status_reg_pie_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~1 (
	.dataa(!\M_iw[14]~q ),
	.datab(!\M_op_eret~2_combout ),
	.datac(!\A_estatus_reg_pie~q ),
	.datad(!\A_bstatus_reg_pie~q ),
	.datae(!\A_status_reg_pie_inst_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~1 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_status_reg_pie_inst_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~2 (
	.dataa(!\M_ctrl_break~q ),
	.datab(!\M_ctrl_exception~q ),
	.datac(!\M_ctrl_crst~q ),
	.datad(!\A_status_reg_pie_inst_nxt~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~2 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~2 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \A_status_reg_pie_inst_nxt~2 .shared_arith = "off";

dffeas A_status_reg_pie(
	.clk(clk_clk),
	.d(\A_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always138~0_combout ),
	.q(\A_status_reg_pie~q ),
	.prn(vcc));
defparam A_status_reg_pie.is_wysiwyg = "true";
defparam A_status_reg_pie.power_up = "low";

dffeas A_valid_wrctl_ienable(
	.clk(clk_clk),
	.d(\A_ienable_reg_irq0_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_valid_wrctl_ienable~q ),
	.prn(vcc));
defparam A_valid_wrctl_ienable.is_wysiwyg = "true";
defparam A_valid_wrctl_ienable.power_up = "low";

cyclonev_lcell_comb \norm_intr_req~0 (
	.dataa(!\A_status_reg_pie~q ),
	.datab(!\A_valid_wrctl_ienable~q ),
	.datac(!\A_ipending_reg_irq0~q ),
	.datad(!\A_ipending_reg_irq1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\norm_intr_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \norm_intr_req~0 .extended_lut = "off";
defparam \norm_intr_req~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \norm_intr_req~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[5]~1 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~1 .extended_lut = "off";
defparam \F_iw[5]~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[5]~1 .shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cyclonev_lcell_comb \Equal169~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal169~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal169~0 .extended_lut = "off";
defparam \Equal169~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \Equal169~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~2 .extended_lut = "off";
defparam \D_ctrl_late_result~2 .lut_mask = 64'hFDFFFFFFFFFDFFFF;
defparam \D_ctrl_late_result~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~0 .extended_lut = "off";
defparam \D_ctrl_late_result~0 .lut_mask = 64'hFFFFF7FBFFFFFFFF;
defparam \D_ctrl_late_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~1 (
	.dataa(!\Equal169~0_combout ),
	.datab(!\Equal152~6_combout ),
	.datac(!\D_ctrl_shift_rot~1_combout ),
	.datad(!\D_ctrl_late_result~2_combout ),
	.datae(!\D_ctrl_late_result~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~1 .extended_lut = "off";
defparam \D_ctrl_late_result~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_late_result~1 .shared_arith = "off";

dffeas E_ctrl_late_result(
	.clk(clk_clk),
	.d(\D_ctrl_late_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_late_result~q ),
	.prn(vcc));
defparam E_ctrl_late_result.is_wysiwyg = "true";
defparam E_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \D_data_depend~0 (
	.dataa(!\E_ctrl_late_result~q ),
	.datab(!\D_ctrl_a_not_src~q ),
	.datac(!\E_regnum_a_cmp_D~q ),
	.datad(!\D_ctrl_b_is_dst~q ),
	.datae(!\E_regnum_b_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~0 .extended_lut = "off";
defparam \D_data_depend~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_data_depend~0 .shared_arith = "off";

cyclonev_lcell_comb D_valid(
	.dataa(!\D_data_depend~0_combout ),
	.datab(!\D_data_depend~1_combout ),
	.datac(!\D_dep_stall~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_valid.extended_lut = "off";
defparam D_valid.lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam D_valid.shared_arith = "off";

dffeas E_valid_from_D(
	.clk(clk_clk),
	.d(\D_valid~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_valid_from_D~q ),
	.prn(vcc));
defparam E_valid_from_D.is_wysiwyg = "true";
defparam E_valid_from_D.power_up = "low";

cyclonev_lcell_comb \E_valid~0 (
	.dataa(!\E_valid_from_D~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~0 .extended_lut = "off";
defparam \E_valid~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \latched_oci_tb_hbreak_req_next~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!hbreak_enabled1),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\hbreak_req~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\latched_oci_tb_hbreak_req_next~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \latched_oci_tb_hbreak_req_next~0 .extended_lut = "off";
defparam \latched_oci_tb_hbreak_req_next~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \latched_oci_tb_hbreak_req_next~0 .shared_arith = "off";

dffeas latched_oci_tb_hbreak_req(
	.clk(clk_clk),
	.d(\latched_oci_tb_hbreak_req_next~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latched_oci_tb_hbreak_req~q ),
	.prn(vcc));
defparam latched_oci_tb_hbreak_req.is_wysiwyg = "true";
defparam latched_oci_tb_hbreak_req.power_up = "low";

cyclonev_lcell_comb \F_iw~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\latched_oci_tb_hbreak_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw~0 .extended_lut = "off";
defparam \F_iw~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[0]~9 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\norm_intr_req~0_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[0]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[0]~9 .extended_lut = "off";
defparam \F_iw[0]~9 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \F_iw[0]~9 .shared_arith = "off";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

dffeas \E_iw[0] (
	.clk(clk_clk),
	.d(\D_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[0]~q ),
	.prn(vcc));
defparam \E_iw[0] .is_wysiwyg = "true";
defparam \E_iw[0] .power_up = "low";

cyclonev_lcell_comb \E_ld_st_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add24~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_bus~0 .extended_lut = "off";
defparam \E_ld_st_bus~0 .lut_mask = 64'hF737FFFFFFFFFFFF;
defparam \E_ld_st_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_bypass(
	.clk(clk_clk),
	.d(\E_ld_st_bus~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_st_bypass.power_up = "low";

dffeas A_ctrl_ld_st_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_ld_st_bypass~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_st_bypass~q ),
	.prn(vcc));
defparam A_ctrl_ld_st_bypass.is_wysiwyg = "true";
defparam A_ctrl_ld_st_bypass.power_up = "low";

cyclonev_lcell_comb A_mem_bypass_pending(
	.dataa(!\A_ctrl_ld_st_bypass~q ),
	.datab(!\A_valid~q ),
	.datac(!\A_stall~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_bypass_pending~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_mem_bypass_pending.extended_lut = "off";
defparam A_mem_bypass_pending.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam A_mem_bypass_pending.shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[0]~0 (
	.dataa(!d_read1),
	.datab(!\A_dc_wb_rd_data_first~q ),
	.datac(!\A_dc_wb_active~q ),
	.datad(!\A_dc_want_fill~q ),
	.datae(!\A_dc_fill_has_started~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[0]~0 .extended_lut = "off";
defparam \d_address_offset_field[0]~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \d_address_offset_field[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add21~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_2),
	.datac(!d_address_offset_field_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add21~0 .extended_lut = "off";
defparam \Add21~0 .lut_mask = 64'h9696969696969696;
defparam \Add21~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[2]~0 (
	.dataa(!\av_addr_accepted~combout ),
	.datab(!\A_mem_bypass_pending~combout ),
	.datac(!\d_address_offset_field[0]~0_combout ),
	.datad(!\A_mem_baddr[4]~q ),
	.datae(!\Add21~0_combout ),
	.dataf(!\M_alu_result[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[2]~0 .extended_lut = "off";
defparam \d_address_offset_field_nxt[2]~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \d_address_offset_field_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[0]~1 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[0]~1 .extended_lut = "off";
defparam \d_address_offset_field[0]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \d_address_offset_field[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[0]~2 (
	.dataa(!rst1),
	.datab(!av_begintransfer),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(!\d_address_offset_field[0]~0_combout ),
	.dataf(!\d_address_offset_field[0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[0]~2 .extended_lut = "off";
defparam \d_address_offset_field[0]~2 .lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam \d_address_offset_field[0]~2 .shared_arith = "off";

cyclonev_lcell_comb A_dc_wb_update_av_writedata(
	.dataa(!rst1),
	.datab(!suppress_change_dest_id),
	.datac(!WideOr01),
	.datad(!\A_dc_wb_wr_starting~combout ),
	.datae(!\A_dc_wb_wr_active~q ),
	.dataf(!\A_dc_wr_data_cnt[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_update_av_writedata~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_update_av_writedata.extended_lut = "off";
defparam A_dc_wb_update_av_writedata.lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam A_dc_wb_update_av_writedata.shared_arith = "off";

dffeas \E_src2_reg[0] (
	.clk(clk_clk),
	.d(\D_src2_reg[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[0]~q ),
	.prn(vcc));
defparam \E_src2_reg[0] .is_wysiwyg = "true";
defparam \E_src2_reg[0] .power_up = "low";

dffeas \M_st_data[0] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[0]~q ),
	.prn(vcc));
defparam \M_st_data[0] .is_wysiwyg = "true";
defparam \M_st_data[0] .power_up = "low";

dffeas \A_st_data[0] (
	.clk(clk_clk),
	.d(\M_st_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[0]~q ),
	.prn(vcc));
defparam \A_st_data[0] .is_wysiwyg = "true";
defparam \A_st_data[0] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[0]~0 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\A_st_data[0]~q ),
	.datae(!\M_st_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[0]~0 .extended_lut = "off";
defparam \d_writedata_nxt[0]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_writedata[14]~0 (
	.dataa(!rst1),
	.datab(!suppress_change_dest_id),
	.datac(!WideOr01),
	.datad(!\A_dc_wb_wr_starting~combout ),
	.datae(!\A_dc_wb_wr_active~q ),
	.dataf(!\A_dc_wr_data_cnt[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata[14]~0 .extended_lut = "off";
defparam \d_writedata[14]~0 .lut_mask = 64'hFFFFFFFFFFFFFDFF;
defparam \d_writedata[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[0]~1 (
	.dataa(!d_address_offset_field_0),
	.datab(!\av_addr_accepted~combout ),
	.datac(!\A_mem_bypass_pending~combout ),
	.datad(!\d_address_offset_field[0]~0_combout ),
	.datae(!\A_mem_baddr[2]~q ),
	.dataf(!\M_alu_result[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[0]~1 .extended_lut = "off";
defparam \d_address_offset_field_nxt[0]~1 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \d_address_offset_field_nxt[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_st_bypass_delayed~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\M_ctrl_st_bypass~q ),
	.datac(!\M_valid_from_E~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_delayed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_st_bypass_delayed~0 .extended_lut = "off";
defparam \A_st_bypass_delayed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_st_bypass_delayed~0 .shared_arith = "off";

dffeas A_st_bypass_delayed(
	.clk(clk_clk),
	.d(\A_st_bypass_delayed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_bypass_delayed~q ),
	.prn(vcc));
defparam A_st_bypass_delayed.is_wysiwyg = "true";
defparam A_st_bypass_delayed.power_up = "low";

cyclonev_lcell_comb \A_st_bypass_delayed_started~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_st_bypass_delayed~q ),
	.datac(!\A_st_bypass_delayed_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_delayed_started~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_st_bypass_delayed_started~0 .extended_lut = "off";
defparam \A_st_bypass_delayed_started~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_st_bypass_delayed_started~0 .shared_arith = "off";

dffeas A_st_bypass_delayed_started(
	.clk(clk_clk),
	.d(\A_st_bypass_delayed_started~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_st_bypass_delayed_started~q ),
	.prn(vcc));
defparam A_st_bypass_delayed_started.is_wysiwyg = "true";
defparam A_st_bypass_delayed_started.power_up = "low";

cyclonev_lcell_comb \d_write_nxt~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_st_bypass_delayed~q ),
	.datac(!\A_st_bypass_delayed_started~q ),
	.datad(!\M_ctrl_st_bypass~q ),
	.datae(!\always138~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~0 .extended_lut = "off";
defparam \d_write_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \d_write_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \d_write_nxt~1 (
	.dataa(!d_write1),
	.datab(!av_waitrequest),
	.datac(!\A_dc_wb_wr_starting~combout ),
	.datad(!\A_dc_wr_data_cnt[3]~q ),
	.datae(!\d_write_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~1 .extended_lut = "off";
defparam \d_write_nxt~1 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \d_write_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb A_dc_wb_wr_want_dmaster(
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_want_dmaster~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_wr_want_dmaster.extended_lut = "off";
defparam A_dc_wb_wr_want_dmaster.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam A_dc_wb_wr_want_dmaster.shared_arith = "off";

dffeas \A_dc_wb_line[0] (
	.clk(clk_clk),
	.d(\A_mem_baddr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[0] .is_wysiwyg = "true";
defparam \A_dc_wb_line[0] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt~0 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(!\A_dc_fill_active~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt~0 .extended_lut = "off";
defparam \d_address_tag_field_nxt~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \d_address_tag_field_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_line_field_nxt[0]~0 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\A_dc_wb_line[0]~q ),
	.datac(!\d_address_tag_field_nxt~0_combout ),
	.datad(!\A_mem_baddr[5]~q ),
	.datae(!\M_alu_result[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[0]~0 .extended_lut = "off";
defparam \d_address_line_field_nxt[0]~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \d_address_line_field_nxt[0]~0 .shared_arith = "off";

dffeas \A_dc_actual_tag[1] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[1]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[1] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[1] .power_up = "low";

dffeas \A_dc_wb_tag[1] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[1] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[1] .power_up = "low";

dffeas \A_mem_baddr[12] (
	.clk(clk_clk),
	.d(\M_alu_result[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[12]~q ),
	.prn(vcc));
defparam \A_mem_baddr[12] .is_wysiwyg = "true";
defparam \A_mem_baddr[12] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[1]~1 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[1]~q ),
	.datad(!\A_mem_baddr[12]~q ),
	.datae(!\M_alu_result[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[1]~1 .extended_lut = "off";
defparam \d_address_tag_field_nxt[1]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[1]~1 .shared_arith = "off";

dffeas \A_dc_actual_tag[0] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[0]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[0] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[0] .power_up = "low";

dffeas \A_dc_wb_tag[0] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[0] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[0] .power_up = "low";

dffeas \A_mem_baddr[11] (
	.clk(clk_clk),
	.d(\M_alu_result[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[11]~q ),
	.prn(vcc));
defparam \A_mem_baddr[11] .is_wysiwyg = "true";
defparam \A_mem_baddr[11] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[0]~2 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[0]~q ),
	.datad(!\A_mem_baddr[11]~q ),
	.datae(!\M_alu_result[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[0]~2 .extended_lut = "off";
defparam \d_address_tag_field_nxt[0]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[0]~2 .shared_arith = "off";

dffeas \A_dc_wb_line[5] (
	.clk(clk_clk),
	.d(\A_mem_baddr[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[5]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[5] .is_wysiwyg = "true";
defparam \A_dc_wb_line[5] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[5]~1 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[5]~q ),
	.datad(!\A_mem_baddr[10]~q ),
	.datae(!\M_alu_result[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[5]~1 .extended_lut = "off";
defparam \d_address_line_field_nxt[5]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[5]~1 .shared_arith = "off";

dffeas \A_dc_wb_line[4] (
	.clk(clk_clk),
	.d(\A_mem_baddr[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[4]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[4] .is_wysiwyg = "true";
defparam \A_dc_wb_line[4] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[4]~2 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[4]~q ),
	.datad(!\A_mem_baddr[9]~q ),
	.datae(!\M_alu_result[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[4]~2 .extended_lut = "off";
defparam \d_address_line_field_nxt[4]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[4]~2 .shared_arith = "off";

dffeas \A_dc_wb_line[3] (
	.clk(clk_clk),
	.d(\A_mem_baddr[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[3]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[3] .is_wysiwyg = "true";
defparam \A_dc_wb_line[3] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[3]~3 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[3]~q ),
	.datad(!\A_mem_baddr[8]~q ),
	.datae(!\M_alu_result[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[3]~3 .extended_lut = "off";
defparam \d_address_line_field_nxt[3]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[3]~3 .shared_arith = "off";

dffeas \A_dc_wb_line[2] (
	.clk(clk_clk),
	.d(\A_mem_baddr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[2] .is_wysiwyg = "true";
defparam \A_dc_wb_line[2] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[2]~4 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[2]~q ),
	.datad(!\A_mem_baddr[7]~q ),
	.datae(!\M_alu_result[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[2]~4 .extended_lut = "off";
defparam \d_address_line_field_nxt[2]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[2]~4 .shared_arith = "off";

dffeas \A_dc_wb_line[1] (
	.clk(clk_clk),
	.d(\A_mem_baddr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[1] .is_wysiwyg = "true";
defparam \A_dc_wb_line[1] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[1]~5 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[1]~q ),
	.datad(!\A_mem_baddr[6]~q ),
	.datae(!\M_alu_result[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[1]~5 .extended_lut = "off";
defparam \d_address_line_field_nxt[1]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[1]~5 .shared_arith = "off";

dffeas \A_dc_actual_tag[5] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[5]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[5] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[5] .power_up = "low";

dffeas \A_dc_wb_tag[5] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[5]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[5] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[5] .power_up = "low";

dffeas \A_mem_baddr[16] (
	.clk(clk_clk),
	.d(\M_alu_result[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[16]~q ),
	.prn(vcc));
defparam \A_mem_baddr[16] .is_wysiwyg = "true";
defparam \A_mem_baddr[16] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[5]~3 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[5]~q ),
	.datad(!\A_mem_baddr[16]~q ),
	.datae(!\M_alu_result[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[5]~3 .extended_lut = "off";
defparam \d_address_tag_field_nxt[5]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[5]~3 .shared_arith = "off";

dffeas \A_dc_actual_tag[4] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[4]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[4] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[4] .power_up = "low";

dffeas \A_dc_wb_tag[4] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[4]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[4] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[4] .power_up = "low";

dffeas \A_mem_baddr[15] (
	.clk(clk_clk),
	.d(\M_alu_result[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[15]~q ),
	.prn(vcc));
defparam \A_mem_baddr[15] .is_wysiwyg = "true";
defparam \A_mem_baddr[15] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[4]~4 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[4]~q ),
	.datad(!\A_mem_baddr[15]~q ),
	.datae(!\M_alu_result[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[4]~4 .extended_lut = "off";
defparam \d_address_tag_field_nxt[4]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[4]~4 .shared_arith = "off";

dffeas \A_dc_actual_tag[3] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[3]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[3] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[3] .power_up = "low";

dffeas \A_dc_wb_tag[3] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[3]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[3] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[3] .power_up = "low";

dffeas \A_mem_baddr[14] (
	.clk(clk_clk),
	.d(\M_alu_result[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[14]~q ),
	.prn(vcc));
defparam \A_mem_baddr[14] .is_wysiwyg = "true";
defparam \A_mem_baddr[14] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[3]~5 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[3]~q ),
	.datad(!\A_mem_baddr[14]~q ),
	.datae(!\M_alu_result[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[3]~5 .extended_lut = "off";
defparam \d_address_tag_field_nxt[3]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[3]~5 .shared_arith = "off";

dffeas \A_dc_actual_tag[2] (
	.clk(clk_clk),
	.d(\Qsys_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[2]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[2] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[2] .power_up = "low";

dffeas \A_dc_wb_tag[2] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[2] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[2] .power_up = "low";

dffeas \A_mem_baddr[13] (
	.clk(clk_clk),
	.d(\M_alu_result[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[13]~q ),
	.prn(vcc));
defparam \A_mem_baddr[13] .is_wysiwyg = "true";
defparam \A_mem_baddr[13] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[2]~6 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[2]~q ),
	.datad(!\A_mem_baddr[13]~q ),
	.datae(!\M_alu_result[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[2]~6 .extended_lut = "off";
defparam \d_address_tag_field_nxt[2]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[1]~2 (
	.dataa(!d_address_offset_field_0),
	.datab(!d_address_offset_field_1),
	.datac(!\A_mem_baddr[3]~q ),
	.datad(!\d_address_offset_field[0]~0_combout ),
	.datae(!\A_mem_bypass_pending~combout ),
	.dataf(!\av_addr_accepted~combout ),
	.datag(!\M_alu_result[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[1]~2 .extended_lut = "on";
defparam \d_address_offset_field_nxt[1]~2 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \d_address_offset_field_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_ld_bypass_delayed~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_ld_bypass~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_delayed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ld_bypass_delayed~0 .extended_lut = "off";
defparam \A_ld_bypass_delayed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_ld_bypass_delayed~0 .shared_arith = "off";

dffeas A_ld_bypass_delayed(
	.clk(clk_clk),
	.d(\A_ld_bypass_delayed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_bypass_delayed~q ),
	.prn(vcc));
defparam A_ld_bypass_delayed.is_wysiwyg = "true";
defparam A_ld_bypass_delayed.power_up = "low";

cyclonev_lcell_comb \A_ld_bypass_delayed_started~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_ld_bypass_delayed~q ),
	.datac(!\A_ld_bypass_delayed_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_delayed_started~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ld_bypass_delayed_started~0 .extended_lut = "off";
defparam \A_ld_bypass_delayed_started~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_ld_bypass_delayed_started~0 .shared_arith = "off";

dffeas A_ld_bypass_delayed_started(
	.clk(clk_clk),
	.d(\A_ld_bypass_delayed_started~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_ld_bypass_delayed_started~q ),
	.prn(vcc));
defparam A_ld_bypass_delayed_started.is_wysiwyg = "true";
defparam A_ld_bypass_delayed_started.power_up = "low";

cyclonev_lcell_comb \d_read_nxt~0 (
	.dataa(!\A_dc_want_fill~q ),
	.datab(!\A_dc_fill_has_started~q ),
	.datac(!\A_ld_bypass_delayed~q ),
	.datad(!\A_ld_bypass_delayed_started~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~0 .extended_lut = "off";
defparam \d_read_nxt~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \d_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \d_read_nxt~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\always138~0_combout ),
	.datac(!\M_ctrl_ld_bypass~q ),
	.datad(!\d_read_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~1 .extended_lut = "off";
defparam \d_read_nxt~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \d_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[0]~3 (
	.dataa(!d_read1),
	.datab(!av_waitrequest),
	.datac(!\A_dc_fill_starting~0_combout ),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt[0]~0 (
	.dataa(!rst1),
	.datab(!d_read1),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr01),
	.datae(!\A_dc_fill_starting~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt[0]~0 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt[0]~0 .lut_mask = 64'hFFFFFFFFFFF7FFFF;
defparam \A_dc_rd_addr_cnt[0]~0 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[0]~0_combout ),
	.q(\A_dc_rd_addr_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[1]~2 (
	.dataa(!d_read1),
	.datab(!av_waitrequest),
	.datac(!\A_dc_rd_addr_cnt[1]~q ),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[0]~0_combout ),
	.q(\A_dc_rd_addr_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[2]~1 (
	.dataa(!d_read1),
	.datab(!av_waitrequest),
	.datac(!\A_dc_rd_addr_cnt[2]~q ),
	.datad(!\A_dc_rd_addr_cnt[1]~q ),
	.datae(!\A_dc_rd_addr_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .lut_mask = 64'hF77F7FF7F77F7FF7;
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[0]~0_combout ),
	.q(\A_dc_rd_addr_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add22~0 (
	.dataa(!\A_dc_rd_addr_cnt[3]~q ),
	.datab(!\A_dc_rd_addr_cnt[2]~q ),
	.datac(!\A_dc_rd_addr_cnt[1]~q ),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add22~0 .extended_lut = "off";
defparam \Add22~0 .lut_mask = 64'h6996699669966996;
defparam \Add22~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[3]~0 (
	.dataa(!d_read1),
	.datab(!av_waitrequest),
	.datac(!\A_dc_fill_starting~0_combout ),
	.datad(!\Add22~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .lut_mask = 64'hF6FFF6FFF6FFF6FF;
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[0]~0_combout ),
	.q(\A_dc_rd_addr_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[3] .power_up = "low";

cyclonev_lcell_comb \d_read_nxt~2 (
	.dataa(!d_read1),
	.datab(!av_waitrequest),
	.datac(!\d_read_nxt~1_combout ),
	.datad(!\A_dc_rd_addr_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~2 .extended_lut = "off";
defparam \d_read_nxt~2 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \d_read_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~0 (
	.dataa(!ic_fill_line_5),
	.datab(!\F_pc[7]~q ),
	.datac(!ic_fill_line_4),
	.datad(!\F_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~0 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~0 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~1 (
	.dataa(!\F_pc[4]~q ),
	.datab(!ic_fill_line_1),
	.datac(!\F_pc[5]~q ),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~1 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~2 (
	.dataa(!ic_fill_tag_1),
	.datab(!ic_fill_tag_0),
	.datac(!\F_pc[10]~q ),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~2 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~2 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~3 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!\F_pc[14]~q ),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~3 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~3 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~3 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~4 (
	.dataa(!ic_fill_tag_2),
	.datab(!\F_pc[12]~q ),
	.datac(!\F_pc[3]~q ),
	.datad(!ic_fill_line_0),
	.datae(!\F_ic_fill_same_tag_line~2_combout ),
	.dataf(!\F_ic_fill_same_tag_line~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~4 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \F_ic_fill_same_tag_line~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~5 (
	.dataa(!\F_pc[6]~q ),
	.datab(!ic_fill_line_3),
	.datac(!\F_ic_fill_same_tag_line~1_combout ),
	.datad(!\F_ic_fill_same_tag_line~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~5 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \F_ic_fill_same_tag_line~5 .shared_arith = "off";

cyclonev_lcell_comb F_ic_fill_same_tag_line(
	.dataa(!ic_fill_line_6),
	.datab(!\F_pc[9]~q ),
	.datac(!\F_ic_fill_same_tag_line~0_combout ),
	.datad(!\F_ic_fill_same_tag_line~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ic_fill_same_tag_line.extended_lut = "off";
defparam F_ic_fill_same_tag_line.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam F_ic_fill_same_tag_line.shared_arith = "off";

dffeas D_ic_fill_same_tag_line(
	.clk(clk_clk),
	.d(\F_ic_fill_same_tag_line~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ic_fill_same_tag_line~q ),
	.prn(vcc));
defparam D_ic_fill_same_tag_line.is_wysiwyg = "true";
defparam D_ic_fill_same_tag_line.power_up = "low";

cyclonev_lcell_comb \E_ctrl_invalidate_i~0 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_iw[11]~q ),
	.datac(!\E_iw[16]~q ),
	.datad(!\E_iw[15]~q ),
	.datae(!\E_iw[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~0 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~0 .lut_mask = 64'h9669699696696996;
defparam \E_ctrl_invalidate_i~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_invalidate_i~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\Equal207~0_combout ),
	.datac(!\E_ctrl_invalidate_i~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~1 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_invalidate_i~1 .shared_arith = "off";

dffeas M_ctrl_invalidate_i(
	.clk(clk_clk),
	.d(\E_ctrl_invalidate_i~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_invalidate_i~q ),
	.prn(vcc));
defparam M_ctrl_invalidate_i.is_wysiwyg = "true";
defparam M_ctrl_invalidate_i.power_up = "low";

cyclonev_lcell_comb \ic_tag_clr_valid_bits_nxt~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_invalidate_i~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \ic_tag_clr_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_prevent_refill_nxt(
	.dataa(!\ic_fill_prevent_refill~q ),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_prevent_refill_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_prevent_refill_nxt.extended_lut = "off";
defparam ic_fill_prevent_refill_nxt.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam ic_fill_prevent_refill_nxt.shared_arith = "off";

dffeas ic_fill_prevent_refill(
	.clk(clk_clk),
	.d(\ic_fill_prevent_refill_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_prevent_refill~q ),
	.prn(vcc));
defparam ic_fill_prevent_refill.is_wysiwyg = "true";
defparam ic_fill_prevent_refill.power_up = "low";

dffeas \ic_fill_initial_offset[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[2] .power_up = "low";

dffeas D_ic_fill_starting_d1(
	.clk(clk_clk),
	.d(\D_ic_fill_starting~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_ic_fill_starting_d1~q ),
	.prn(vcc));
defparam D_ic_fill_starting_d1.is_wysiwyg = "true";
defparam D_ic_fill_starting_d1.power_up = "low";

dffeas \ic_fill_initial_offset[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[0]~1 (
	.dataa(!\ic_fill_initial_offset[0]~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(!\ic_fill_dp_offset[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \ic_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

dffeas i_readdatavalid_d1(
	.clk(clk_clk),
	.d(WideOr11),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdatavalid_d1~q ),
	.prn(vcc));
defparam i_readdatavalid_d1.is_wysiwyg = "true";
defparam i_readdatavalid_d1.power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_en~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_en~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_en~0 .lut_mask = 64'h7777777777777777;
defparam \ic_fill_dp_offset_en~0 .shared_arith = "off";

dffeas \ic_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[0] .power_up = "low";

dffeas \ic_fill_initial_offset[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[1]~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_initial_offset[1]~q ),
	.datad(!\ic_fill_dp_offset[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[1]~2 .lut_mask = 64'h9F6F9F6F9F6F9F6F;
defparam \ic_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[1] .power_up = "low";

dffeas \ic_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[2]~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_dp_offset[1]~q ),
	.datad(!\ic_fill_initial_offset[2]~q ),
	.datae(!\ic_fill_dp_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[2]~0 .lut_mask = 64'h69FF96FF69FF96FF;
defparam \ic_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_fill_initial_offset[0]~q ),
	.datac(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datad(!\ic_fill_initial_offset[1]~q ),
	.datae(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~0 .extended_lut = "off";
defparam \ic_fill_active_nxt~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_active_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~1 (
	.dataa(!\ic_fill_active~q ),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_fill_initial_offset[2]~q ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_active_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~1 .extended_lut = "off";
defparam \ic_fill_active_nxt~1 .lut_mask = 64'hFFFF7FF7FFFF7FF7;
defparam \ic_fill_active_nxt~1 .shared_arith = "off";

dffeas ic_fill_active(
	.clk(clk_clk),
	.d(\ic_fill_active_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_active~q ),
	.prn(vcc));
defparam ic_fill_active.is_wysiwyg = "true";
defparam ic_fill_active.power_up = "low";

cyclonev_lcell_comb \D_ic_fill_starting~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_ic_fill_same_tag_line~q ),
	.datac(!\ic_fill_prevent_refill~q ),
	.datad(!\ic_fill_active~q ),
	.datae(!\D_iw_valid~q ),
	.dataf(!\D_kill~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ic_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ic_fill_starting~0 .extended_lut = "off";
defparam \D_ic_fill_starting~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \D_ic_fill_starting~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[0]~3 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[0]~3 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[0]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \ic_fill_ap_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_cnt[3]~0 (
	.dataa(!save_dest_id),
	.datab(!WideOr0),
	.datac(!\D_ic_fill_starting~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt[3]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt[3]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ic_fill_ap_cnt[3]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(\ic_fill_ap_cnt[0]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[1]~q ),
	.datac(!\ic_fill_ap_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \ic_fill_ap_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(\ic_fill_ap_cnt[1]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[2]~q ),
	.datac(!\ic_fill_ap_cnt[1]~q ),
	.datad(!\ic_fill_ap_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \ic_fill_ap_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(\ic_fill_ap_cnt[2]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[3]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[3]~q ),
	.datac(!\ic_fill_ap_cnt[2]~q ),
	.datad(!\ic_fill_ap_cnt[1]~q ),
	.datae(!\ic_fill_ap_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[3]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[3]~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_ap_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[3] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[3]~0_combout ),
	.q(\ic_fill_ap_cnt[3]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[3] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[3] .power_up = "low";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!rst1),
	.datab(!has_pending_responses),
	.datac(!suppress_change_dest_id1),
	.datad(!\ic_fill_active~q ),
	.datae(!\ic_fill_ap_cnt[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~1 (
	.dataa(!i_read1),
	.datab(!WideOr0),
	.datac(!\D_ic_fill_starting~0_combout ),
	.datad(!\i_read_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~1 .extended_lut = "off";
defparam \i_read_nxt~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \i_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~0 (
	.dataa(!ic_fill_line_6),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\D_pc[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~0 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~0 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\M_ctrl_break~q ),
	.datac(!\M_iw[14]~q ),
	.datad(!\M_op_eret~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~0 .extended_lut = "off";
defparam \hbreak_enabled~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \hbreak_enabled~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~1 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_5),
	.datac(!\D_pc[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~1 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~1 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~2 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_4),
	.datac(!\D_pc[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~2 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~2 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~3 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_3),
	.datac(!\D_pc[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~3 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~3 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~4 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_1),
	.datac(!\D_pc[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~4 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~4 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~5 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_2),
	.datac(!\D_pc[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~5 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~5 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~6 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_0),
	.datac(!\D_pc[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~6 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~6 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~6 .shared_arith = "off";

dffeas \E_src2_reg[7] (
	.clk(clk_clk),
	.d(\D_src2_reg[7]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[7]~q ),
	.prn(vcc));
defparam \E_src2_reg[7] .is_wysiwyg = "true";
defparam \E_src2_reg[7] .power_up = "low";

dffeas \M_st_data[7] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[7]~q ),
	.prn(vcc));
defparam \M_st_data[7] .is_wysiwyg = "true";
defparam \M_st_data[7] .power_up = "low";

dffeas \A_st_data[7] (
	.clk(clk_clk),
	.d(\M_st_data[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[7]~q ),
	.prn(vcc));
defparam \A_st_data[7] .is_wysiwyg = "true";
defparam \A_st_data[7] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[7]~1 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[7]~q ),
	.datad(!\A_st_data[7]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[7]~1 .extended_lut = "off";
defparam \d_writedata_nxt[7]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[0]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!\D_pc[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[0]~0 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[0]~0 .lut_mask = 64'h8D8D8D8D8D8D8D8D;
defparam \ic_fill_ap_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!ic_fill_ap_offset_2),
	.datad(!ic_fill_ap_offset_1),
	.datae(!\D_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[2]~1 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \ic_fill_ap_offset_nxt[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!ic_fill_ap_offset_1),
	.datad(!\D_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[1]~2 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \ic_fill_ap_offset_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add24~69_sumout ),
	.datad(!\Add24~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \E_mem_byte_en~0 .shared_arith = "off";

dffeas \M_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[0]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[0] .is_wysiwyg = "true";
defparam \M_mem_byte_en[0] .power_up = "low";

dffeas \A_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[0]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[0] .is_wysiwyg = "true";
defparam \A_mem_byte_en[0] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[0]~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\A_dc_wb_wr_want_dmaster~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[0]~0 .extended_lut = "off";
defparam \d_byteenable_nxt[0]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \d_byteenable_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_byteenable_nxt[0]~1 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\M_mem_byte_en[0]~q ),
	.datac(!\A_mem_byte_en[0]~q ),
	.datad(!\d_byteenable_nxt[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[0]~1 .extended_lut = "off";
defparam \d_byteenable_nxt[0]~1 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \d_byteenable_nxt[0]~1 .shared_arith = "off";

dffeas \E_src2_reg[3] (
	.clk(clk_clk),
	.d(\D_src2_reg[3]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[3]~q ),
	.prn(vcc));
defparam \E_src2_reg[3] .is_wysiwyg = "true";
defparam \E_src2_reg[3] .power_up = "low";

dffeas \M_st_data[3] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[3]~q ),
	.prn(vcc));
defparam \M_st_data[3] .is_wysiwyg = "true";
defparam \M_st_data[3] .power_up = "low";

dffeas \A_st_data[3] (
	.clk(clk_clk),
	.d(\M_st_data[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[3]~q ),
	.prn(vcc));
defparam \A_st_data[3] .is_wysiwyg = "true";
defparam \A_st_data[3] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[3]~2 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[3]~q ),
	.datad(!\A_st_data[3]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[3]~2 .extended_lut = "off";
defparam \d_writedata_nxt[3]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[3]~2 .shared_arith = "off";

dffeas \E_src2_reg[1] (
	.clk(clk_clk),
	.d(\D_src2_reg[1]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[1]~q ),
	.prn(vcc));
defparam \E_src2_reg[1] .is_wysiwyg = "true";
defparam \E_src2_reg[1] .power_up = "low";

dffeas \M_st_data[1] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[1]~q ),
	.prn(vcc));
defparam \M_st_data[1] .is_wysiwyg = "true";
defparam \M_st_data[1] .power_up = "low";

dffeas \A_st_data[1] (
	.clk(clk_clk),
	.d(\M_st_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[1]~q ),
	.prn(vcc));
defparam \A_st_data[1] .is_wysiwyg = "true";
defparam \A_st_data[1] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[1]~3 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[1]~q ),
	.datad(!\A_st_data[1]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[1]~3 .extended_lut = "off";
defparam \d_writedata_nxt[1]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[1]~3 .shared_arith = "off";

dffeas \E_src2_reg[4] (
	.clk(clk_clk),
	.d(\D_src2_reg[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[4]~q ),
	.prn(vcc));
defparam \E_src2_reg[4] .is_wysiwyg = "true";
defparam \E_src2_reg[4] .power_up = "low";

dffeas \M_st_data[4] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[4]~q ),
	.prn(vcc));
defparam \M_st_data[4] .is_wysiwyg = "true";
defparam \M_st_data[4] .power_up = "low";

dffeas \A_st_data[4] (
	.clk(clk_clk),
	.d(\M_st_data[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[4]~q ),
	.prn(vcc));
defparam \A_st_data[4] .is_wysiwyg = "true";
defparam \A_st_data[4] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[4]~4 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[4]~q ),
	.datad(!\A_st_data[4]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[4]~4 .extended_lut = "off";
defparam \d_writedata_nxt[4]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[4]~4 .shared_arith = "off";

dffeas \E_src2_reg[20] (
	.clk(clk_clk),
	.d(\D_src2_reg[20]~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[20]~q ),
	.prn(vcc));
defparam \E_src2_reg[20] .is_wysiwyg = "true";
defparam \E_src2_reg[20] .power_up = "low";

dffeas \M_st_data[20] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[20]~q ),
	.prn(vcc));
defparam \M_st_data[20] .is_wysiwyg = "true";
defparam \M_st_data[20] .power_up = "low";

dffeas \A_st_data[20] (
	.clk(clk_clk),
	.d(\M_st_data[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[20]~q ),
	.prn(vcc));
defparam \A_st_data[20] .is_wysiwyg = "true";
defparam \A_st_data[20] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[20]~5 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[20]~q ),
	.datad(!\A_st_data[20]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[20]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[20]~5 .extended_lut = "off";
defparam \d_writedata_nxt[20]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[20]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add24~69_sumout ),
	.datad(!\Add24~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~1 .extended_lut = "off";
defparam \E_mem_byte_en[2]~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_mem_byte_en[2]~1 .shared_arith = "off";

dffeas \M_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[2]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[2] .is_wysiwyg = "true";
defparam \M_mem_byte_en[2] .power_up = "low";

dffeas \A_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[2]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[2] .is_wysiwyg = "true";
defparam \A_mem_byte_en[2] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[2]~2 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\M_mem_byte_en[2]~q ),
	.datac(!\A_mem_byte_en[2]~q ),
	.datad(!\d_byteenable_nxt[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[2]~2 .extended_lut = "off";
defparam \d_byteenable_nxt[2]~2 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \d_byteenable_nxt[2]~2 .shared_arith = "off";

dffeas \E_src2_reg[12] (
	.clk(clk_clk),
	.d(\D_src2_reg[12]~127_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[12]~q ),
	.prn(vcc));
defparam \E_src2_reg[12] .is_wysiwyg = "true";
defparam \E_src2_reg[12] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7777777777777777;
defparam \Equal0~0 .shared_arith = "off";

dffeas \M_st_data[12] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[12]~q ),
	.prn(vcc));
defparam \M_st_data[12] .is_wysiwyg = "true";
defparam \M_st_data[12] .power_up = "low";

dffeas \A_st_data[12] (
	.clk(clk_clk),
	.d(\M_st_data[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[12]~q ),
	.prn(vcc));
defparam \A_st_data[12] .is_wysiwyg = "true";
defparam \A_st_data[12] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[12]~6 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[12]~q ),
	.datad(!\A_st_data[12]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[12]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[12]~6 .extended_lut = "off";
defparam \d_writedata_nxt[12]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[12]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[1]~2 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add24~69_sumout ),
	.datad(!\Add24~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~2 .extended_lut = "off";
defparam \E_mem_byte_en[1]~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \E_mem_byte_en[1]~2 .shared_arith = "off";

dffeas \M_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[1]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[1] .is_wysiwyg = "true";
defparam \M_mem_byte_en[1] .power_up = "low";

dffeas \A_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[1]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[1] .is_wysiwyg = "true";
defparam \A_mem_byte_en[1] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[1]~3 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\A_mem_byte_en[1]~q ),
	.datad(!\d_byteenable_nxt[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[1]~3 .extended_lut = "off";
defparam \d_byteenable_nxt[1]~3 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \d_byteenable_nxt[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~62 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~62 .extended_lut = "off";
defparam \D_src2_reg[28]~62 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[28]~62 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~63 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~18_combout ),
	.datad(!\Add24~85_sumout ),
	.datae(!\D_src2_reg[28]~62_combout ),
	.dataf(!\D_src2_reg[28]~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~63 .extended_lut = "off";
defparam \D_src2_reg[28]~63 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[28]~63 .shared_arith = "off";

dffeas \E_src2_reg[28] (
	.clk(clk_clk),
	.d(\D_src2_reg[28]~63_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[28]~q ),
	.prn(vcc));
defparam \E_src2_reg[28] .is_wysiwyg = "true";
defparam \E_src2_reg[28] .power_up = "low";

cyclonev_lcell_comb \E_st_data[28]~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[4]~q ),
	.datad(!\E_src2_reg[12]~q ),
	.datae(!\E_src2_reg[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~0 .extended_lut = "off";
defparam \E_st_data[28]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[28]~0 .shared_arith = "off";

dffeas \M_st_data[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[28]~q ),
	.prn(vcc));
defparam \M_st_data[28] .is_wysiwyg = "true";
defparam \M_st_data[28] .power_up = "low";

dffeas \A_st_data[28] (
	.clk(clk_clk),
	.d(\M_st_data[28]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[28]~q ),
	.prn(vcc));
defparam \A_st_data[28] .is_wysiwyg = "true";
defparam \A_st_data[28] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[28]~7 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[28]~q ),
	.datad(!\A_st_data[28]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[28]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[28]~7 .extended_lut = "off";
defparam \d_writedata_nxt[28]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[28]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add24~69_sumout ),
	.datad(!\Add24~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~3 .extended_lut = "off";
defparam \E_mem_byte_en[3]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_mem_byte_en[3]~3 .shared_arith = "off";

dffeas \M_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[3]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[3] .is_wysiwyg = "true";
defparam \M_mem_byte_en[3] .power_up = "low";

dffeas \A_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[3]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[3] .is_wysiwyg = "true";
defparam \A_mem_byte_en[3] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[3]~4 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\A_mem_byte_en[3]~q ),
	.datad(!\d_byteenable_nxt[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[3]~4 .extended_lut = "off";
defparam \d_byteenable_nxt[3]~4 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \d_byteenable_nxt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[16]~64 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[16]~23_combout ),
	.datad(!\E_alu_result[16]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~64 .extended_lut = "off";
defparam \D_src2_reg[16]~64 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[16]~64 .shared_arith = "off";

dffeas \E_src2_reg[16] (
	.clk(clk_clk),
	.d(\D_src2_reg[16]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[16]~q ),
	.prn(vcc));
defparam \E_src2_reg[16] .is_wysiwyg = "true";
defparam \E_src2_reg[16] .power_up = "low";

dffeas \M_st_data[16] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[16]~q ),
	.prn(vcc));
defparam \M_st_data[16] .is_wysiwyg = "true";
defparam \M_st_data[16] .power_up = "low";

dffeas \A_st_data[16] (
	.clk(clk_clk),
	.d(\M_st_data[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[16]~q ),
	.prn(vcc));
defparam \A_st_data[16] .is_wysiwyg = "true";
defparam \A_st_data[16] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[16]~8 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[16]~q ),
	.datad(!\A_st_data[16]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[16]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[16]~8 .extended_lut = "off";
defparam \d_writedata_nxt[16]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[16]~8 .shared_arith = "off";

dffeas \E_src2_reg[8] (
	.clk(clk_clk),
	.d(\D_src2_reg[8]~111_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[8]~q ),
	.prn(vcc));
defparam \E_src2_reg[8] .is_wysiwyg = "true";
defparam \E_src2_reg[8] .power_up = "low";

dffeas \M_st_data[8] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[8]~q ),
	.prn(vcc));
defparam \M_st_data[8] .is_wysiwyg = "true";
defparam \M_st_data[8] .power_up = "low";

dffeas \A_st_data[8] (
	.clk(clk_clk),
	.d(\M_st_data[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[8]~q ),
	.prn(vcc));
defparam \A_st_data[8] .is_wysiwyg = "true";
defparam \A_st_data[8] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[8]~9 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[8]~q ),
	.datad(!\A_st_data[8]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[8]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[8]~9 .extended_lut = "off";
defparam \d_writedata_nxt[8]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[8]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~65 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~65 .extended_lut = "off";
defparam \D_src2_reg[24]~65 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[24]~65 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~66 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~29_combout ),
	.datad(!\Add24~125_sumout ),
	.datae(!\D_src2_reg[24]~65_combout ),
	.dataf(!\D_src2_reg[24]~57_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~66 .extended_lut = "off";
defparam \D_src2_reg[24]~66 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[24]~66 .shared_arith = "off";

dffeas \E_src2_reg[24] (
	.clk(clk_clk),
	.d(\D_src2_reg[24]~66_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[24]~q ),
	.prn(vcc));
defparam \E_src2_reg[24] .is_wysiwyg = "true";
defparam \E_src2_reg[24] .power_up = "low";

cyclonev_lcell_comb \E_st_data[24]~1 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[0]~q ),
	.datad(!\E_src2_reg[8]~q ),
	.datae(!\E_src2_reg[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~1 .extended_lut = "off";
defparam \E_st_data[24]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[24]~1 .shared_arith = "off";

dffeas \M_st_data[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[24]~q ),
	.prn(vcc));
defparam \M_st_data[24] .is_wysiwyg = "true";
defparam \M_st_data[24] .power_up = "low";

dffeas \A_st_data[24] (
	.clk(clk_clk),
	.d(\M_st_data[24]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[24]~q ),
	.prn(vcc));
defparam \A_st_data[24] .is_wysiwyg = "true";
defparam \A_st_data[24] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[24]~10 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[24]~q ),
	.datad(!\A_st_data[24]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[24]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[24]~10 .extended_lut = "off";
defparam \d_writedata_nxt[24]~10 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[24]~10 .shared_arith = "off";

dffeas \E_src2_reg[2] (
	.clk(clk_clk),
	.d(\D_src2_reg[2]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[2]~q ),
	.prn(vcc));
defparam \E_src2_reg[2] .is_wysiwyg = "true";
defparam \E_src2_reg[2] .power_up = "low";

dffeas \M_st_data[2] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[2]~q ),
	.prn(vcc));
defparam \M_st_data[2] .is_wysiwyg = "true";
defparam \M_st_data[2] .power_up = "low";

dffeas \A_st_data[2] (
	.clk(clk_clk),
	.d(\M_st_data[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[2]~q ),
	.prn(vcc));
defparam \A_st_data[2] .is_wysiwyg = "true";
defparam \A_st_data[2] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[2]~11 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[2]~q ),
	.datad(!\A_st_data[2]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[2]~11 .extended_lut = "off";
defparam \d_writedata_nxt[2]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~67 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[18]~54_combout ),
	.datad(!\E_alu_result[18]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~67 .extended_lut = "off";
defparam \D_src2_reg[18]~67 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[18]~67 .shared_arith = "off";

dffeas \E_src2_reg[18] (
	.clk(clk_clk),
	.d(\D_src2_reg[18]~67_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[18]~q ),
	.prn(vcc));
defparam \E_src2_reg[18] .is_wysiwyg = "true";
defparam \E_src2_reg[18] .power_up = "low";

dffeas \M_st_data[18] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[18]~q ),
	.prn(vcc));
defparam \M_st_data[18] .is_wysiwyg = "true";
defparam \M_st_data[18] .power_up = "low";

dffeas \A_st_data[18] (
	.clk(clk_clk),
	.d(\M_st_data[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[18]~q ),
	.prn(vcc));
defparam \A_st_data[18] .is_wysiwyg = "true";
defparam \A_st_data[18] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[18]~12 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[18]~q ),
	.datad(!\A_st_data[18]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[18]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[18]~12 .extended_lut = "off";
defparam \d_writedata_nxt[18]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[18]~12 .shared_arith = "off";

dffeas \E_src2_reg[10] (
	.clk(clk_clk),
	.d(\D_src2_reg[10]~119_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[10]~q ),
	.prn(vcc));
defparam \E_src2_reg[10] .is_wysiwyg = "true";
defparam \E_src2_reg[10] .power_up = "low";

dffeas \M_st_data[10] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[10]~q ),
	.prn(vcc));
defparam \M_st_data[10] .is_wysiwyg = "true";
defparam \M_st_data[10] .power_up = "low";

dffeas \A_st_data[10] (
	.clk(clk_clk),
	.d(\M_st_data[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[10]~q ),
	.prn(vcc));
defparam \A_st_data[10] .is_wysiwyg = "true";
defparam \A_st_data[10] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[10]~13 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[10]~q ),
	.datad(!\A_st_data[10]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[10]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[10]~13 .extended_lut = "off";
defparam \d_writedata_nxt[10]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[10]~13 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~68 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~68 .extended_lut = "off";
defparam \D_src2_reg[26]~68 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[26]~68 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~69 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~21_combout ),
	.datad(!\Add24~93_sumout ),
	.datae(!\D_src2_reg[26]~68_combout ),
	.dataf(!\D_src2_reg[26]~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~69 .extended_lut = "off";
defparam \D_src2_reg[26]~69 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[26]~69 .shared_arith = "off";

dffeas \E_src2_reg[26] (
	.clk(clk_clk),
	.d(\D_src2_reg[26]~69_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[26]~q ),
	.prn(vcc));
defparam \E_src2_reg[26] .is_wysiwyg = "true";
defparam \E_src2_reg[26] .power_up = "low";

cyclonev_lcell_comb \E_st_data[26]~2 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[2]~q ),
	.datad(!\E_src2_reg[10]~q ),
	.datae(!\E_src2_reg[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~2 .extended_lut = "off";
defparam \E_st_data[26]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[26]~2 .shared_arith = "off";

dffeas \M_st_data[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[26]~q ),
	.prn(vcc));
defparam \M_st_data[26] .is_wysiwyg = "true";
defparam \M_st_data[26] .power_up = "low";

dffeas \A_st_data[26] (
	.clk(clk_clk),
	.d(\M_st_data[26]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[26]~q ),
	.prn(vcc));
defparam \A_st_data[26] .is_wysiwyg = "true";
defparam \A_st_data[26] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[26]~14 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[26]~q ),
	.datad(!\A_st_data[26]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[26]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[26]~14 .extended_lut = "off";
defparam \d_writedata_nxt[26]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[26]~14 .shared_arith = "off";

dffeas \E_src2_reg[5] (
	.clk(clk_clk),
	.d(\D_src2_reg[5]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[5]~q ),
	.prn(vcc));
defparam \E_src2_reg[5] .is_wysiwyg = "true";
defparam \E_src2_reg[5] .power_up = "low";

dffeas \M_st_data[5] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[5]~q ),
	.prn(vcc));
defparam \M_st_data[5] .is_wysiwyg = "true";
defparam \M_st_data[5] .power_up = "low";

dffeas \A_st_data[5] (
	.clk(clk_clk),
	.d(\M_st_data[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[5]~q ),
	.prn(vcc));
defparam \A_st_data[5] .is_wysiwyg = "true";
defparam \A_st_data[5] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[5]~15 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[5]~q ),
	.datad(!\A_st_data[5]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[5]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[5]~15 .extended_lut = "off";
defparam \d_writedata_nxt[5]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[5]~15 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~70 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~70 .extended_lut = "off";
defparam \D_src2_reg[21]~70 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[21]~70 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~71 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~26_combout ),
	.datad(!\Add24~113_sumout ),
	.datae(!\D_src2_reg[21]~70_combout ),
	.dataf(!\D_src2_reg[21]~52_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~71 .extended_lut = "off";
defparam \D_src2_reg[21]~71 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[21]~71 .shared_arith = "off";

dffeas \E_src2_reg[21] (
	.clk(clk_clk),
	.d(\D_src2_reg[21]~71_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[21]~q ),
	.prn(vcc));
defparam \E_src2_reg[21] .is_wysiwyg = "true";
defparam \E_src2_reg[21] .power_up = "low";

dffeas \M_st_data[21] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[21]~q ),
	.prn(vcc));
defparam \M_st_data[21] .is_wysiwyg = "true";
defparam \M_st_data[21] .power_up = "low";

dffeas \A_st_data[21] (
	.clk(clk_clk),
	.d(\M_st_data[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[21]~q ),
	.prn(vcc));
defparam \A_st_data[21] .is_wysiwyg = "true";
defparam \A_st_data[21] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[21]~16 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[21]~q ),
	.datad(!\A_st_data[21]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[21]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[21]~16 .extended_lut = "off";
defparam \d_writedata_nxt[21]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[21]~16 .shared_arith = "off";

dffeas \E_src2_reg[13] (
	.clk(clk_clk),
	.d(\D_src2_reg[13]~99_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[13]~q ),
	.prn(vcc));
defparam \E_src2_reg[13] .is_wysiwyg = "true";
defparam \E_src2_reg[13] .power_up = "low";

dffeas \M_st_data[13] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[13]~q ),
	.prn(vcc));
defparam \M_st_data[13] .is_wysiwyg = "true";
defparam \M_st_data[13] .power_up = "low";

dffeas \A_st_data[13] (
	.clk(clk_clk),
	.d(\M_st_data[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[13]~q ),
	.prn(vcc));
defparam \A_st_data[13] .is_wysiwyg = "true";
defparam \A_st_data[13] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[13]~17 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[13]~q ),
	.datad(!\A_st_data[13]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[13]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[13]~17 .extended_lut = "off";
defparam \d_writedata_nxt[13]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[13]~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~72 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~72 .extended_lut = "off";
defparam \D_src2_reg[29]~72 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[29]~72 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~73 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~17_combout ),
	.datad(!\Add24~81_sumout ),
	.datae(!\D_src2_reg[29]~72_combout ),
	.dataf(!\D_src2_reg[29]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~73 .extended_lut = "off";
defparam \D_src2_reg[29]~73 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[29]~73 .shared_arith = "off";

dffeas \E_src2_reg[29] (
	.clk(clk_clk),
	.d(\D_src2_reg[29]~73_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[29]~q ),
	.prn(vcc));
defparam \E_src2_reg[29] .is_wysiwyg = "true";
defparam \E_src2_reg[29] .power_up = "low";

cyclonev_lcell_comb \E_st_data[29]~3 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[5]~q ),
	.datad(!\E_src2_reg[13]~q ),
	.datae(!\E_src2_reg[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~3 .extended_lut = "off";
defparam \E_st_data[29]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[29]~3 .shared_arith = "off";

dffeas \M_st_data[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[29]~q ),
	.prn(vcc));
defparam \M_st_data[29] .is_wysiwyg = "true";
defparam \M_st_data[29] .power_up = "low";

dffeas \A_st_data[29] (
	.clk(clk_clk),
	.d(\M_st_data[29]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[29]~q ),
	.prn(vcc));
defparam \A_st_data[29] .is_wysiwyg = "true";
defparam \A_st_data[29] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[29]~18 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[29]~q ),
	.datad(!\A_st_data[29]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[29]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[29]~18 .extended_lut = "off";
defparam \d_writedata_nxt[29]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[29]~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~74 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~74 .extended_lut = "off";
defparam \D_src2_reg[23]~74 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[23]~74 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~75 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~30_combout ),
	.datad(!\Add24~129_sumout ),
	.datae(!\D_src2_reg[23]~74_combout ),
	.dataf(!\D_src2_reg[23]~59_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~75 .extended_lut = "off";
defparam \D_src2_reg[23]~75 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[23]~75 .shared_arith = "off";

dffeas \E_src2_reg[23] (
	.clk(clk_clk),
	.d(\D_src2_reg[23]~75_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[23]~q ),
	.prn(vcc));
defparam \E_src2_reg[23] .is_wysiwyg = "true";
defparam \E_src2_reg[23] .power_up = "low";

dffeas \M_st_data[23] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[23]~q ),
	.prn(vcc));
defparam \M_st_data[23] .is_wysiwyg = "true";
defparam \M_st_data[23] .power_up = "low";

dffeas \A_st_data[23] (
	.clk(clk_clk),
	.d(\M_st_data[23]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[23]~q ),
	.prn(vcc));
defparam \A_st_data[23] .is_wysiwyg = "true";
defparam \A_st_data[23] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[23]~19 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[23]~q ),
	.datad(!\A_st_data[23]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[23]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[23]~19 .extended_lut = "off";
defparam \d_writedata_nxt[23]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[23]~19 .shared_arith = "off";

dffeas \E_src2_reg[15] (
	.clk(clk_clk),
	.d(\D_src2_reg[15]~107_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[15]~q ),
	.prn(vcc));
defparam \E_src2_reg[15] .is_wysiwyg = "true";
defparam \E_src2_reg[15] .power_up = "low";

dffeas \M_st_data[15] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[15]~q ),
	.prn(vcc));
defparam \M_st_data[15] .is_wysiwyg = "true";
defparam \M_st_data[15] .power_up = "low";

dffeas \A_st_data[15] (
	.clk(clk_clk),
	.d(\M_st_data[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[15]~q ),
	.prn(vcc));
defparam \A_st_data[15] .is_wysiwyg = "true";
defparam \A_st_data[15] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[15]~20 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[15]~q ),
	.datad(!\A_st_data[15]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[15]~20 .extended_lut = "off";
defparam \d_writedata_nxt[15]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[15]~20 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~76 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~76 .extended_lut = "off";
defparam \D_src2_reg[31]~76 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_src2_reg[31]~76 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~77 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add24~37_sumout ),
	.datac(!\D_src2_reg[0]~31_combout ),
	.datad(!\E_alu_result~31_combout ),
	.datae(!\D_src2_reg[31]~76_combout ),
	.dataf(!\D_src2_reg[31]~61_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~77 .extended_lut = "off";
defparam \D_src2_reg[31]~77 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[31]~77 .shared_arith = "off";

dffeas \E_src2_reg[31] (
	.clk(clk_clk),
	.d(\D_src2_reg[31]~77_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[31]~q ),
	.prn(vcc));
defparam \E_src2_reg[31] .is_wysiwyg = "true";
defparam \E_src2_reg[31] .power_up = "low";

cyclonev_lcell_comb \E_st_data[31]~4 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[7]~q ),
	.datad(!\E_src2_reg[15]~q ),
	.datae(!\E_src2_reg[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~4 .extended_lut = "off";
defparam \E_st_data[31]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[31]~4 .shared_arith = "off";

dffeas \M_st_data[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[31]~q ),
	.prn(vcc));
defparam \M_st_data[31] .is_wysiwyg = "true";
defparam \M_st_data[31] .power_up = "low";

dffeas \A_st_data[31] (
	.clk(clk_clk),
	.d(\M_st_data[31]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[31]~q ),
	.prn(vcc));
defparam \A_st_data[31] .is_wysiwyg = "true";
defparam \A_st_data[31] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[31]~21 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[31]~q ),
	.datad(!\A_st_data[31]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[31]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[31]~21 .extended_lut = "off";
defparam \d_writedata_nxt[31]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[31]~21 .shared_arith = "off";

dffeas \E_src2_reg[11] (
	.clk(clk_clk),
	.d(\D_src2_reg[11]~123_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[11]~q ),
	.prn(vcc));
defparam \E_src2_reg[11] .is_wysiwyg = "true";
defparam \E_src2_reg[11] .power_up = "low";

dffeas \M_st_data[11] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[11]~q ),
	.prn(vcc));
defparam \M_st_data[11] .is_wysiwyg = "true";
defparam \M_st_data[11] .power_up = "low";

dffeas \A_st_data[11] (
	.clk(clk_clk),
	.d(\M_st_data[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[11]~q ),
	.prn(vcc));
defparam \A_st_data[11] .is_wysiwyg = "true";
defparam \A_st_data[11] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[11]~22 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[11]~q ),
	.datad(!\A_st_data[11]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[11]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[11]~22 .extended_lut = "off";
defparam \d_writedata_nxt[11]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[11]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~78 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~78 .extended_lut = "off";
defparam \D_src2_reg[27]~78 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[27]~78 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~79 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~19_combout ),
	.datad(!\Add24~89_sumout ),
	.datae(!\D_src2_reg[27]~78_combout ),
	.dataf(!\D_src2_reg[27]~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~79 .extended_lut = "off";
defparam \D_src2_reg[27]~79 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[27]~79 .shared_arith = "off";

dffeas \E_src2_reg[27] (
	.clk(clk_clk),
	.d(\D_src2_reg[27]~79_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[27]~q ),
	.prn(vcc));
defparam \E_src2_reg[27] .is_wysiwyg = "true";
defparam \E_src2_reg[27] .power_up = "low";

cyclonev_lcell_comb \E_st_data[27]~5 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[3]~q ),
	.datad(!\E_src2_reg[11]~q ),
	.datae(!\E_src2_reg[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~5 .extended_lut = "off";
defparam \E_st_data[27]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[27]~5 .shared_arith = "off";

dffeas \M_st_data[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[27]~q ),
	.prn(vcc));
defparam \M_st_data[27] .is_wysiwyg = "true";
defparam \M_st_data[27] .power_up = "low";

dffeas \A_st_data[27] (
	.clk(clk_clk),
	.d(\M_st_data[27]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[27]~q ),
	.prn(vcc));
defparam \A_st_data[27] .is_wysiwyg = "true";
defparam \A_st_data[27] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[27]~23 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[27]~q ),
	.datad(!\A_st_data[27]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[27]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[27]~23 .extended_lut = "off";
defparam \d_writedata_nxt[27]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[27]~23 .shared_arith = "off";

dffeas \E_src2_reg[9] (
	.clk(clk_clk),
	.d(\D_src2_reg[9]~115_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[9]~q ),
	.prn(vcc));
defparam \E_src2_reg[9] .is_wysiwyg = "true";
defparam \E_src2_reg[9] .power_up = "low";

dffeas \M_st_data[9] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[9]~q ),
	.prn(vcc));
defparam \M_st_data[9] .is_wysiwyg = "true";
defparam \M_st_data[9] .power_up = "low";

dffeas \A_st_data[9] (
	.clk(clk_clk),
	.d(\M_st_data[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[9]~q ),
	.prn(vcc));
defparam \A_st_data[9] .is_wysiwyg = "true";
defparam \A_st_data[9] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[9]~24 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[9]~q ),
	.datad(!\A_st_data[9]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[9]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[9]~24 .extended_lut = "off";
defparam \d_writedata_nxt[9]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[9]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~80 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~80 .extended_lut = "off";
defparam \D_src2_reg[25]~80 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[25]~80 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~81 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~22_combout ),
	.datad(!\Add24~97_sumout ),
	.datae(!\D_src2_reg[25]~80_combout ),
	.dataf(!\D_src2_reg[25]~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~81 .extended_lut = "off";
defparam \D_src2_reg[25]~81 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[25]~81 .shared_arith = "off";

dffeas \E_src2_reg[25] (
	.clk(clk_clk),
	.d(\D_src2_reg[25]~81_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[25]~q ),
	.prn(vcc));
defparam \E_src2_reg[25] .is_wysiwyg = "true";
defparam \E_src2_reg[25] .power_up = "low";

cyclonev_lcell_comb \E_st_data[25]~6 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[1]~q ),
	.datad(!\E_src2_reg[9]~q ),
	.datae(!\E_src2_reg[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~6 .extended_lut = "off";
defparam \E_st_data[25]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[25]~6 .shared_arith = "off";

dffeas \M_st_data[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[25]~q ),
	.prn(vcc));
defparam \M_st_data[25] .is_wysiwyg = "true";
defparam \M_st_data[25] .power_up = "low";

dffeas \A_st_data[25] (
	.clk(clk_clk),
	.d(\M_st_data[25]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[25]~q ),
	.prn(vcc));
defparam \A_st_data[25] .is_wysiwyg = "true";
defparam \A_st_data[25] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[25]~25 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[25]~q ),
	.datad(!\A_st_data[25]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[25]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[25]~25 .extended_lut = "off";
defparam \d_writedata_nxt[25]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[25]~25 .shared_arith = "off";

dffeas \E_src2_reg[6] (
	.clk(clk_clk),
	.d(\D_src2_reg[6]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[6]~q ),
	.prn(vcc));
defparam \E_src2_reg[6] .is_wysiwyg = "true";
defparam \E_src2_reg[6] .power_up = "low";

dffeas \M_st_data[6] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[6]~q ),
	.prn(vcc));
defparam \M_st_data[6] .is_wysiwyg = "true";
defparam \M_st_data[6] .power_up = "low";

dffeas \A_st_data[6] (
	.clk(clk_clk),
	.d(\M_st_data[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[6]~q ),
	.prn(vcc));
defparam \A_st_data[6] .is_wysiwyg = "true";
defparam \A_st_data[6] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[6]~26 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[6]~q ),
	.datad(!\A_st_data[6]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[6]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[6]~26 .extended_lut = "off";
defparam \d_writedata_nxt[6]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[6]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~82 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~82 .extended_lut = "off";
defparam \D_src2_reg[22]~82 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[22]~82 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~83 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\E_alu_result~25_combout ),
	.datad(!\Add24~109_sumout ),
	.datae(!\D_src2_reg[22]~82_combout ),
	.dataf(!\D_src2_reg[22]~50_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~83 .extended_lut = "off";
defparam \D_src2_reg[22]~83 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[22]~83 .shared_arith = "off";

dffeas \E_src2_reg[22] (
	.clk(clk_clk),
	.d(\D_src2_reg[22]~83_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[22]~q ),
	.prn(vcc));
defparam \E_src2_reg[22] .is_wysiwyg = "true";
defparam \E_src2_reg[22] .power_up = "low";

dffeas \M_st_data[22] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[22]~q ),
	.prn(vcc));
defparam \M_st_data[22] .is_wysiwyg = "true";
defparam \M_st_data[22] .power_up = "low";

dffeas \A_st_data[22] (
	.clk(clk_clk),
	.d(\M_st_data[22]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[22]~q ),
	.prn(vcc));
defparam \A_st_data[22] .is_wysiwyg = "true";
defparam \A_st_data[22] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[22]~27 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[22]~q ),
	.datad(!\A_st_data[22]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[22]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[22]~27 .extended_lut = "off";
defparam \d_writedata_nxt[22]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[22]~27 .shared_arith = "off";

dffeas \E_src2_reg[14] (
	.clk(clk_clk),
	.d(\D_src2_reg[14]~103_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[14]~q ),
	.prn(vcc));
defparam \E_src2_reg[14] .is_wysiwyg = "true";
defparam \E_src2_reg[14] .power_up = "low";

dffeas \M_st_data[14] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[14]~q ),
	.prn(vcc));
defparam \M_st_data[14] .is_wysiwyg = "true";
defparam \M_st_data[14] .power_up = "low";

dffeas \A_st_data[14] (
	.clk(clk_clk),
	.d(\M_st_data[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[14]~q ),
	.prn(vcc));
defparam \A_st_data[14] .is_wysiwyg = "true";
defparam \A_st_data[14] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[14]~28 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[14]~q ),
	.datad(!\A_st_data[14]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[14]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[14]~28 .extended_lut = "off";
defparam \d_writedata_nxt[14]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[14]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~84 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[29]~0_combout ),
	.datad(!\Equal299~0_combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~84 .extended_lut = "off";
defparam \D_src2_reg[30]~84 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_src2_reg[30]~84 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~85 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~31_combout ),
	.datac(!\Add24~77_sumout ),
	.datad(!\E_alu_result~20_combout ),
	.datae(!\D_src2_reg[30]~84_combout ),
	.dataf(!\D_src2_reg[30]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~85 .extended_lut = "off";
defparam \D_src2_reg[30]~85 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \D_src2_reg[30]~85 .shared_arith = "off";

dffeas \E_src2_reg[30] (
	.clk(clk_clk),
	.d(\D_src2_reg[30]~85_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[30]~q ),
	.prn(vcc));
defparam \E_src2_reg[30] .is_wysiwyg = "true";
defparam \E_src2_reg[30] .power_up = "low";

cyclonev_lcell_comb \E_st_data[30]~7 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[6]~q ),
	.datad(!\E_src2_reg[14]~q ),
	.datae(!\E_src2_reg[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~7 .extended_lut = "off";
defparam \E_st_data[30]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[30]~7 .shared_arith = "off";

dffeas \M_st_data[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[30]~q ),
	.prn(vcc));
defparam \M_st_data[30] .is_wysiwyg = "true";
defparam \M_st_data[30] .power_up = "low";

dffeas \A_st_data[30] (
	.clk(clk_clk),
	.d(\M_st_data[30]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[30]~q ),
	.prn(vcc));
defparam \A_st_data[30] .is_wysiwyg = "true";
defparam \A_st_data[30] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[30]~29 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[30]~q ),
	.datad(!\A_st_data[30]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[30]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[30]~29 .extended_lut = "off";
defparam \d_writedata_nxt[30]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[30]~29 .shared_arith = "off";

dffeas \E_src2_reg[19] (
	.clk(clk_clk),
	.d(\D_src2_reg[19]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[19]~q ),
	.prn(vcc));
defparam \E_src2_reg[19] .is_wysiwyg = "true";
defparam \E_src2_reg[19] .power_up = "low";

dffeas \M_st_data[19] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[19]~q ),
	.prn(vcc));
defparam \M_st_data[19] .is_wysiwyg = "true";
defparam \M_st_data[19] .power_up = "low";

dffeas \A_st_data[19] (
	.clk(clk_clk),
	.d(\M_st_data[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[19]~q ),
	.prn(vcc));
defparam \A_st_data[19] .is_wysiwyg = "true";
defparam \A_st_data[19] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[19]~30 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[19]~q ),
	.datad(!\A_st_data[19]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[19]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[19]~30 .extended_lut = "off";
defparam \d_writedata_nxt[19]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[19]~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[17]~86 (
	.dataa(!\D_src2_reg[29]~1_combout ),
	.datab(!\D_src2_reg[29]~2_combout ),
	.datac(!\D_src2_reg[17]~47_combout ),
	.datad(!\E_alu_result[17]~combout ),
	.datae(!\Qsys_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~86 .extended_lut = "off";
defparam \D_src2_reg[17]~86 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[17]~86 .shared_arith = "off";

dffeas \E_src2_reg[17] (
	.clk(clk_clk),
	.d(\D_src2_reg[17]~86_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[17]~q ),
	.prn(vcc));
defparam \E_src2_reg[17] .is_wysiwyg = "true";
defparam \E_src2_reg[17] .power_up = "low";

dffeas \M_st_data[17] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[17]~q ),
	.prn(vcc));
defparam \M_st_data[17] .is_wysiwyg = "true";
defparam \M_st_data[17] .power_up = "low";

dffeas \A_st_data[17] (
	.clk(clk_clk),
	.d(\M_st_data[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[17]~q ),
	.prn(vcc));
defparam \A_st_data[17] .is_wysiwyg = "true";
defparam \A_st_data[17] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[17]~31 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[17]~q ),
	.datad(!\A_st_data[17]~q ),
	.datae(!\Qsys_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[17]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[17]~31 .extended_lut = "off";
defparam \d_writedata_nxt[17]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[17]~31 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_bht_module (
	q_b_1,
	q_b_0,
	F_stall,
	M_bht_wr_en_unfiltered,
	M_bht_wr_data_unfiltered_1,
	M_bht_ptr_unfiltered_0,
	M_bht_ptr_unfiltered_1,
	M_bht_ptr_unfiltered_2,
	M_bht_ptr_unfiltered_3,
	M_bht_ptr_unfiltered_4,
	M_bht_ptr_unfiltered_5,
	M_bht_ptr_unfiltered_6,
	M_bht_ptr_unfiltered_7,
	F_bht_ptr_nxt_0,
	F_bht_ptr_nxt_1,
	F_bht_ptr_nxt_2,
	F_bht_ptr_nxt_3,
	F_bht_ptr_nxt_4,
	F_bht_ptr_nxt_5,
	F_bht_ptr_nxt_6,
	F_bht_ptr_nxt_7,
	M_br_mispredict,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
input 	F_stall;
input 	M_bht_wr_en_unfiltered;
input 	M_bht_wr_data_unfiltered_1;
input 	M_bht_ptr_unfiltered_0;
input 	M_bht_ptr_unfiltered_1;
input 	M_bht_ptr_unfiltered_2;
input 	M_bht_ptr_unfiltered_3;
input 	M_bht_ptr_unfiltered_4;
input 	M_bht_ptr_unfiltered_5;
input 	M_bht_ptr_unfiltered_6;
input 	M_bht_ptr_unfiltered_7;
input 	F_bht_ptr_nxt_0;
input 	F_bht_ptr_nxt_1;
input 	F_bht_ptr_nxt_2;
input 	F_bht_ptr_nxt_3;
input 	F_bht_ptr_nxt_4;
input 	F_bht_ptr_nxt_5;
input 	F_bht_ptr_nxt_6;
input 	F_bht_ptr_nxt_7;
input 	M_br_mispredict;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_1 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_1,q_b_0}),
	.rden_b(F_stall),
	.wren_a(M_bht_wr_en_unfiltered),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,M_bht_wr_data_unfiltered_1,M_br_mispredict}),
	.address_a({gnd,gnd,gnd,gnd,gnd,M_bht_ptr_unfiltered_7,M_bht_ptr_unfiltered_6,M_bht_ptr_unfiltered_5,M_bht_ptr_unfiltered_4,M_bht_ptr_unfiltered_3,M_bht_ptr_unfiltered_2,M_bht_ptr_unfiltered_1,M_bht_ptr_unfiltered_0}),
	.address_b({gnd,gnd,F_bht_ptr_nxt_7,F_bht_ptr_nxt_6,F_bht_ptr_nxt_5,F_bht_ptr_nxt_4,F_bht_ptr_nxt_3,F_bht_ptr_nxt_2,F_bht_ptr_nxt_1,F_bht_ptr_nxt_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_f4o1 auto_generated(
	.q_b({q_b[1],q_b[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_f4o1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[1:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[1:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_bht_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_bht_module:Qsys_system_nios2_qsys_0_bht|altsyncram:the_altsyncram|altsyncram_f4o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 2;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 2;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "47FA19FCB2124EB3FB783923FDBBAA3EC40C758C6F9E56B3BBC04C1B566B8EEE";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_bht_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_bht_module:Qsys_system_nios2_qsys_0_bht|altsyncram:the_altsyncram|altsyncram_f4o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 2;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "E85DFB4B53DA445E12F71630B1B6463EF6602B57E2A6B55EA0889FF222FAD437";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_dc_data_module (
	q_b_0,
	q_b_4,
	q_b_20,
	q_b_12,
	q_b_28,
	q_b_16,
	q_b_8,
	q_b_24,
	q_b_2,
	q_b_18,
	q_b_10,
	q_b_26,
	q_b_5,
	q_b_21,
	q_b_13,
	q_b_29,
	q_b_7,
	q_b_23,
	q_b_15,
	q_b_31,
	q_b_11,
	q_b_27,
	q_b_9,
	q_b_25,
	q_b_6,
	q_b_22,
	q_b_14,
	q_b_30,
	q_b_3,
	q_b_19,
	q_b_1,
	q_b_17,
	dc_data_wr_port_en,
	dc_data_wr_port_data_0,
	dc_data_wr_port_addr_0,
	dc_data_wr_port_addr_1,
	dc_data_wr_port_addr_2,
	dc_data_wr_port_addr_3,
	dc_data_wr_port_addr_4,
	dc_data_wr_port_addr_5,
	dc_data_wr_port_addr_6,
	dc_data_wr_port_addr_7,
	dc_data_wr_port_addr_8,
	dc_data_rd_port_addr_0,
	dc_data_rd_port_addr_1,
	dc_data_rd_port_addr_2,
	dc_data_rd_port_addr_3,
	dc_data_rd_port_addr_4,
	dc_data_rd_port_addr_5,
	dc_data_rd_port_addr_6,
	dc_data_rd_port_addr_7,
	dc_data_rd_port_addr_8,
	dc_data_wr_port_data_4,
	dc_data_wr_port_data_20,
	dc_data_wr_port_data_12,
	dc_data_wr_port_data_28,
	dc_data_wr_port_data_16,
	dc_data_wr_port_data_8,
	dc_data_wr_port_data_24,
	dc_data_wr_port_data_2,
	dc_data_wr_port_data_18,
	dc_data_wr_port_data_10,
	dc_data_wr_port_data_26,
	dc_data_wr_port_data_5,
	dc_data_wr_port_data_21,
	dc_data_wr_port_data_13,
	dc_data_wr_port_data_29,
	dc_data_wr_port_data_7,
	dc_data_wr_port_data_23,
	dc_data_wr_port_data_15,
	dc_data_wr_port_data_31,
	dc_data_wr_port_data_11,
	dc_data_wr_port_data_27,
	dc_data_wr_port_data_9,
	dc_data_wr_port_data_25,
	dc_data_wr_port_data_6,
	dc_data_wr_port_data_22,
	dc_data_wr_port_data_14,
	dc_data_wr_port_data_30,
	dc_data_wr_port_data_3,
	dc_data_wr_port_data_19,
	dc_data_wr_port_data_1,
	dc_data_wr_port_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_4;
output 	q_b_20;
output 	q_b_12;
output 	q_b_28;
output 	q_b_16;
output 	q_b_8;
output 	q_b_24;
output 	q_b_2;
output 	q_b_18;
output 	q_b_10;
output 	q_b_26;
output 	q_b_5;
output 	q_b_21;
output 	q_b_13;
output 	q_b_29;
output 	q_b_7;
output 	q_b_23;
output 	q_b_15;
output 	q_b_31;
output 	q_b_11;
output 	q_b_27;
output 	q_b_9;
output 	q_b_25;
output 	q_b_6;
output 	q_b_22;
output 	q_b_14;
output 	q_b_30;
output 	q_b_3;
output 	q_b_19;
output 	q_b_1;
output 	q_b_17;
input 	dc_data_wr_port_en;
input 	dc_data_wr_port_data_0;
input 	dc_data_wr_port_addr_0;
input 	dc_data_wr_port_addr_1;
input 	dc_data_wr_port_addr_2;
input 	dc_data_wr_port_addr_3;
input 	dc_data_wr_port_addr_4;
input 	dc_data_wr_port_addr_5;
input 	dc_data_wr_port_addr_6;
input 	dc_data_wr_port_addr_7;
input 	dc_data_wr_port_addr_8;
input 	dc_data_rd_port_addr_0;
input 	dc_data_rd_port_addr_1;
input 	dc_data_rd_port_addr_2;
input 	dc_data_rd_port_addr_3;
input 	dc_data_rd_port_addr_4;
input 	dc_data_rd_port_addr_5;
input 	dc_data_rd_port_addr_6;
input 	dc_data_rd_port_addr_7;
input 	dc_data_rd_port_addr_8;
input 	dc_data_wr_port_data_4;
input 	dc_data_wr_port_data_20;
input 	dc_data_wr_port_data_12;
input 	dc_data_wr_port_data_28;
input 	dc_data_wr_port_data_16;
input 	dc_data_wr_port_data_8;
input 	dc_data_wr_port_data_24;
input 	dc_data_wr_port_data_2;
input 	dc_data_wr_port_data_18;
input 	dc_data_wr_port_data_10;
input 	dc_data_wr_port_data_26;
input 	dc_data_wr_port_data_5;
input 	dc_data_wr_port_data_21;
input 	dc_data_wr_port_data_13;
input 	dc_data_wr_port_data_29;
input 	dc_data_wr_port_data_7;
input 	dc_data_wr_port_data_23;
input 	dc_data_wr_port_data_15;
input 	dc_data_wr_port_data_31;
input 	dc_data_wr_port_data_11;
input 	dc_data_wr_port_data_27;
input 	dc_data_wr_port_data_9;
input 	dc_data_wr_port_data_25;
input 	dc_data_wr_port_data_6;
input 	dc_data_wr_port_data_22;
input 	dc_data_wr_port_data_14;
input 	dc_data_wr_port_data_30;
input 	dc_data_wr_port_data_3;
input 	dc_data_wr_port_data_19;
input 	dc_data_wr_port_data_1;
input 	dc_data_wr_port_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(dc_data_wr_port_en),
	.data_a({dc_data_wr_port_data_31,dc_data_wr_port_data_30,dc_data_wr_port_data_29,dc_data_wr_port_data_28,dc_data_wr_port_data_27,dc_data_wr_port_data_26,dc_data_wr_port_data_25,dc_data_wr_port_data_24,dc_data_wr_port_data_23,dc_data_wr_port_data_22,dc_data_wr_port_data_21,
dc_data_wr_port_data_20,dc_data_wr_port_data_19,dc_data_wr_port_data_18,dc_data_wr_port_data_17,dc_data_wr_port_data_16,dc_data_wr_port_data_15,dc_data_wr_port_data_14,dc_data_wr_port_data_13,dc_data_wr_port_data_12,dc_data_wr_port_data_11,dc_data_wr_port_data_10,
dc_data_wr_port_data_9,dc_data_wr_port_data_8,dc_data_wr_port_data_7,dc_data_wr_port_data_6,dc_data_wr_port_data_5,dc_data_wr_port_data_4,dc_data_wr_port_data_3,dc_data_wr_port_data_2,dc_data_wr_port_data_1,dc_data_wr_port_data_0}),
	.address_a({gnd,gnd,gnd,gnd,dc_data_wr_port_addr_8,dc_data_wr_port_addr_7,dc_data_wr_port_addr_6,dc_data_wr_port_addr_5,dc_data_wr_port_addr_4,dc_data_wr_port_addr_3,dc_data_wr_port_addr_2,dc_data_wr_port_addr_1,dc_data_wr_port_addr_0}),
	.address_b({gnd,dc_data_rd_port_addr_8,dc_data_rd_port_addr_7,dc_data_rd_port_addr_6,dc_data_rd_port_addr_5,dc_data_rd_port_addr_4,dc_data_rd_port_addr_3,dc_data_rd_port_addr_2,dc_data_rd_port_addr_1,dc_data_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_40j1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_40j1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 9;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 511;
defparam ram_block1a4.port_a_logical_ram_depth = 512;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 9;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 511;
defparam ram_block1a4.port_b_logical_ram_depth = 512;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 9;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 511;
defparam ram_block1a20.port_a_logical_ram_depth = 512;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 9;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 511;
defparam ram_block1a20.port_b_logical_ram_depth = 512;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 9;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 511;
defparam ram_block1a12.port_a_logical_ram_depth = 512;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 9;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 511;
defparam ram_block1a12.port_b_logical_ram_depth = 512;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 9;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 511;
defparam ram_block1a28.port_a_logical_ram_depth = 512;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 9;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 511;
defparam ram_block1a28.port_b_logical_ram_depth = 512;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 9;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 511;
defparam ram_block1a16.port_a_logical_ram_depth = 512;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 9;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 511;
defparam ram_block1a16.port_b_logical_ram_depth = 512;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 9;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 511;
defparam ram_block1a8.port_a_logical_ram_depth = 512;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 9;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 511;
defparam ram_block1a8.port_b_logical_ram_depth = 512;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 9;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 511;
defparam ram_block1a24.port_a_logical_ram_depth = 512;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 9;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 511;
defparam ram_block1a24.port_b_logical_ram_depth = 512;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 9;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 511;
defparam ram_block1a2.port_a_logical_ram_depth = 512;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 9;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 511;
defparam ram_block1a2.port_b_logical_ram_depth = 512;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 9;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 511;
defparam ram_block1a18.port_a_logical_ram_depth = 512;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 9;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 511;
defparam ram_block1a18.port_b_logical_ram_depth = 512;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 9;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 511;
defparam ram_block1a10.port_a_logical_ram_depth = 512;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 9;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 511;
defparam ram_block1a10.port_b_logical_ram_depth = 512;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 9;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 511;
defparam ram_block1a26.port_a_logical_ram_depth = 512;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 9;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 511;
defparam ram_block1a26.port_b_logical_ram_depth = 512;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 9;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 511;
defparam ram_block1a5.port_a_logical_ram_depth = 512;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 9;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 511;
defparam ram_block1a5.port_b_logical_ram_depth = 512;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 9;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 511;
defparam ram_block1a21.port_a_logical_ram_depth = 512;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 9;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 511;
defparam ram_block1a21.port_b_logical_ram_depth = 512;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 9;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 511;
defparam ram_block1a13.port_a_logical_ram_depth = 512;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 9;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 511;
defparam ram_block1a13.port_b_logical_ram_depth = 512;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 9;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 511;
defparam ram_block1a29.port_a_logical_ram_depth = 512;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 9;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 511;
defparam ram_block1a29.port_b_logical_ram_depth = 512;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 9;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 511;
defparam ram_block1a7.port_a_logical_ram_depth = 512;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 9;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 511;
defparam ram_block1a7.port_b_logical_ram_depth = 512;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 9;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 511;
defparam ram_block1a23.port_a_logical_ram_depth = 512;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 9;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 511;
defparam ram_block1a23.port_b_logical_ram_depth = 512;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 9;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 511;
defparam ram_block1a15.port_a_logical_ram_depth = 512;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 9;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 511;
defparam ram_block1a15.port_b_logical_ram_depth = 512;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 9;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 511;
defparam ram_block1a31.port_a_logical_ram_depth = 512;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 9;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 511;
defparam ram_block1a31.port_b_logical_ram_depth = 512;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 9;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 511;
defparam ram_block1a11.port_a_logical_ram_depth = 512;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 9;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 511;
defparam ram_block1a11.port_b_logical_ram_depth = 512;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 9;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 511;
defparam ram_block1a27.port_a_logical_ram_depth = 512;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 9;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 511;
defparam ram_block1a27.port_b_logical_ram_depth = 512;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 9;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 511;
defparam ram_block1a9.port_a_logical_ram_depth = 512;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 9;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 511;
defparam ram_block1a9.port_b_logical_ram_depth = 512;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 9;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 511;
defparam ram_block1a25.port_a_logical_ram_depth = 512;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 9;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 511;
defparam ram_block1a25.port_b_logical_ram_depth = 512;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 9;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 511;
defparam ram_block1a6.port_a_logical_ram_depth = 512;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 9;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 511;
defparam ram_block1a6.port_b_logical_ram_depth = 512;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 9;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 511;
defparam ram_block1a22.port_a_logical_ram_depth = 512;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 9;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 511;
defparam ram_block1a22.port_b_logical_ram_depth = 512;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 9;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 511;
defparam ram_block1a14.port_a_logical_ram_depth = 512;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 9;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 511;
defparam ram_block1a14.port_b_logical_ram_depth = 512;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 9;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 511;
defparam ram_block1a30.port_a_logical_ram_depth = 512;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 9;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 511;
defparam ram_block1a30.port_b_logical_ram_depth = 512;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 9;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 511;
defparam ram_block1a3.port_a_logical_ram_depth = 512;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 9;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 511;
defparam ram_block1a3.port_b_logical_ram_depth = 512;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 9;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 511;
defparam ram_block1a19.port_a_logical_ram_depth = 512;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 9;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 511;
defparam ram_block1a19.port_b_logical_ram_depth = 512;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_data_module:Qsys_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 9;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 511;
defparam ram_block1a17.port_a_logical_ram_depth = 512;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 9;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 511;
defparam ram_block1a17.port_b_logical_ram_depth = 512;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_dc_tag_module (
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_7,
	dc_tag_wr_port_en,
	dc_tag_wr_port_data_4,
	dc_tag_wr_port_addr_0,
	dc_tag_wr_port_addr_1,
	dc_tag_wr_port_addr_2,
	dc_tag_wr_port_addr_3,
	dc_tag_wr_port_addr_4,
	dc_tag_wr_port_addr_5,
	dc_tag_rd_port_addr_0,
	dc_tag_rd_port_addr_1,
	dc_tag_rd_port_addr_2,
	dc_tag_rd_port_addr_3,
	dc_tag_rd_port_addr_4,
	dc_tag_rd_port_addr_5,
	dc_tag_wr_port_data_5,
	dc_tag_wr_port_data_6,
	dc_tag_wr_port_data_0,
	dc_tag_wr_port_data_1,
	dc_tag_wr_port_data_2,
	dc_tag_wr_port_data_3,
	dc_tag_wr_port_data_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_7;
input 	dc_tag_wr_port_en;
input 	dc_tag_wr_port_data_4;
input 	dc_tag_wr_port_addr_0;
input 	dc_tag_wr_port_addr_1;
input 	dc_tag_wr_port_addr_2;
input 	dc_tag_wr_port_addr_3;
input 	dc_tag_wr_port_addr_4;
input 	dc_tag_wr_port_addr_5;
input 	dc_tag_rd_port_addr_0;
input 	dc_tag_rd_port_addr_1;
input 	dc_tag_rd_port_addr_2;
input 	dc_tag_rd_port_addr_3;
input 	dc_tag_rd_port_addr_4;
input 	dc_tag_rd_port_addr_5;
input 	dc_tag_wr_port_data_5;
input 	dc_tag_wr_port_data_6;
input 	dc_tag_wr_port_data_0;
input 	dc_tag_wr_port_data_1;
input 	dc_tag_wr_port_data_2;
input 	dc_tag_wr_port_data_3;
input 	dc_tag_wr_port_data_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_3 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(dc_tag_wr_port_en),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dc_tag_wr_port_data_7,dc_tag_wr_port_data_6,dc_tag_wr_port_data_5,dc_tag_wr_port_data_4,dc_tag_wr_port_data_3,dc_tag_wr_port_data_2,dc_tag_wr_port_data_1,dc_tag_wr_port_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,dc_tag_wr_port_addr_5,dc_tag_wr_port_addr_4,dc_tag_wr_port_addr_3,dc_tag_wr_port_addr_2,dc_tag_wr_port_addr_1,dc_tag_wr_port_addr_0}),
	.address_b({gnd,gnd,gnd,gnd,dc_tag_rd_port_addr_5,dc_tag_rd_port_addr_4,dc_tag_rd_port_addr_3,dc_tag_rd_port_addr_2,dc_tag_rd_port_addr_1,dc_tag_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_bmn1 auto_generated(
	.q_b({q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_bmn1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "213D88B7D0F0E5B1";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "A3CC6CAD97DF7A85";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "A4D8522DE84C47AD";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "2BD4632004610FB3";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FB6F31394B5E9B8D";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "F8A16A39AD4A669B";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "B080F4B85A47B308";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_tag_module:Qsys_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_bmn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "8691A9DB70998817";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_dc_victim_module (
	q_b_0,
	A_dc_xfer_wr_data_0,
	q_b_7,
	q_b_3,
	A_dc_xfer_wr_data_7,
	q_b_1,
	A_dc_xfer_wr_data_3,
	q_b_4,
	q_b_20,
	q_b_12,
	q_b_28,
	q_b_16,
	q_b_8,
	q_b_24,
	q_b_2,
	q_b_18,
	q_b_10,
	q_b_26,
	q_b_5,
	q_b_21,
	q_b_13,
	q_b_29,
	q_b_23,
	q_b_15,
	q_b_31,
	q_b_11,
	q_b_27,
	q_b_9,
	q_b_25,
	q_b_6,
	q_b_22,
	q_b_14,
	q_b_30,
	q_b_19,
	A_dc_xfer_wr_data_1,
	q_b_17,
	A_dc_xfer_wr_data_4,
	A_dc_xfer_wr_data_20,
	A_dc_xfer_wr_data_12,
	A_dc_xfer_wr_data_28,
	A_dc_xfer_wr_data_16,
	A_dc_xfer_wr_data_8,
	A_dc_xfer_wr_data_24,
	A_dc_xfer_wr_data_2,
	A_dc_xfer_wr_data_18,
	A_dc_xfer_wr_data_10,
	A_dc_xfer_wr_data_26,
	A_dc_xfer_wr_data_5,
	A_dc_xfer_wr_data_21,
	A_dc_xfer_wr_data_13,
	A_dc_xfer_wr_data_29,
	A_dc_xfer_wr_data_23,
	A_dc_xfer_wr_data_15,
	A_dc_xfer_wr_data_31,
	A_dc_xfer_wr_data_11,
	A_dc_xfer_wr_data_27,
	A_dc_xfer_wr_data_9,
	A_dc_xfer_wr_data_25,
	A_dc_xfer_wr_data_6,
	A_dc_xfer_wr_data_22,
	A_dc_xfer_wr_data_14,
	A_dc_xfer_wr_data_30,
	A_dc_xfer_wr_data_19,
	A_dc_xfer_wr_data_17,
	A_dc_xfer_wr_active,
	A_dc_wb_rd_en,
	A_dc_xfer_wr_offset_0,
	A_dc_xfer_wr_offset_1,
	A_dc_xfer_wr_offset_2,
	A_dc_wb_rd_addr_offset_0,
	A_dc_wb_rd_addr_offset_1,
	A_dc_wb_rd_addr_offset_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
input 	A_dc_xfer_wr_data_0;
output 	q_b_7;
output 	q_b_3;
input 	A_dc_xfer_wr_data_7;
output 	q_b_1;
input 	A_dc_xfer_wr_data_3;
output 	q_b_4;
output 	q_b_20;
output 	q_b_12;
output 	q_b_28;
output 	q_b_16;
output 	q_b_8;
output 	q_b_24;
output 	q_b_2;
output 	q_b_18;
output 	q_b_10;
output 	q_b_26;
output 	q_b_5;
output 	q_b_21;
output 	q_b_13;
output 	q_b_29;
output 	q_b_23;
output 	q_b_15;
output 	q_b_31;
output 	q_b_11;
output 	q_b_27;
output 	q_b_9;
output 	q_b_25;
output 	q_b_6;
output 	q_b_22;
output 	q_b_14;
output 	q_b_30;
output 	q_b_19;
input 	A_dc_xfer_wr_data_1;
output 	q_b_17;
input 	A_dc_xfer_wr_data_4;
input 	A_dc_xfer_wr_data_20;
input 	A_dc_xfer_wr_data_12;
input 	A_dc_xfer_wr_data_28;
input 	A_dc_xfer_wr_data_16;
input 	A_dc_xfer_wr_data_8;
input 	A_dc_xfer_wr_data_24;
input 	A_dc_xfer_wr_data_2;
input 	A_dc_xfer_wr_data_18;
input 	A_dc_xfer_wr_data_10;
input 	A_dc_xfer_wr_data_26;
input 	A_dc_xfer_wr_data_5;
input 	A_dc_xfer_wr_data_21;
input 	A_dc_xfer_wr_data_13;
input 	A_dc_xfer_wr_data_29;
input 	A_dc_xfer_wr_data_23;
input 	A_dc_xfer_wr_data_15;
input 	A_dc_xfer_wr_data_31;
input 	A_dc_xfer_wr_data_11;
input 	A_dc_xfer_wr_data_27;
input 	A_dc_xfer_wr_data_9;
input 	A_dc_xfer_wr_data_25;
input 	A_dc_xfer_wr_data_6;
input 	A_dc_xfer_wr_data_22;
input 	A_dc_xfer_wr_data_14;
input 	A_dc_xfer_wr_data_30;
input 	A_dc_xfer_wr_data_19;
input 	A_dc_xfer_wr_data_17;
input 	A_dc_xfer_wr_active;
input 	A_dc_wb_rd_en;
input 	A_dc_xfer_wr_offset_0;
input 	A_dc_xfer_wr_offset_1;
input 	A_dc_xfer_wr_offset_2;
input 	A_dc_wb_rd_addr_offset_0;
input 	A_dc_wb_rd_addr_offset_1;
input 	A_dc_wb_rd_addr_offset_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_4 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_dc_xfer_wr_data_31,A_dc_xfer_wr_data_30,A_dc_xfer_wr_data_29,A_dc_xfer_wr_data_28,A_dc_xfer_wr_data_27,A_dc_xfer_wr_data_26,A_dc_xfer_wr_data_25,A_dc_xfer_wr_data_24,A_dc_xfer_wr_data_23,A_dc_xfer_wr_data_22,A_dc_xfer_wr_data_21,A_dc_xfer_wr_data_20,
A_dc_xfer_wr_data_19,A_dc_xfer_wr_data_18,A_dc_xfer_wr_data_17,A_dc_xfer_wr_data_16,A_dc_xfer_wr_data_15,A_dc_xfer_wr_data_14,A_dc_xfer_wr_data_13,A_dc_xfer_wr_data_12,A_dc_xfer_wr_data_11,A_dc_xfer_wr_data_10,A_dc_xfer_wr_data_9,A_dc_xfer_wr_data_8,
A_dc_xfer_wr_data_7,A_dc_xfer_wr_data_6,A_dc_xfer_wr_data_5,A_dc_xfer_wr_data_4,A_dc_xfer_wr_data_3,A_dc_xfer_wr_data_2,A_dc_xfer_wr_data_1,A_dc_xfer_wr_data_0}),
	.wren_a(A_dc_xfer_wr_active),
	.rden_b(A_dc_wb_rd_en),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dc_xfer_wr_offset_2,A_dc_xfer_wr_offset_1,A_dc_xfer_wr_offset_0}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dc_wb_rd_addr_offset_2,A_dc_wb_rd_addr_offset_1,A_dc_wb_rd_addr_offset_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_4 (
	q_b,
	data_a,
	wren_a,
	rden_b,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	rden_b;
input 	[12:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_baj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.rden_b(rden_b),
	.address_a({address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_baj1 (
	q_b,
	data_a,
	wren_a,
	rden_b,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	rden_b;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 3;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 7;
defparam ram_block1a20.port_a_logical_ram_depth = 8;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 3;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 7;
defparam ram_block1a20.port_b_logical_ram_depth = 8;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 3;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 7;
defparam ram_block1a28.port_a_logical_ram_depth = 8;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 3;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 7;
defparam ram_block1a28.port_b_logical_ram_depth = 8;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 3;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 7;
defparam ram_block1a16.port_a_logical_ram_depth = 8;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 3;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 7;
defparam ram_block1a24.port_a_logical_ram_depth = 8;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 3;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 7;
defparam ram_block1a24.port_b_logical_ram_depth = 8;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 3;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 7;
defparam ram_block1a18.port_a_logical_ram_depth = 8;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 3;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 7;
defparam ram_block1a26.port_a_logical_ram_depth = 8;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 3;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 7;
defparam ram_block1a26.port_b_logical_ram_depth = 8;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 3;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 7;
defparam ram_block1a21.port_a_logical_ram_depth = 8;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 3;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 7;
defparam ram_block1a21.port_b_logical_ram_depth = 8;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 3;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 7;
defparam ram_block1a29.port_a_logical_ram_depth = 8;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 3;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 7;
defparam ram_block1a29.port_b_logical_ram_depth = 8;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 3;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 7;
defparam ram_block1a23.port_a_logical_ram_depth = 8;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 3;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 7;
defparam ram_block1a23.port_b_logical_ram_depth = 8;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 3;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 7;
defparam ram_block1a31.port_a_logical_ram_depth = 8;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 3;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 7;
defparam ram_block1a31.port_b_logical_ram_depth = 8;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 3;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 7;
defparam ram_block1a27.port_a_logical_ram_depth = 8;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 3;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 7;
defparam ram_block1a27.port_b_logical_ram_depth = 8;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 3;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 7;
defparam ram_block1a25.port_a_logical_ram_depth = 8;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 3;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 7;
defparam ram_block1a25.port_b_logical_ram_depth = 8;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 3;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 7;
defparam ram_block1a22.port_a_logical_ram_depth = 8;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 3;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 7;
defparam ram_block1a22.port_b_logical_ram_depth = 8;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 3;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 7;
defparam ram_block1a30.port_a_logical_ram_depth = 8;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 3;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 7;
defparam ram_block1a30.port_b_logical_ram_depth = 8;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 3;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 7;
defparam ram_block1a19.port_a_logical_ram_depth = 8;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_dc_victim_module:Qsys_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 3;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 7;
defparam ram_block1a17.port_a_logical_ram_depth = 8;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_ic_data_module (
	q_b_5,
	q_b_3,
	q_b_1,
	q_b_4,
	q_b_2,
	q_b_28,
	q_b_30,
	q_b_31,
	q_b_27,
	q_b_29,
	q_b_0,
	q_b_23,
	q_b_25,
	q_b_26,
	q_b_22,
	q_b_24,
	q_b_16,
	q_b_15,
	q_b_13,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_8,
	q_b_18,
	q_b_17,
	q_b_21,
	q_b_6,
	q_b_20,
	q_b_19,
	q_b_9,
	q_b_7,
	ic_fill_line_6,
	ic_fill_line_5,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_0,
	F_stall,
	ic_fill_dp_offset_0,
	ic_fill_dp_offset_1,
	ic_fill_dp_offset_2,
	i_readdatavalid_d1,
	F_ic_tag_rd_addr_nxt_6,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_0,
	i_readdata_d1_5,
	F_ic_data_rd_addr_nxt_0,
	F_ic_data_rd_addr_nxt_1,
	F_ic_data_rd_addr_nxt_2,
	i_readdata_d1_3,
	i_readdata_d1_1,
	i_readdata_d1_4,
	i_readdata_d1_2,
	i_readdata_d1_28,
	i_readdata_d1_30,
	i_readdata_d1_31,
	i_readdata_d1_27,
	i_readdata_d1_29,
	i_readdata_d1_0,
	i_readdata_d1_23,
	i_readdata_d1_25,
	i_readdata_d1_26,
	i_readdata_d1_22,
	i_readdata_d1_24,
	i_readdata_d1_16,
	i_readdata_d1_15,
	i_readdata_d1_13,
	i_readdata_d1_14,
	i_readdata_d1_12,
	i_readdata_d1_11,
	i_readdata_d1_10,
	i_readdata_d1_8,
	i_readdata_d1_18,
	i_readdata_d1_17,
	i_readdata_d1_21,
	i_readdata_d1_6,
	i_readdata_d1_20,
	i_readdata_d1_19,
	i_readdata_d1_9,
	i_readdata_d1_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_3;
output 	q_b_1;
output 	q_b_4;
output 	q_b_2;
output 	q_b_28;
output 	q_b_30;
output 	q_b_31;
output 	q_b_27;
output 	q_b_29;
output 	q_b_0;
output 	q_b_23;
output 	q_b_25;
output 	q_b_26;
output 	q_b_22;
output 	q_b_24;
output 	q_b_16;
output 	q_b_15;
output 	q_b_13;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_8;
output 	q_b_18;
output 	q_b_17;
output 	q_b_21;
output 	q_b_6;
output 	q_b_20;
output 	q_b_19;
output 	q_b_9;
output 	q_b_7;
input 	ic_fill_line_6;
input 	ic_fill_line_5;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_0;
input 	F_stall;
input 	ic_fill_dp_offset_0;
input 	ic_fill_dp_offset_1;
input 	ic_fill_dp_offset_2;
input 	i_readdatavalid_d1;
input 	F_ic_tag_rd_addr_nxt_6;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_0;
input 	i_readdata_d1_5;
input 	F_ic_data_rd_addr_nxt_0;
input 	F_ic_data_rd_addr_nxt_1;
input 	F_ic_data_rd_addr_nxt_2;
input 	i_readdata_d1_3;
input 	i_readdata_d1_1;
input 	i_readdata_d1_4;
input 	i_readdata_d1_2;
input 	i_readdata_d1_28;
input 	i_readdata_d1_30;
input 	i_readdata_d1_31;
input 	i_readdata_d1_27;
input 	i_readdata_d1_29;
input 	i_readdata_d1_0;
input 	i_readdata_d1_23;
input 	i_readdata_d1_25;
input 	i_readdata_d1_26;
input 	i_readdata_d1_22;
input 	i_readdata_d1_24;
input 	i_readdata_d1_16;
input 	i_readdata_d1_15;
input 	i_readdata_d1_13;
input 	i_readdata_d1_14;
input 	i_readdata_d1_12;
input 	i_readdata_d1_11;
input 	i_readdata_d1_10;
input 	i_readdata_d1_8;
input 	i_readdata_d1_18;
input 	i_readdata_d1_17;
input 	i_readdata_d1_21;
input 	i_readdata_d1_6;
input 	i_readdata_d1_20;
input 	i_readdata_d1_19;
input 	i_readdata_d1_9;
input 	i_readdata_d1_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_5 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({gnd,gnd,gnd,ic_fill_line_6,ic_fill_line_5,ic_fill_line_4,ic_fill_line_3,ic_fill_line_2,ic_fill_line_1,ic_fill_line_0,ic_fill_dp_offset_2,ic_fill_dp_offset_1,ic_fill_dp_offset_0}),
	.rden_b(F_stall),
	.wren_a(i_readdatavalid_d1),
	.address_b({F_ic_tag_rd_addr_nxt_6,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0,F_ic_data_rd_addr_nxt_2,F_ic_data_rd_addr_nxt_1,F_ic_data_rd_addr_nxt_0}),
	.data_a({i_readdata_d1_31,i_readdata_d1_30,i_readdata_d1_29,i_readdata_d1_28,i_readdata_d1_27,i_readdata_d1_26,i_readdata_d1_25,i_readdata_d1_24,i_readdata_d1_23,i_readdata_d1_22,i_readdata_d1_21,i_readdata_d1_20,i_readdata_d1_19,i_readdata_d1_18,i_readdata_d1_17,i_readdata_d1_16,
i_readdata_d1_15,i_readdata_d1_14,i_readdata_d1_13,i_readdata_d1_12,i_readdata_d1_11,i_readdata_d1_10,i_readdata_d1_9,i_readdata_d1_8,i_readdata_d1_7,i_readdata_d1_6,i_readdata_d1_5,i_readdata_d1_4,i_readdata_d1_3,i_readdata_d1_2,i_readdata_d1_1,i_readdata_d1_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_5 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[12:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[9:0] address_b;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_spj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.address_b({address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_spj1 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[9:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[9:0] address_b;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 10;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 1023;
defparam ram_block1a5.port_a_logical_ram_depth = 1024;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 10;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 1023;
defparam ram_block1a5.port_b_logical_ram_depth = 1024;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 10;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 1023;
defparam ram_block1a3.port_a_logical_ram_depth = 1024;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 10;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 1023;
defparam ram_block1a3.port_b_logical_ram_depth = 1024;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 10;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 1023;
defparam ram_block1a1.port_a_logical_ram_depth = 1024;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 10;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 1023;
defparam ram_block1a1.port_b_logical_ram_depth = 1024;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 10;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 1023;
defparam ram_block1a4.port_a_logical_ram_depth = 1024;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 10;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 1023;
defparam ram_block1a4.port_b_logical_ram_depth = 1024;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 10;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 1023;
defparam ram_block1a2.port_a_logical_ram_depth = 1024;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 10;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 1023;
defparam ram_block1a2.port_b_logical_ram_depth = 1024;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 10;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 1023;
defparam ram_block1a28.port_a_logical_ram_depth = 1024;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 10;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 1023;
defparam ram_block1a28.port_b_logical_ram_depth = 1024;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 10;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 1023;
defparam ram_block1a30.port_a_logical_ram_depth = 1024;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 10;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 1023;
defparam ram_block1a30.port_b_logical_ram_depth = 1024;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 10;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 1023;
defparam ram_block1a31.port_a_logical_ram_depth = 1024;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 10;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 1023;
defparam ram_block1a31.port_b_logical_ram_depth = 1024;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 10;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 1023;
defparam ram_block1a27.port_a_logical_ram_depth = 1024;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 10;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 1023;
defparam ram_block1a27.port_b_logical_ram_depth = 1024;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 10;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 1023;
defparam ram_block1a29.port_a_logical_ram_depth = 1024;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 10;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 1023;
defparam ram_block1a29.port_b_logical_ram_depth = 1024;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 10;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 1023;
defparam ram_block1a0.port_a_logical_ram_depth = 1024;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 10;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 1023;
defparam ram_block1a0.port_b_logical_ram_depth = 1024;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 10;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 1023;
defparam ram_block1a23.port_a_logical_ram_depth = 1024;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 10;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 1023;
defparam ram_block1a23.port_b_logical_ram_depth = 1024;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 10;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 1023;
defparam ram_block1a25.port_a_logical_ram_depth = 1024;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 10;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 1023;
defparam ram_block1a25.port_b_logical_ram_depth = 1024;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 10;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 1023;
defparam ram_block1a26.port_a_logical_ram_depth = 1024;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 10;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 1023;
defparam ram_block1a26.port_b_logical_ram_depth = 1024;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 10;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 1023;
defparam ram_block1a22.port_a_logical_ram_depth = 1024;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 10;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 1023;
defparam ram_block1a22.port_b_logical_ram_depth = 1024;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 10;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 1023;
defparam ram_block1a24.port_a_logical_ram_depth = 1024;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 10;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 1023;
defparam ram_block1a24.port_b_logical_ram_depth = 1024;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 10;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 1023;
defparam ram_block1a16.port_a_logical_ram_depth = 1024;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 10;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 1023;
defparam ram_block1a16.port_b_logical_ram_depth = 1024;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 10;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 1023;
defparam ram_block1a15.port_a_logical_ram_depth = 1024;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 10;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 1023;
defparam ram_block1a15.port_b_logical_ram_depth = 1024;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 10;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 1023;
defparam ram_block1a13.port_a_logical_ram_depth = 1024;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 10;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 1023;
defparam ram_block1a13.port_b_logical_ram_depth = 1024;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 10;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 1023;
defparam ram_block1a14.port_a_logical_ram_depth = 1024;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 10;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 1023;
defparam ram_block1a14.port_b_logical_ram_depth = 1024;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 10;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 1023;
defparam ram_block1a12.port_a_logical_ram_depth = 1024;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 10;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 1023;
defparam ram_block1a12.port_b_logical_ram_depth = 1024;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 10;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 1023;
defparam ram_block1a11.port_a_logical_ram_depth = 1024;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 10;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 1023;
defparam ram_block1a11.port_b_logical_ram_depth = 1024;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 10;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 1023;
defparam ram_block1a10.port_a_logical_ram_depth = 1024;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 10;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 1023;
defparam ram_block1a10.port_b_logical_ram_depth = 1024;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 10;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 1023;
defparam ram_block1a8.port_a_logical_ram_depth = 1024;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 10;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 1023;
defparam ram_block1a8.port_b_logical_ram_depth = 1024;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 10;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 1023;
defparam ram_block1a18.port_a_logical_ram_depth = 1024;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 10;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 1023;
defparam ram_block1a18.port_b_logical_ram_depth = 1024;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 10;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 1023;
defparam ram_block1a17.port_a_logical_ram_depth = 1024;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 10;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 1023;
defparam ram_block1a17.port_b_logical_ram_depth = 1024;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 10;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 1023;
defparam ram_block1a21.port_a_logical_ram_depth = 1024;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 10;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 1023;
defparam ram_block1a21.port_b_logical_ram_depth = 1024;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 10;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 1023;
defparam ram_block1a6.port_a_logical_ram_depth = 1024;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 10;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 1023;
defparam ram_block1a6.port_b_logical_ram_depth = 1024;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 10;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 1023;
defparam ram_block1a20.port_a_logical_ram_depth = 1024;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 10;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 1023;
defparam ram_block1a20.port_b_logical_ram_depth = 1024;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 10;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 1023;
defparam ram_block1a19.port_a_logical_ram_depth = 1024;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 10;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 1023;
defparam ram_block1a19.port_b_logical_ram_depth = 1024;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 10;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 1023;
defparam ram_block1a9.port_a_logical_ram_depth = 1024;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 10;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 1023;
defparam ram_block1a9.port_b_logical_ram_depth = 1024;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_data_module:Qsys_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 10;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 1023;
defparam ram_block1a7.port_a_logical_ram_depth = 1024;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 10;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 1023;
defparam ram_block1a7.port_b_logical_ram_depth = 1024;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_ic_tag_module (
	q_b_2,
	q_b_0,
	q_b_1,
	q_b_3,
	q_b_4,
	q_b_10,
	q_b_12,
	q_b_9,
	q_b_11,
	ic_fill_valid_bits_5,
	ic_fill_valid_bits_7,
	ic_fill_valid_bits_4,
	q_b_6,
	q_b_8,
	q_b_5,
	q_b_7,
	ic_fill_valid_bits_6,
	ic_fill_valid_bits_1,
	ic_fill_valid_bits_3,
	ic_fill_valid_bits_0,
	ic_fill_valid_bits_2,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	F_stall,
	F_ic_tag_rd_addr_nxt_6,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_0,
	ic_tag_wren,
	ic_tag_wraddress_0,
	ic_tag_wraddress_1,
	ic_tag_wraddress_2,
	ic_tag_wraddress_3,
	ic_tag_wraddress_4,
	ic_tag_wraddress_5,
	ic_tag_wraddress_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_2;
output 	q_b_0;
output 	q_b_1;
output 	q_b_3;
output 	q_b_4;
output 	q_b_10;
output 	q_b_12;
output 	q_b_9;
output 	q_b_11;
input 	ic_fill_valid_bits_5;
input 	ic_fill_valid_bits_7;
input 	ic_fill_valid_bits_4;
output 	q_b_6;
output 	q_b_8;
output 	q_b_5;
output 	q_b_7;
input 	ic_fill_valid_bits_6;
input 	ic_fill_valid_bits_1;
input 	ic_fill_valid_bits_3;
input 	ic_fill_valid_bits_0;
input 	ic_fill_valid_bits_2;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	F_stall;
input 	F_ic_tag_rd_addr_nxt_6;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_0;
input 	ic_tag_wren;
input 	ic_tag_wraddress_0;
input 	ic_tag_wraddress_1;
input 	ic_tag_wraddress_2;
input 	ic_tag_wraddress_3;
input 	ic_tag_wraddress_4;
input 	ic_tag_wraddress_5;
input 	ic_tag_wraddress_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_6 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_fill_valid_bits_7,ic_fill_valid_bits_6,ic_fill_valid_bits_5,ic_fill_valid_bits_4,ic_fill_valid_bits_3,ic_fill_valid_bits_2,ic_fill_valid_bits_1,ic_fill_valid_bits_0,ic_fill_tag_4,ic_fill_tag_3,ic_fill_tag_2,
ic_fill_tag_1,ic_fill_tag_0}),
	.rden_b(F_stall),
	.address_b({gnd,gnd,gnd,F_ic_tag_rd_addr_nxt_6,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0}),
	.wren_a(ic_tag_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,ic_tag_wraddress_6,ic_tag_wraddress_5,ic_tag_wraddress_4,ic_tag_wraddress_3,ic_tag_wraddress_2,ic_tag_wraddress_1,ic_tag_wraddress_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_6 (
	q_b,
	data_a,
	rden_b,
	address_b,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	rden_b;
input 	[9:0] address_b;
input 	wren_a;
input 	[12:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_mgo1 auto_generated(
	.q_b({q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.rden_b(rden_b),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_mgo1 (
	q_b,
	data_a,
	rden_b,
	address_b,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[12:0] q_b;
input 	[12:0] data_a;
input 	rden_b;
input 	[6:0] address_b;
input 	wren_a;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 13;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 13;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "F8D03CE85CB189A866F33435CC960198";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 13;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 13;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "B57EB627EACE9E3DB4E2FBAE751F1E7B";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 13;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 13;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "C3FCF92EBBCC2B6A198D03846DA98D04";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 13;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 13;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "73D9443D590D805932C19C540815BA17";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 13;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 13;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "9EC4F7C0395A71D9C7150B3DCE44583B";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 13;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 13;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "C78EA19A15635D63B7985C4CB0BBC968";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 13;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 13;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "EE1F708F423E6F94E0EC38012A3EDBCD";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 13;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 13;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "09415291511A5F780D6F81A0DC328FD6";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 13;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 13;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "617B4B0894A9F3BD864713E5C66BCE07";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 13;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 13;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "F440ECAC4FFB1F094F2996DA16385CF2";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 13;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 13;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "416DB8FE334D30A9F63F2250392C148C";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 13;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 13;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "9BF506141D38FED27209A6A81568A156";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_ic_tag_module:Qsys_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_mgo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 13;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 13;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "92357571045DDED040349E904F8351BF";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_mult_cell (
	Add0,
	Add01,
	Add02,
	Add03,
	Add04,
	Add05,
	Add06,
	Add07,
	Add08,
	Add09,
	Add010,
	Add011,
	Add012,
	Add013,
	Add014,
	Add015,
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	r_sync_rst,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	Add0;
output 	Add01;
output 	Add02;
output 	Add03;
output 	Add04;
output 	Add05;
output 	Add06;
output 	Add07;
output 	Add08;
output 	Add09;
output 	Add010;
output 	Add011;
output 	Add012;
output 	Add013;
output 	Add014;
output 	Add015;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	r_sync_rst;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ;
wire \Add0~2 ;
wire \Add0~6 ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~18 ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~30 ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~50 ;
wire \Add0~54 ;
wire \Add0~58 ;


Qsys_system_altera_mult_add the_altmult_add_part_1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_16(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.data_out_wire_29(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.data_out_wire_28(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.data_out_wire_27(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.data_out_wire_30(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.data_out_wire_26(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.data_out_wire_25(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.data_out_wire_19(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.data_out_wire_17(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.data_out_wire_22(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.data_out_wire_21(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.data_out_wire_20(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.data_out_wire_18(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.data_out_wire_24(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.data_out_wire_23(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.data_out_wire_31(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.clk_clk(clk_clk));

Qsys_system_altera_mult_add_1 the_altmult_add_part_2(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_0(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_13(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_12(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_11(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_14(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_10(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_9(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_3(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_1(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_6(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_5(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_4(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_2(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_8(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_7(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_15(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.clk_clk(clk_clk));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add0),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add01),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add02),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add03),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add04),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add05),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add06),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add07),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add08),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add09),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add010),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add011),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add012),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add013),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add014),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add015),
	.cout(),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

endmodule

module Qsys_system_altera_mult_add (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	r_sync_rst,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_16,
	data_out_wire_29,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_30,
	data_out_wire_26,
	data_out_wire_25,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_22,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_18,
	data_out_wire_24,
	data_out_wire_23,
	data_out_wire_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	r_sync_rst;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_16;
output 	data_out_wire_29;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_30;
output 	data_out_wire_26;
output 	data_out_wire_25;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_22;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_18;
output 	data_out_wire_24;
output 	data_out_wire_23;
output 	data_out_wire_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altera_mult_add_ujt2 auto_generated(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_31(data_out_wire_31),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_altera_mult_add_ujt2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	r_sync_rst,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_16,
	data_out_wire_29,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_30,
	data_out_wire_26,
	data_out_wire_25,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_22,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_18,
	data_out_wire_24,
	data_out_wire_23,
	data_out_wire_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	r_sync_rst;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_16;
output 	data_out_wire_29;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_30;
output 	data_out_wire_26;
output 	data_out_wire_25;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_22;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_18;
output 	data_out_wire_24;
output 	data_out_wire_23;
output 	data_out_wire_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altera_mult_add_rtl_1 altera_mult_add_rtl1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_31(data_out_wire_31),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_altera_mult_add_rtl_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	r_sync_rst,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_16,
	data_out_wire_29,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_30,
	data_out_wire_26,
	data_out_wire_25,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_22,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_18,
	data_out_wire_24,
	data_out_wire_23,
	data_out_wire_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	r_sync_rst;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_16;
output 	data_out_wire_29;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_30;
output 	data_out_wire_26;
output 	data_out_wire_25;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_22;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_18;
output 	data_out_wire_24;
output 	data_out_wire_23;
output 	data_out_wire_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_ama_multiplier_function multiplier_block(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_31(data_out_wire_31),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_ama_multiplier_function (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	r_sync_rst,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_16,
	data_out_wire_29,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_30,
	data_out_wire_26,
	data_out_wire_25,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_22,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_18,
	data_out_wire_24,
	data_out_wire_23,
	data_out_wire_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	r_sync_rst;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_16;
output 	data_out_wire_29;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_30;
output 	data_out_wire_26;
output 	data_out_wire_25;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_22;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_18;
output 	data_out_wire_24;
output 	data_out_wire_23;
output 	data_out_wire_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \data_out_wire_0[16] ;
wire \data_out_wire_0[17] ;
wire \data_out_wire_0[18] ;
wire \data_out_wire_0[19] ;
wire \data_out_wire_0[20] ;
wire \data_out_wire_0[21] ;
wire \data_out_wire_0[22] ;
wire \data_out_wire_0[23] ;
wire \data_out_wire_0[24] ;
wire \data_out_wire_0[25] ;
wire \data_out_wire_0[26] ;
wire \data_out_wire_0[27] ;
wire \data_out_wire_0[28] ;
wire \data_out_wire_0[29] ;
wire \data_out_wire_0[30] ;
wire \data_out_wire_0[31] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \data_out_wire_0[16]  = \Mult0~mac_RESULTA_bus [16];
assign \data_out_wire_0[17]  = \Mult0~mac_RESULTA_bus [17];
assign \data_out_wire_0[18]  = \Mult0~mac_RESULTA_bus [18];
assign \data_out_wire_0[19]  = \Mult0~mac_RESULTA_bus [19];
assign \data_out_wire_0[20]  = \Mult0~mac_RESULTA_bus [20];
assign \data_out_wire_0[21]  = \Mult0~mac_RESULTA_bus [21];
assign \data_out_wire_0[22]  = \Mult0~mac_RESULTA_bus [22];
assign \data_out_wire_0[23]  = \Mult0~mac_RESULTA_bus [23];
assign \data_out_wire_0[24]  = \Mult0~mac_RESULTA_bus [24];
assign \data_out_wire_0[25]  = \Mult0~mac_RESULTA_bus [25];
assign \data_out_wire_0[26]  = \Mult0~mac_RESULTA_bus [26];
assign \data_out_wire_0[27]  = \Mult0~mac_RESULTA_bus [27];
assign \data_out_wire_0[28]  = \Mult0~mac_RESULTA_bus [28];
assign \data_out_wire_0[29]  = \Mult0~mac_RESULTA_bus [29];
assign \data_out_wire_0[30]  = \Mult0~mac_RESULTA_bus [30];
assign \data_out_wire_0[31]  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [63];

Qsys_system_ama_register_function_12 multiplier_register_block_0(
	.data_in({gnd,gnd,\data_out_wire_0[31] ,\data_out_wire_0[30] ,\data_out_wire_0[29] ,\data_out_wire_0[28] ,\data_out_wire_0[27] ,\data_out_wire_0[26] ,\data_out_wire_0[25] ,\data_out_wire_0[24] ,\data_out_wire_0[23] ,\data_out_wire_0[22] ,\data_out_wire_0[21] ,
\data_out_wire_0[20] ,\data_out_wire_0[19] ,\data_out_wire_0[18] ,\data_out_wire_0[17] ,\data_out_wire_0[16] ,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,
\data_out_wire_0[8] ,\data_out_wire_0[7] ,\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,r_sync_rst}),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_31(data_out_wire_31),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src2_15,A_mul_src2_14,A_mul_src2_13,A_mul_src2_12,A_mul_src2_11,A_mul_src2_10,A_mul_src2_9,A_mul_src2_8,A_mul_src2_7,A_mul_src2_6,A_mul_src2_5,A_mul_src2_4,A_mul_src2_3,A_mul_src2_2,A_mul_src2_1,A_mul_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src1_15,A_mul_src1_14,A_mul_src1_13,A_mul_src1_12,A_mul_src1_11,A_mul_src1_10,A_mul_src1_9,A_mul_src1_8,A_mul_src1_7,A_mul_src1_6,A_mul_src1_5,A_mul_src1_4,A_mul_src1_3,A_mul_src1_2,A_mul_src1_1,A_mul_src1_0}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module Qsys_system_ama_register_function_12 (
	data_in,
	aclr,
	data_out_wire_4,
	data_out_wire_0,
	data_out_wire_2,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_13,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_16,
	data_out_wire_29,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_30,
	data_out_wire_26,
	data_out_wire_25,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_22,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_18,
	data_out_wire_24,
	data_out_wire_23,
	data_out_wire_31,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
output 	data_out_wire_4;
output 	data_out_wire_0;
output 	data_out_wire_2;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_13;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_16;
output 	data_out_wire_29;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_30;
output 	data_out_wire_26;
output 	data_out_wire_25;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_22;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_18;
output 	data_out_wire_24;
output 	data_out_wire_23;
output 	data_out_wire_31;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[16] (
	.clk(clock[0]),
	.d(data_in[16]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_16),
	.prn(vcc));
defparam \data_out_wire[16] .is_wysiwyg = "true";
defparam \data_out_wire[16] .power_up = "low";

dffeas \data_out_wire[29] (
	.clk(clock[0]),
	.d(data_in[29]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_29),
	.prn(vcc));
defparam \data_out_wire[29] .is_wysiwyg = "true";
defparam \data_out_wire[29] .power_up = "low";

dffeas \data_out_wire[28] (
	.clk(clock[0]),
	.d(data_in[28]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_28),
	.prn(vcc));
defparam \data_out_wire[28] .is_wysiwyg = "true";
defparam \data_out_wire[28] .power_up = "low";

dffeas \data_out_wire[27] (
	.clk(clock[0]),
	.d(data_in[27]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_27),
	.prn(vcc));
defparam \data_out_wire[27] .is_wysiwyg = "true";
defparam \data_out_wire[27] .power_up = "low";

dffeas \data_out_wire[30] (
	.clk(clock[0]),
	.d(data_in[30]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_30),
	.prn(vcc));
defparam \data_out_wire[30] .is_wysiwyg = "true";
defparam \data_out_wire[30] .power_up = "low";

dffeas \data_out_wire[26] (
	.clk(clock[0]),
	.d(data_in[26]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_26),
	.prn(vcc));
defparam \data_out_wire[26] .is_wysiwyg = "true";
defparam \data_out_wire[26] .power_up = "low";

dffeas \data_out_wire[25] (
	.clk(clock[0]),
	.d(data_in[25]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_25),
	.prn(vcc));
defparam \data_out_wire[25] .is_wysiwyg = "true";
defparam \data_out_wire[25] .power_up = "low";

dffeas \data_out_wire[19] (
	.clk(clock[0]),
	.d(data_in[19]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_19),
	.prn(vcc));
defparam \data_out_wire[19] .is_wysiwyg = "true";
defparam \data_out_wire[19] .power_up = "low";

dffeas \data_out_wire[17] (
	.clk(clock[0]),
	.d(data_in[17]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_17),
	.prn(vcc));
defparam \data_out_wire[17] .is_wysiwyg = "true";
defparam \data_out_wire[17] .power_up = "low";

dffeas \data_out_wire[22] (
	.clk(clock[0]),
	.d(data_in[22]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_22),
	.prn(vcc));
defparam \data_out_wire[22] .is_wysiwyg = "true";
defparam \data_out_wire[22] .power_up = "low";

dffeas \data_out_wire[21] (
	.clk(clock[0]),
	.d(data_in[21]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_21),
	.prn(vcc));
defparam \data_out_wire[21] .is_wysiwyg = "true";
defparam \data_out_wire[21] .power_up = "low";

dffeas \data_out_wire[20] (
	.clk(clock[0]),
	.d(data_in[20]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_20),
	.prn(vcc));
defparam \data_out_wire[20] .is_wysiwyg = "true";
defparam \data_out_wire[20] .power_up = "low";

dffeas \data_out_wire[18] (
	.clk(clock[0]),
	.d(data_in[18]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_18),
	.prn(vcc));
defparam \data_out_wire[18] .is_wysiwyg = "true";
defparam \data_out_wire[18] .power_up = "low";

dffeas \data_out_wire[24] (
	.clk(clock[0]),
	.d(data_in[24]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_24),
	.prn(vcc));
defparam \data_out_wire[24] .is_wysiwyg = "true";
defparam \data_out_wire[24] .power_up = "low";

dffeas \data_out_wire[23] (
	.clk(clock[0]),
	.d(data_in[23]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_23),
	.prn(vcc));
defparam \data_out_wire[23] .is_wysiwyg = "true";
defparam \data_out_wire[23] .power_up = "low";

dffeas \data_out_wire[31] (
	.clk(clock[0]),
	.d(data_in[31]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_31),
	.prn(vcc));
defparam \data_out_wire[31] .is_wysiwyg = "true";
defparam \data_out_wire[31] .power_up = "low";

endmodule

module Qsys_system_altera_mult_add_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	r_sync_rst,
	data_out_wire_0,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_14,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_2,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	r_sync_rst;
output 	data_out_wire_0;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_14;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_2;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altera_mult_add_0kt2 auto_generated(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_15(data_out_wire_15),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_altera_mult_add_0kt2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	r_sync_rst,
	data_out_wire_0,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_14,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_2,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	r_sync_rst;
output 	data_out_wire_0;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_14;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_2;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altera_mult_add_rtl_2 altera_mult_add_rtl1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_15(data_out_wire_15),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_altera_mult_add_rtl_2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	r_sync_rst,
	data_out_wire_0,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_14,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_2,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	r_sync_rst;
output 	data_out_wire_0;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_14;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_2;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_ama_multiplier_function_1 multiplier_block(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.r_sync_rst(r_sync_rst),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_15(data_out_wire_15),
	.clk_clk(clk_clk));

endmodule

module Qsys_system_ama_multiplier_function_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	r_sync_rst,
	data_out_wire_0,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_14,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_2,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	r_sync_rst;
output 	data_out_wire_0;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_14;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_2;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;
wire \Mult0~40 ;
wire \Mult0~41 ;
wire \Mult0~42 ;
wire \Mult0~43 ;
wire \Mult0~44 ;
wire \Mult0~45 ;
wire \Mult0~46 ;
wire \Mult0~47 ;
wire \Mult0~48 ;
wire \Mult0~49 ;
wire \Mult0~50 ;
wire \Mult0~51 ;
wire \Mult0~52 ;
wire \Mult0~53 ;
wire \Mult0~54 ;
wire \Mult0~55 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [16];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [17];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [18];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [19];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [20];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [21];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [22];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [23];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [24];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [25];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [26];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [27];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [28];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [29];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [30];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~40  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~41  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~42  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~43  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~44  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~45  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~46  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~47  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~48  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~49  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~50  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~51  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~52  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~53  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~54  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~55  = \Mult0~mac_RESULTA_bus [63];

Qsys_system_ama_register_function_31 multiplier_register_block_0(
	.data_in({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,\data_out_wire_0[8] ,\data_out_wire_0[7] ,
\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,r_sync_rst}),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_15(data_out_wire_15),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src2_15,A_mul_src2_14,A_mul_src2_13,A_mul_src2_12,A_mul_src2_11,A_mul_src2_10,A_mul_src2_9,A_mul_src2_8,A_mul_src2_7,A_mul_src2_6,A_mul_src2_5,A_mul_src2_4,A_mul_src2_3,A_mul_src2_2,A_mul_src2_1,A_mul_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src1_31,A_mul_src1_30,A_mul_src1_29,A_mul_src1_28,A_mul_src1_27,A_mul_src1_26,A_mul_src1_25,A_mul_src1_24,A_mul_src1_23,A_mul_src1_22,A_mul_src1_21,A_mul_src1_20,A_mul_src1_19,A_mul_src1_18,A_mul_src1_17,A_mul_src1_16}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module Qsys_system_ama_register_function_31 (
	data_in,
	aclr,
	data_out_wire_0,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_14,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_2,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_15,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
output 	data_out_wire_0;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_14;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_2;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_15;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci (
	readdata_4,
	readdata_20,
	readdata_12,
	readdata_28,
	readdata_16,
	readdata_8,
	readdata_24,
	readdata_2,
	readdata_18,
	readdata_10,
	readdata_26,
	readdata_5,
	readdata_21,
	readdata_13,
	readdata_29,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_11,
	readdata_27,
	readdata_9,
	readdata_25,
	readdata_6,
	readdata_22,
	readdata_14,
	readdata_30,
	readdata_3,
	readdata_19,
	readdata_17,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_write,
	r_sync_rst,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	WideOr1,
	rf_source_valid,
	hbreak_enabled,
	jtag_break,
	address_nxt,
	oci_single_step_mode,
	r_early_rst,
	writedata_nxt,
	debugaccess_nxt,
	byteenable_nxt,
	oci_ienable_0,
	oci_ienable_1,
	readdata_0,
	resetrequest,
	readdata_1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_4;
output 	readdata_20;
output 	readdata_12;
output 	readdata_28;
output 	readdata_16;
output 	readdata_8;
output 	readdata_24;
output 	readdata_2;
output 	readdata_18;
output 	readdata_10;
output 	readdata_26;
output 	readdata_5;
output 	readdata_21;
output 	readdata_13;
output 	readdata_29;
output 	readdata_7;
output 	readdata_23;
output 	readdata_15;
output 	readdata_31;
output 	readdata_11;
output 	readdata_27;
output 	readdata_9;
output 	readdata_25;
output 	readdata_6;
output 	readdata_22;
output 	readdata_14;
output 	readdata_30;
output 	readdata_3;
output 	readdata_19;
output 	readdata_17;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	d_write;
input 	r_sync_rst;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	WideOr1;
input 	rf_source_valid;
input 	hbreak_enabled;
output 	jtag_break;
input 	[8:0] address_nxt;
output 	oci_single_step_mode;
input 	r_early_rst;
input 	[31:0] writedata_nxt;
input 	debugaccess_nxt;
input 	[3:0] byteenable_nxt;
output 	oci_ienable_0;
output 	oci_ienable_1;
output 	readdata_0;
output 	resetrequest;
output 	readdata_1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ;
wire \write~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ;
wire \read~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \address[0]~q ;
wire \address[3]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \address[4]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal0~1_combout ;
wire \debugaccess~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ;
wire \byteenable[0]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ;
wire \writedata[3]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal1~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ;
wire \writedata[16]~q ;
wire \byteenable[2]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ;
wire \writedata[4]~q ;
wire \writedata[26]~q ;
wire \writedata[27]~q ;
wire \writedata[25]~q ;
wire \writedata[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[21]~q ;
wire \writedata[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \byteenable[1]~q ;
wire \writedata[28]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \writedata[10]~q ;
wire \writedata[5]~q ;
wire \writedata[13]~q ;
wire \writedata[29]~q ;
wire \writedata[7]~q ;
wire \writedata[23]~q ;
wire \writedata[15]~q ;
wire \writedata[31]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ;
wire \writedata[11]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \writedata[6]~q ;
wire \writedata[22]~q ;
wire \the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \writedata[30]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ;
wire \address[8]~q ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata[0]~0_combout ;
wire \readdata[0]~1_combout ;
wire \readdata~2_combout ;
wire \readdata~5_combout ;


Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper(
	.break_readreg_0(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ),
	.break_readreg_2(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_20(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ),
	.break_readreg_24(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_26(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_27(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_25(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_17(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ),
	.break_readreg_21(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ),
	.MonDReg_21(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_18(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_5(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_29(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ),
	.MonDReg_30(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_30(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_22(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ),
	.MonDReg_22(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ),
	.break_readreg_6(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ),
	.MonDReg_6(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ),
	.break_readreg_15(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ),
	.MonDReg_23(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_10(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_13(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_7(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ),
	.break_readreg_7(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_8(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_14(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_13(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_11(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.MonDReg_0(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ),
	.hbreak_enabled(hbreak_enabled),
	.monitor_ready(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.jdo_0(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ),
	.ir_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.jdo_35(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_b(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_34(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.MonDReg_2(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_27(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_28(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_26(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.MonDReg_3(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_29(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ),
	.MonDReg_16(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ),
	.monitor_error(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.MonDReg_4(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.jdo_16(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ),
	.jdo_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.MonDReg_5(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ),
	.resetlatch(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ),
	.jdo_8(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.MonDReg_15(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_12(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_8(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_11(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_9(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_14(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ),
	.jdo_9(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_15(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_11(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_13(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_10(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci_break the_Qsys_system_nios2_qsys_0_nios2_oci_break(
	.break_readreg_0(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_20(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_24(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_26(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_27(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_25(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_17(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_21(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_5(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_22(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_6(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_8(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_14(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_13(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_11(\the_Qsys_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ),
	.jdo_0(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ),
	.ir_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.jdo_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_27(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_28(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_26(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_2(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_29(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_6(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.jdo_16(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.jdo_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.jdo_7(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.jdo_8(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_9(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_15(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_11(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_13(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_10(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_nios2_avalon_reg the_Qsys_system_nios2_qsys_0_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.oci_single_step_mode1(oci_single_step_mode),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.Equal0(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal0~1_combout ),
	.debugaccess(\debugaccess~q ),
	.take_action_ocireg(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.writedata_3(\writedata[3]~q ),
	.writedata_1(\writedata[1]~q ),
	.oci_ienable_0(oci_ienable_0),
	.oci_ienable_1(oci_ienable_1),
	.Equal1(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal1~0_combout ),
	.oci_reg_readdata(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_nios2_ocimem the_Qsys_system_nios2_qsys_0_nios2_ocimem(
	.MonDReg_1(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ),
	.q_a_0(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.MonDReg_20(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_24(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ),
	.q_a_3(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.MonDReg_26(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_27(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_25(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_17(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ),
	.q_a_16(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.MonDReg_21(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ),
	.q_a_20(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_24(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_4(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.MonDReg_28(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_30(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ),
	.q_a_26(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_27(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_25(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_17(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.MonDReg_22(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ),
	.q_a_21(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_12(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_8(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_5(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_13(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_7(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_9(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_6(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.MonDReg_6(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_23(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_10(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_13(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_7(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.jdo_35(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_b(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_34(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_no_action_ocimem_a(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.debugaccess(\debugaccess~q ),
	.MonDReg_2(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_27(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_28(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_26(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.writedata_3(\writedata[3]~q ),
	.jdo_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.MonDReg_3(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_29(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ),
	.MonDReg_16(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_4(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.jdo_16(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ),
	.jdo_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.MonDReg_5(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ),
	.writedata_16(\writedata[16]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.jdo_8(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.writedata_4(\writedata[4]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_17(\writedata[17]~q ),
	.MonDReg_15(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_18(\writedata[18]~q ),
	.MonDReg_12(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.writedata_28(\writedata[28]~q ),
	.MonDReg_8(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_7(\writedata[7]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_31(\writedata[31]~q ),
	.MonDReg_11(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ),
	.writedata_11(\writedata[11]~q ),
	.MonDReg_9(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_22(\writedata[22]~q ),
	.MonDReg_14(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.writedata_30(\writedata[30]~q ),
	.jdo_9(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_15(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_11(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_13(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_10(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci_debug the_Qsys_system_nios2_qsys_0_nios2_oci_debug(
	.r_sync_rst(r_sync_rst),
	.jtag_break1(jtag_break),
	.monitor_ready1(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.jdo_35(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.jdo_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.resetrequest1(resetrequest),
	.jdo_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper|the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.resetlatch1(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ),
	.monitor_go1(\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!d_write),
	.datab(!saved_grant_0),
	.datac(!waitrequest),
	.datad(!mem_used_1),
	.datae(!WideOr1),
	.dataf(!\write~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFF3FFFFF7F7FFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!\read~q ),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \read~0 .shared_arith = "off";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~4_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclonev_lcell_comb \readdata~3 (
	.dataa(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal0~1_combout ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datac(!\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~3 .extended_lut = "off";
defparam \readdata~3 .lut_mask = 64'h2727272727272727;
defparam \readdata~3 .shared_arith = "off";

cyclonev_lcell_comb \readdata~4 (
	.dataa(!oci_single_step_mode),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal0~1_combout ),
	.datac(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~4 .extended_lut = "off";
defparam \readdata~4 .lut_mask = 64'h4747474747474747;
defparam \readdata~4 .shared_arith = "off";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!\address[8]~q ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \readdata[0]~1 (
	.dataa(!\address[8]~q ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_avalon_reg|Equal0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~1 .extended_lut = "off";
defparam \readdata[0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \readdata[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.datac(!oci_ienable_0),
	.datad(!\readdata[0]~0_combout ),
	.datae(!\readdata[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \readdata~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata~5 (
	.dataa(!\the_Qsys_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.datab(!\the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.datac(!oci_ienable_1),
	.datad(!\readdata[0]~0_combout ),
	.datae(!\readdata[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~5 .extended_lut = "off";
defparam \readdata~5 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \readdata~5 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_wrapper (
	break_readreg_0,
	break_readreg_1,
	MonDReg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_16,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	break_readreg_26,
	MonDReg_26,
	break_readreg_27,
	MonDReg_27,
	break_readreg_25,
	MonDReg_25,
	break_readreg_17,
	MonDReg_17,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	break_readreg_22,
	MonDReg_22,
	break_readreg_6,
	MonDReg_6,
	break_readreg_15,
	break_readreg_23,
	MonDReg_23,
	MonDReg_10,
	MonDReg_13,
	MonDReg_7,
	break_readreg_7,
	break_readreg_8,
	break_readreg_9,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	MonDReg_0,
	hbreak_enabled,
	monitor_ready,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_35,
	take_action_ocimem_a,
	take_action_ocimem_b,
	jdo_3,
	jdo_17,
	jdo_34,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_21,
	jdo_20,
	jdo_25,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_27,
	jdo_28,
	jdo_26,
	jdo_19,
	jdo_18,
	MonDReg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	MonDReg_16,
	monitor_error,
	MonDReg_4,
	jdo_6,
	jdo_16,
	jdo_23,
	jdo_22,
	MonDReg_18,
	jdo_24,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	resetlatch,
	jdo_8,
	MonDReg_15,
	MonDReg_12,
	MonDReg_8,
	MonDReg_11,
	MonDReg_9,
	MonDReg_14,
	jdo_9,
	jdo_15,
	jdo_11,
	jdo_13,
	jdo_10,
	jdo_14,
	jdo_12,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	break_readreg_1;
input 	MonDReg_1;
input 	break_readreg_2;
input 	break_readreg_3;
input 	break_readreg_16;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_22;
input 	MonDReg_22;
input 	break_readreg_6;
input 	MonDReg_6;
input 	break_readreg_15;
input 	break_readreg_23;
input 	MonDReg_23;
input 	MonDReg_10;
input 	MonDReg_13;
input 	MonDReg_7;
input 	break_readreg_7;
input 	break_readreg_8;
input 	break_readreg_9;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_13;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	MonDReg_0;
input 	hbreak_enabled;
input 	monitor_ready;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	jdo_35;
output 	take_action_ocimem_a;
output 	take_action_ocimem_b;
output 	jdo_3;
output 	jdo_17;
output 	jdo_34;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	jdo_21;
output 	jdo_20;
output 	jdo_25;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_27;
output 	jdo_28;
output 	jdo_26;
output 	jdo_19;
output 	jdo_18;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
input 	MonDReg_16;
input 	monitor_error;
input 	MonDReg_4;
output 	jdo_6;
output 	jdo_16;
output 	jdo_23;
output 	jdo_22;
input 	MonDReg_18;
output 	jdo_24;
input 	MonDReg_5;
output 	jdo_7;
input 	MonDReg_29;
input 	resetlatch;
output 	jdo_8;
input 	MonDReg_15;
input 	MonDReg_12;
input 	MonDReg_8;
input 	MonDReg_11;
input 	MonDReg_9;
input 	MonDReg_14;
output 	jdo_9;
output 	jdo_15;
output 	jdo_11;
output 	jdo_13;
output 	jdo_10;
output 	jdo_14;
output 	jdo_12;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ;
wire \Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ;
wire \Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ;
wire \Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ;
wire \Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ;
wire \the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ;


Qsys_system_sld_virtual_jtag_basic_1 Qsys_system_nios2_qsys_0_jtag_debug_module_phy(
	.virtual_state_sdr(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk the_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk(
	.sr_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ),
	.sr_3(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ),
	.sr_4(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ),
	.sr_17(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ),
	.sr_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ),
	.sr_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ),
	.sr_27(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ),
	.sr_28(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ),
	.sr_26(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ),
	.sr_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ),
	.sr_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ),
	.sr_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ),
	.sr_6(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ),
	.sr_29(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ),
	.sr_30(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ),
	.sr_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ),
	.sr_16(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ),
	.sr_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ),
	.sr_8(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ),
	.sr_9(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ),
	.sr_10(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ),
	.sr_11(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ),
	.sr_13(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ),
	.sr_14(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ),
	.sr_12(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_35(jdo_35),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.jdo_3(jdo_3),
	.jdo_17(jdo_17),
	.jdo_34(jdo_34),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ),
	.sr_35(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ),
	.jdo_27(jdo_27),
	.jdo_28(jdo_28),
	.jdo_26(jdo_26),
	.sr_34(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_6(jdo_6),
	.sr_31(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ),
	.jdo_16(jdo_16),
	.jdo_23(jdo_23),
	.jdo_22(jdo_22),
	.jdo_24(jdo_24),
	.sr_7(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.virtual_state_udr(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.jdo_8(jdo_8),
	.jdo_9(jdo_9),
	.jdo_15(jdo_15),
	.jdo_11(jdo_11),
	.jdo_13(jdo_13),
	.jdo_10(jdo_10),
	.jdo_14(jdo_14),
	.jdo_12(jdo_12),
	.sr_15(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_tck the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck(
	.sr_1(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.sr_3(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.sr_4(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.sr_17(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ),
	.sr_21(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ),
	.sr_25(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_27(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ),
	.sr_28(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ),
	.sr_26(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ),
	.sr_18(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.sr_22(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.sr_29(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ),
	.sr_30(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.sr_23(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.MonDReg_21(MonDReg_21),
	.break_readreg_18(break_readreg_18),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_29(break_readreg_29),
	.MonDReg_30(MonDReg_30),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.sr_16(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ),
	.sr_24(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.MonDReg_22(MonDReg_22),
	.sr_8(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.MonDReg_6(MonDReg_6),
	.break_readreg_15(break_readreg_15),
	.break_readreg_23(break_readreg_23),
	.MonDReg_23(MonDReg_23),
	.MonDReg_10(MonDReg_10),
	.MonDReg_13(MonDReg_13),
	.MonDReg_7(MonDReg_7),
	.sr_9(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ),
	.break_readreg_7(break_readreg_7),
	.sr_10(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ),
	.break_readreg_8(break_readreg_8),
	.sr_11(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ),
	.sr_13(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ),
	.sr_14(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ),
	.sr_12(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ),
	.break_readreg_9(break_readreg_9),
	.break_readreg_14(break_readreg_14),
	.break_readreg_10(break_readreg_10),
	.break_readreg_12(break_readreg_12),
	.break_readreg_13(break_readreg_13),
	.break_readreg_11(break_readreg_11),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.hbreak_enabled(hbreak_enabled),
	.monitor_ready(monitor_ready),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ),
	.sr_35(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ),
	.sr_34(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ),
	.MonDReg_3(MonDReg_3),
	.virtual_state_cdr(\Qsys_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.MonDReg_16(MonDReg_16),
	.monitor_error(monitor_error),
	.MonDReg_4(MonDReg_4),
	.sr_31(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ),
	.MonDReg_18(MonDReg_18),
	.sr_7(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ),
	.MonDReg_5(MonDReg_5),
	.MonDReg_29(MonDReg_29),
	.resetlatch(resetlatch),
	.MonDReg_15(MonDReg_15),
	.MonDReg_12(MonDReg_12),
	.MonDReg_8(MonDReg_8),
	.MonDReg_11(MonDReg_11),
	.MonDReg_9(MonDReg_9),
	.MonDReg_14(MonDReg_14),
	.sr_15(\the_Qsys_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_4,
	sr_17,
	sr_21,
	sr_20,
	sr_25,
	sr_5,
	sr_27,
	sr_28,
	sr_26,
	sr_18,
	sr_22,
	sr_19,
	sr_6,
	sr_29,
	sr_30,
	sr_32,
	sr_23,
	sr_16,
	sr_24,
	sr_8,
	sr_9,
	sr_10,
	sr_11,
	sr_13,
	sr_14,
	sr_12,
	sr_0,
	virtual_state_uir,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe1,
	jdo_35,
	take_action_ocimem_a1,
	take_action_ocimem_b1,
	jdo_3,
	jdo_17,
	jdo_34,
	take_action_ocimem_a2,
	take_action_ocimem_a3,
	jdo_21,
	jdo_20,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	sr_35,
	jdo_27,
	jdo_28,
	jdo_26,
	sr_34,
	jdo_19,
	jdo_18,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_6,
	sr_31,
	sr_33,
	jdo_16,
	jdo_23,
	jdo_22,
	jdo_24,
	sr_7,
	jdo_7,
	virtual_state_udr,
	jdo_8,
	jdo_9,
	jdo_15,
	jdo_11,
	jdo_13,
	jdo_10,
	jdo_14,
	jdo_12,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_4;
input 	sr_17;
input 	sr_21;
input 	sr_20;
input 	sr_25;
input 	sr_5;
input 	sr_27;
input 	sr_28;
input 	sr_26;
input 	sr_18;
input 	sr_22;
input 	sr_19;
input 	sr_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_23;
input 	sr_16;
input 	sr_24;
input 	sr_8;
input 	sr_9;
input 	sr_10;
input 	sr_11;
input 	sr_13;
input 	sr_14;
input 	sr_12;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	jdo_35;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_b1;
output 	jdo_3;
output 	jdo_17;
output 	jdo_34;
output 	take_action_ocimem_a2;
output 	take_action_ocimem_a3;
output 	jdo_21;
output 	jdo_20;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
input 	sr_35;
output 	jdo_27;
output 	jdo_28;
output 	jdo_26;
input 	sr_34;
output 	jdo_19;
output 	jdo_18;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
output 	jdo_16;
output 	jdo_23;
output 	jdo_22;
output 	jdo_24;
input 	sr_7;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_8;
output 	jdo_9;
output 	jdo_15;
output 	jdo_11;
output 	jdo_13;
output 	jdo_10;
output 	jdo_14;
output 	jdo_12;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


Qsys_system_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

Qsys_system_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_b(
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_b1),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_b.extended_lut = "off";
defparam take_action_ocimem_b.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_b.shared_arith = "off";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!take_action_ocimem_a2),
	.datab(!jdo_34),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module Qsys_system_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module Qsys_system_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_jtag_debug_module_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	sr_4,
	break_readreg_2,
	sr_17,
	sr_21,
	sr_20,
	sr_25,
	sr_5,
	break_readreg_3,
	sr_27,
	sr_28,
	sr_26,
	sr_18,
	break_readreg_16,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	sr_29,
	sr_30,
	sr_32,
	break_readreg_26,
	MonDReg_26,
	break_readreg_27,
	MonDReg_27,
	break_readreg_25,
	MonDReg_25,
	break_readreg_17,
	MonDReg_17,
	sr_23,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	sr_16,
	sr_24,
	break_readreg_22,
	MonDReg_22,
	sr_8,
	break_readreg_6,
	MonDReg_6,
	break_readreg_15,
	break_readreg_23,
	MonDReg_23,
	MonDReg_10,
	MonDReg_13,
	MonDReg_7,
	sr_9,
	break_readreg_7,
	sr_10,
	break_readreg_8,
	sr_11,
	sr_13,
	sr_14,
	sr_12,
	break_readreg_9,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	MonDReg_0,
	virtual_state_uir,
	hbreak_enabled,
	monitor_ready,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_35,
	sr_34,
	MonDReg_3,
	virtual_state_cdr,
	MonDReg_16,
	monitor_error,
	MonDReg_4,
	sr_31,
	sr_33,
	MonDReg_18,
	sr_7,
	MonDReg_5,
	MonDReg_29,
	resetlatch,
	MonDReg_15,
	MonDReg_12,
	MonDReg_8,
	MonDReg_11,
	MonDReg_9,
	MonDReg_14,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
output 	sr_4;
input 	break_readreg_2;
output 	sr_17;
output 	sr_21;
output 	sr_20;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
output 	sr_27;
output 	sr_28;
output 	sr_26;
output 	sr_18;
input 	break_readreg_16;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
output 	sr_29;
output 	sr_30;
output 	sr_32;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_17;
input 	MonDReg_17;
output 	sr_23;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
output 	sr_16;
output 	sr_24;
input 	break_readreg_22;
input 	MonDReg_22;
output 	sr_8;
input 	break_readreg_6;
input 	MonDReg_6;
input 	break_readreg_15;
input 	break_readreg_23;
input 	MonDReg_23;
input 	MonDReg_10;
input 	MonDReg_13;
input 	MonDReg_7;
output 	sr_9;
input 	break_readreg_7;
output 	sr_10;
input 	break_readreg_8;
output 	sr_11;
output 	sr_13;
output 	sr_14;
output 	sr_12;
input 	break_readreg_9;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_13;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	MonDReg_0;
input 	virtual_state_uir;
input 	hbreak_enabled;
input 	monitor_ready;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_35;
output 	sr_34;
input 	MonDReg_3;
input 	virtual_state_cdr;
input 	MonDReg_16;
input 	monitor_error;
input 	MonDReg_4;
output 	sr_31;
output 	sr_33;
input 	MonDReg_18;
output 	sr_7;
input 	MonDReg_5;
input 	MonDReg_29;
input 	resetlatch;
input 	MonDReg_15;
input 	MonDReg_12;
input 	MonDReg_8;
input 	MonDReg_11;
input 	MonDReg_9;
input 	MonDReg_14;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[5]~9_combout ;
wire \sr[5]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~13_combout ;
wire \sr~18_combout ;
wire \sr[24]~19_combout ;
wire \sr[24]~20_combout ;
wire \sr~22_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~39_combout ;
wire \sr~41_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \sr~14_combout ;
wire \sr[36]~15_combout ;
wire \sr~16_combout ;
wire \Mux37~0_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~17_combout ;
wire \sr~21_combout ;
wire \sr[24]~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~40_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr[24]~55_combout ;
wire \DRsize.010~q ;
wire \sr~49_combout ;
wire \sr~50_combout ;


Qsys_system_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

Qsys_system_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[24]~19_combout ),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[5]~9_combout ),
	.sload(gnd),
	.ena(\sr[5]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~15_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~15_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[24]~20_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[5]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[5]~9 .extended_lut = "off";
defparam \sr[5]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[5]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[5]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[5]~10 .extended_lut = "off";
defparam \sr[5]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~13 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr[24]~19 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[24]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[24]~19 .extended_lut = "off";
defparam \sr[24]~19 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[24]~19 .shared_arith = "off";

cyclonev_lcell_comb \sr[24]~20 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[24]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[24]~20 .extended_lut = "off";
defparam \sr[24]~20 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[24]~20 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_19),
	.datad(!break_readreg_17),
	.datae(!MonDReg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_23),
	.datad(!break_readreg_21),
	.datae(!MonDReg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_20),
	.datad(!break_readreg_18),
	.datae(!MonDReg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~32 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_7),
	.datad(!break_readreg_5),
	.datae(!MonDReg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~32 .extended_lut = "off";
defparam \sr~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~33 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_30),
	.datad(!break_readreg_28),
	.datae(!MonDReg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~33 .extended_lut = "off";
defparam \sr~33 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_31),
	.datad(!break_readreg_29),
	.datae(!MonDReg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_33),
	.datad(!break_readreg_31),
	.datae(!MonDReg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_24),
	.datad(!break_readreg_22),
	.datae(!MonDReg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_17),
	.datad(!break_readreg_15),
	.datae(!MonDReg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_25),
	.datad(!break_readreg_23),
	.datae(!MonDReg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_7),
	.datad(!sr_9),
	.datae(!break_readreg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~51 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~54 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \sr~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~14 .extended_lut = "off";
defparam \sr~14 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~14 .shared_arith = "off";

cyclonev_lcell_comb \sr[36]~15 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[36]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[36]~15 .extended_lut = "off";
defparam \sr[36]~15 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[36]~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_2),
	.datad(!irf_reg_1_2),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~17 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~17 .extended_lut = "off";
defparam \sr~17 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~17 .shared_arith = "off";

cyclonev_lcell_comb \sr~21 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~21 .extended_lut = "off";
defparam \sr~21 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~21 .shared_arith = "off";

cyclonev_lcell_comb \sr[24]~35 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[24]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[24]~35 .extended_lut = "off";
defparam \sr[24]~35 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[24]~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~36 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~36 .extended_lut = "off";
defparam \sr~36 .lut_mask = 64'h2727272727272727;
defparam \sr~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[24]~35_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~36_combout ),
	.dataf(!\sr~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!irf_reg_1_2),
	.datab(!break_readreg_6),
	.datac(!MonDReg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'h2727272727272727;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_2),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~42_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr[24]~55 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[24]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[24]~55 .extended_lut = "off";
defparam \sr[24]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[24]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[24]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_2),
	.datac(!irf_reg_1_2),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~49 .shared_arith = "off";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~50 .shared_arith = "off";

endmodule

module Qsys_system_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module Qsys_system_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module Qsys_system_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	oci_single_step_mode1,
	writedata_0,
	address_0,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	debugaccess,
	take_action_ocireg,
	writedata_3,
	writedata_1,
	oci_ienable_0,
	oci_ienable_1,
	Equal1,
	oci_reg_readdata,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
output 	oci_single_step_mode1;
input 	writedata_0;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
output 	Equal0;
input 	debugaccess;
output 	take_action_ocireg;
input 	writedata_3;
input 	writedata_1;
output 	oci_ienable_0;
output 	oci_ienable_1;
output 	Equal1;
output 	oci_reg_readdata;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_single_step_mode~0_combout ;
wire \Equal0~0_combout ;
wire \oci_ienable[0]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[1]~1_combout ;
wire \oci_ienable[31]~q ;


dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!write),
	.datab(!Equal0),
	.datac(!debugaccess),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(\oci_ienable[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas \oci_ienable[1] (
	.clk(clk_clk),
	.d(\oci_ienable[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_reg_readdata~0 (
	.dataa(!Equal1),
	.datab(!\oci_ienable[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~0 .extended_lut = "off";
defparam \oci_reg_readdata~0 .lut_mask = 64'h7777777777777777;
defparam \oci_reg_readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!oci_single_step_mode1),
	.datab(!take_action_ocireg),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h4747474747474747;
defparam \oci_single_step_mode~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(!address_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[0]~0 (
	.dataa(!writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[0]~0 .extended_lut = "off";
defparam \oci_ienable[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(!write),
	.datab(!debugaccess),
	.datac(!Equal1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_oci_intr_mask_reg~0 .extended_lut = "off";
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_oci_intr_mask_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[1]~1 (
	.dataa(!writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[1]~1 .extended_lut = "off";
defparam \oci_ienable[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[1]~1 .shared_arith = "off";

dffeas \oci_ienable[31] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(\oci_ienable[31]~q ),
	.prn(vcc));
defparam \oci_ienable[31] .is_wysiwyg = "true";
defparam \oci_ienable[31] .power_up = "low";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_16,
	break_readreg_20,
	break_readreg_19,
	break_readreg_24,
	break_readreg_4,
	break_readreg_26,
	break_readreg_27,
	break_readreg_25,
	break_readreg_17,
	break_readreg_21,
	break_readreg_18,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_22,
	break_readreg_6,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_8,
	break_readreg_9,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_3,
	jdo_17,
	jdo_21,
	jdo_20,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_27,
	jdo_28,
	jdo_26,
	jdo_19,
	jdo_18,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_6,
	jdo_16,
	jdo_23,
	jdo_22,
	jdo_24,
	jdo_7,
	jdo_8,
	jdo_9,
	jdo_15,
	jdo_11,
	jdo_13,
	jdo_10,
	jdo_14,
	jdo_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_3;
output 	break_readreg_16;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_26;
output 	break_readreg_27;
output 	break_readreg_25;
output 	break_readreg_17;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_5;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_22;
output 	break_readreg_6;
output 	break_readreg_15;
output 	break_readreg_23;
output 	break_readreg_7;
output 	break_readreg_8;
output 	break_readreg_9;
output 	break_readreg_14;
output 	break_readreg_10;
output 	break_readreg_12;
output 	break_readreg_13;
output 	break_readreg_11;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_27;
input 	jdo_28;
input 	jdo_26;
input 	jdo_19;
input 	jdo_18;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_6;
input 	jdo_16;
input 	jdo_23;
input 	jdo_22;
input 	jdo_24;
input 	jdo_7;
input 	jdo_8;
input 	jdo_9;
input 	jdo_15;
input 	jdo_11;
input 	jdo_13;
input 	jdo_10;
input 	jdo_14;
input 	jdo_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[10]~0_combout ;
wire \break_readreg[10]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[10]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[10]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

cyclonev_lcell_comb \break_readreg[10]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[10]~0 .extended_lut = "off";
defparam \break_readreg[10]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[10]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[10]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[10]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[10]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[10]~1 .extended_lut = "off";
defparam \break_readreg[10]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[10]~1 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_nios2_oci_debug (
	r_sync_rst,
	jtag_break1,
	monitor_ready1,
	jdo_35,
	take_action_ocimem_a,
	jdo_34,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	jdo_25,
	writedata_0,
	take_action_ocireg,
	jdo_19,
	jdo_18,
	writedata_1,
	monitor_error1,
	jdo_23,
	jdo_22,
	resetrequest1,
	jdo_24,
	resetlatch1,
	monitor_go1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	jtag_break1;
output 	monitor_ready1;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
input 	jdo_25;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_19;
input 	jdo_18;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_23;
input 	jdo_22;
output 	resetrequest1;
input 	jdo_24;
output 	resetlatch1;
output 	monitor_go1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \resetlatch~0_combout ;
wire \monitor_go~0_combout ;


Qsys_system_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas resetrequest(
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(resetrequest1),
	.prn(vcc));
defparam resetrequest.is_wysiwyg = "true";
defparam resetrequest.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!\break_on_reset~q ),
	.datab(!jdo_19),
	.datac(!jdo_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!monitor_ready1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_25),
	.datad(!writedata_0),
	.datae(!take_action_ocireg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_25),
	.datac(!take_action_ocireg),
	.datad(!writedata_1),
	.datae(!monitor_error1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(!jdo_34),
	.datad(!jdo_23),
	.datae(!monitor_go1),
	.dataf(!state_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \monitor_go~0 .shared_arith = "off";

endmodule

module Qsys_system_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_nios2_ocimem (
	MonDReg_1,
	q_a_0,
	q_a_1,
	q_a_2,
	MonDReg_20,
	MonDReg_19,
	MonDReg_24,
	q_a_3,
	MonDReg_26,
	MonDReg_27,
	MonDReg_25,
	MonDReg_17,
	q_a_16,
	MonDReg_21,
	q_a_20,
	q_a_19,
	q_a_24,
	q_a_4,
	MonDReg_28,
	MonDReg_30,
	MonDReg_31,
	q_a_26,
	q_a_27,
	q_a_25,
	q_a_17,
	MonDReg_22,
	q_a_21,
	q_a_18,
	q_a_12,
	q_a_28,
	q_a_8,
	q_a_10,
	q_a_5,
	q_a_13,
	q_a_29,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_9,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	MonDReg_6,
	MonDReg_23,
	MonDReg_10,
	MonDReg_13,
	MonDReg_7,
	waitrequest1,
	MonDReg_0,
	write,
	address_8,
	read,
	jdo_35,
	take_action_ocimem_a,
	take_action_ocimem_b,
	jdo_3,
	jdo_17,
	jdo_34,
	take_no_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	jdo_25,
	writedata_0,
	address_0,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	debugaccess,
	MonDReg_2,
	jdo_4,
	r_early_rst,
	byteenable_0,
	jdo_27,
	jdo_28,
	jdo_26,
	writedata_3,
	jdo_19,
	jdo_18,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	MonDReg_16,
	MonDReg_4,
	jdo_6,
	writedata_2,
	jdo_16,
	jdo_23,
	jdo_22,
	MonDReg_18,
	jdo_24,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	writedata_16,
	byteenable_2,
	writedata_20,
	writedata_19,
	writedata_24,
	byteenable_3,
	jdo_8,
	writedata_4,
	writedata_26,
	writedata_27,
	writedata_25,
	writedata_17,
	MonDReg_15,
	writedata_21,
	writedata_18,
	MonDReg_12,
	writedata_12,
	byteenable_1,
	writedata_28,
	MonDReg_8,
	writedata_8,
	writedata_10,
	writedata_5,
	writedata_13,
	writedata_29,
	writedata_7,
	writedata_23,
	writedata_15,
	writedata_31,
	MonDReg_11,
	writedata_11,
	MonDReg_9,
	writedata_9,
	writedata_6,
	writedata_22,
	MonDReg_14,
	writedata_14,
	writedata_30,
	jdo_9,
	jdo_15,
	jdo_11,
	jdo_13,
	jdo_10,
	jdo_14,
	jdo_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_24;
output 	q_a_3;
output 	MonDReg_26;
output 	MonDReg_27;
output 	MonDReg_25;
output 	MonDReg_17;
output 	q_a_16;
output 	MonDReg_21;
output 	q_a_20;
output 	q_a_19;
output 	q_a_24;
output 	q_a_4;
output 	MonDReg_28;
output 	MonDReg_30;
output 	MonDReg_31;
output 	q_a_26;
output 	q_a_27;
output 	q_a_25;
output 	q_a_17;
output 	MonDReg_22;
output 	q_a_21;
output 	q_a_18;
output 	q_a_12;
output 	q_a_28;
output 	q_a_8;
output 	q_a_10;
output 	q_a_5;
output 	q_a_13;
output 	q_a_29;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_9;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	MonDReg_6;
output 	MonDReg_23;
output 	MonDReg_10;
output 	MonDReg_13;
output 	MonDReg_7;
output 	waitrequest1;
output 	MonDReg_0;
input 	write;
input 	address_8;
input 	read;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	take_action_ocimem_b;
input 	jdo_3;
input 	jdo_17;
input 	jdo_34;
input 	take_no_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
input 	jdo_25;
input 	writedata_0;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	debugaccess;
output 	MonDReg_2;
input 	jdo_4;
input 	r_early_rst;
input 	byteenable_0;
input 	jdo_27;
input 	jdo_28;
input 	jdo_26;
input 	writedata_3;
input 	jdo_19;
input 	jdo_18;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
output 	MonDReg_16;
output 	MonDReg_4;
input 	jdo_6;
input 	writedata_2;
input 	jdo_16;
input 	jdo_23;
input 	jdo_22;
output 	MonDReg_18;
input 	jdo_24;
output 	MonDReg_5;
input 	jdo_7;
output 	MonDReg_29;
input 	writedata_16;
input 	byteenable_2;
input 	writedata_20;
input 	writedata_19;
input 	writedata_24;
input 	byteenable_3;
input 	jdo_8;
input 	writedata_4;
input 	writedata_26;
input 	writedata_27;
input 	writedata_25;
input 	writedata_17;
output 	MonDReg_15;
input 	writedata_21;
input 	writedata_18;
output 	MonDReg_12;
input 	writedata_12;
input 	byteenable_1;
input 	writedata_28;
output 	MonDReg_8;
input 	writedata_8;
input 	writedata_10;
input 	writedata_5;
input 	writedata_13;
input 	writedata_29;
input 	writedata_7;
input 	writedata_23;
input 	writedata_15;
input 	writedata_31;
output 	MonDReg_11;
input 	writedata_11;
output 	MonDReg_9;
input 	writedata_9;
input 	writedata_6;
input 	writedata_22;
output 	MonDReg_14;
input 	writedata_14;
input 	writedata_30;
input 	jdo_9;
input 	jdo_15;
input 	jdo_11;
input 	jdo_13;
input 	jdo_10;
input 	jdo_14;
input 	jdo_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[3]~3_combout ;
wire \ociram_wr_data[16]~4_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[20]~5_combout ;
wire \ociram_wr_data[19]~6_combout ;
wire \ociram_wr_data[24]~7_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[4]~8_combout ;
wire \ociram_wr_data[26]~9_combout ;
wire \ociram_wr_data[27]~10_combout ;
wire \ociram_wr_data[25]~11_combout ;
wire \ociram_wr_data[17]~12_combout ;
wire \ociram_wr_data[21]~13_combout ;
wire \ociram_wr_data[18]~14_combout ;
wire \ociram_wr_data[12]~15_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[28]~16_combout ;
wire \ociram_wr_data[8]~17_combout ;
wire \ociram_wr_data[10]~18_combout ;
wire \ociram_wr_data[5]~19_combout ;
wire \ociram_wr_data[13]~20_combout ;
wire \ociram_wr_data[29]~21_combout ;
wire \ociram_wr_data[7]~22_combout ;
wire \ociram_wr_data[23]~23_combout ;
wire \ociram_wr_data[15]~24_combout ;
wire \ociram_wr_data[31]~25_combout ;
wire \ociram_wr_data[11]~26_combout ;
wire \ociram_wr_data[9]~27_combout ;
wire \ociram_wr_data[6]~28_combout ;
wire \ociram_wr_data[22]~29_combout ;
wire \ociram_wr_data[14]~30_combout ;
wire \ociram_wr_data[30]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~13_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~14 ;
wire \Add0~5_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~10 ;
wire \Add0~21_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~34 ;
wire \Add0~17_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[6]~3_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~2_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~0_combout ;
wire \MonDReg~1_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg~7_combout ;
wire \MonDReg~8_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~11_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;


Qsys_system_Qsys_system_nios2_qsys_0_ociram_sp_ram_module Qsys_system_nios2_qsys_0_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_16(q_a_16),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_24(q_a_24),
	.q_a_4(q_a_4),
	.q_a_26(q_a_26),
	.q_a_27(q_a_27),
	.q_a_25(q_a_25),
	.q_a_17(q_a_17),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.q_a_12(q_a_12),
	.q_a_28(q_a_28),
	.q_a_8(q_a_8),
	.q_a_10(q_a_10),
	.q_a_5(q_a_5),
	.q_a_13(q_a_13),
	.q_a_29(q_a_29),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_11(q_a_11),
	.q_a_9(q_a_9),
	.q_a_6(q_a_6),
	.q_a_22(q_a_22),
	.q_a_14(q_a_14),
	.q_a_30(q_a_30),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~3_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~4_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~5_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~6_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~7_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~8_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~9_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~10_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~11_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~12_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~13_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~14_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~15_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~16_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~17_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~18_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~19_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~20_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~21_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~22_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~23_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~24_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~25_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~26_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~27_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~28_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~29_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~30_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!write),
	.datab(!address_8),
	.datac(!\jtag_ram_access~q ),
	.datad(!debugaccess),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!address_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[5]~q ),
	.datac(!address_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[6]~q ),
	.datac(!address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[7]~q ),
	.datac(!address_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[8]~q ),
	.datac(!address_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[9]~q ),
	.datac(!address_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_1),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!take_action_ocimem_b),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'h7777777777777777;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!writedata_3),
	.datac(!MonDReg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~3 .extended_lut = "off";
defparam \ociram_wr_data[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_16),
	.datac(!writedata_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~4 .extended_lut = "off";
defparam \ociram_wr_data[16]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~1 .extended_lut = "off";
defparam \ociram_byteenable[2]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~5 .extended_lut = "off";
defparam \ociram_wr_data[20]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~6 .extended_lut = "off";
defparam \ociram_wr_data[19]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~7 .extended_lut = "off";
defparam \ociram_wr_data[24]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~2 .extended_lut = "off";
defparam \ociram_byteenable[3]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~8 .extended_lut = "off";
defparam \ociram_wr_data[4]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~9 .extended_lut = "off";
defparam \ociram_wr_data[26]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~10 .extended_lut = "off";
defparam \ociram_wr_data[27]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~11 .extended_lut = "off";
defparam \ociram_wr_data[25]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~12 .extended_lut = "off";
defparam \ociram_wr_data[17]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~13 .extended_lut = "off";
defparam \ociram_wr_data[21]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~14 .extended_lut = "off";
defparam \ociram_wr_data[18]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~15 .extended_lut = "off";
defparam \ociram_wr_data[12]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~3 .extended_lut = "off";
defparam \ociram_byteenable[1]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~16 .extended_lut = "off";
defparam \ociram_wr_data[28]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~17 .extended_lut = "off";
defparam \ociram_wr_data[8]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~18 .extended_lut = "off";
defparam \ociram_wr_data[10]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~19 .extended_lut = "off";
defparam \ociram_wr_data[5]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~20 .extended_lut = "off";
defparam \ociram_wr_data[13]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~21 .extended_lut = "off";
defparam \ociram_wr_data[29]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~22 .extended_lut = "off";
defparam \ociram_wr_data[7]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~23 .extended_lut = "off";
defparam \ociram_wr_data[23]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~24 .extended_lut = "off";
defparam \ociram_wr_data[15]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~25 .extended_lut = "off";
defparam \ociram_wr_data[31]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~26 .extended_lut = "off";
defparam \ociram_wr_data[11]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~27 .extended_lut = "off";
defparam \ociram_wr_data[9]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~28 .extended_lut = "off";
defparam \ociram_wr_data[6]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~29 .extended_lut = "off";
defparam \ociram_wr_data[22]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~30 .extended_lut = "off";
defparam \ociram_wr_data[14]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~31 .extended_lut = "off";
defparam \ociram_wr_data[30]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~31 .shared_arith = "off";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(q_a_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(q_a_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(q_a_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(q_a_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[6]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(\MonDReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!take_no_action_ocimem_a),
	.datab(!jdo_17),
	.datac(!jdo_34),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[6]~3 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[6]~3 .extended_lut = "off";
defparam \MonDReg[6]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg[6]~3 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_no_action_ocimem_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~2 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~2 .extended_lut = "off";
defparam \MonDReg[0]~2 .lut_mask = 64'h4747474747474747;
defparam \MonDReg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(!jdo_17),
	.datad(!jdo_34),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hF7FBFFFFF7FBFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~0 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~0 .extended_lut = "off";
defparam \MonDReg~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \MonDReg~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~1 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_3),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!q_a_0),
	.datae(!\MonDReg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~1 .extended_lut = "off";
defparam \MonDReg~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!jdo_5),
	.datad(!\MonDReg~4_combout ),
	.datae(!q_a_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~6 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~4_combout ),
	.datad(!jdo_6),
	.datae(!q_a_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~6 .extended_lut = "off";
defparam \MonDReg~6 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~7 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~7 .extended_lut = "off";
defparam \MonDReg~7 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \MonDReg~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~8 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!jdo_19),
	.datad(!q_a_16),
	.datae(!\MonDReg~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~8 .extended_lut = "off";
defparam \MonDReg~8 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~8 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~9 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!jdo_7),
	.datae(!q_a_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~9 .extended_lut = "off";
defparam \MonDReg~9 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~9 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~20 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!q_a_18),
	.datad(!jdo_21),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~20 .extended_lut = "on";
defparam \MonDReg~20 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \MonDReg~20 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~10 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~10 .extended_lut = "off";
defparam \MonDReg~10 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \MonDReg~10 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~11 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!q_a_5),
	.datad(!jdo_8),
	.datae(!\MonDReg~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~11 .extended_lut = "off";
defparam \MonDReg~11 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~11 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~12 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~4_combout ),
	.datad(!jdo_32),
	.datae(!q_a_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~12 .extended_lut = "off";
defparam \MonDReg~12 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~12 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~13 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!jdo_18),
	.datad(!q_a_15),
	.datae(!\MonDReg~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~13 .extended_lut = "off";
defparam \MonDReg~13 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~13 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~14 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_12),
	.datae(!jdo_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~14 .extended_lut = "off";
defparam \MonDReg~14 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~14 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~15 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(!q_a_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~15 .extended_lut = "off";
defparam \MonDReg~15 .lut_mask = 64'hEDDEFFFFEDDEFFFF;
defparam \MonDReg~15 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~16 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_rd_d1~q ),
	.datac(!MonDReg_8),
	.datad(!jdo_11),
	.datae(!\MonDReg~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~16 .extended_lut = "off";
defparam \MonDReg~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~16 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~17 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~4_combout ),
	.datad(!q_a_11),
	.datae(!jdo_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~17 .extended_lut = "off";
defparam \MonDReg~17 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~17 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~18 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~4_combout ),
	.datad(!q_a_9),
	.datae(!jdo_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~18 .extended_lut = "off";
defparam \MonDReg~18 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~18 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~19 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!jdo_17),
	.datad(!\MonDReg~7_combout ),
	.datae(!q_a_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~19 .extended_lut = "off";
defparam \MonDReg~19 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~19 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_16,
	q_a_20,
	q_a_19,
	q_a_24,
	q_a_4,
	q_a_26,
	q_a_27,
	q_a_25,
	q_a_17,
	q_a_21,
	q_a_18,
	q_a_12,
	q_a_28,
	q_a_8,
	q_a_10,
	q_a_5,
	q_a_13,
	q_a_29,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_9,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_3,
	ociram_wr_data_16,
	ociram_byteenable_2,
	ociram_wr_data_20,
	ociram_wr_data_19,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_4,
	ociram_wr_data_26,
	ociram_wr_data_27,
	ociram_wr_data_25,
	ociram_wr_data_17,
	ociram_wr_data_21,
	ociram_wr_data_18,
	ociram_wr_data_12,
	ociram_byteenable_1,
	ociram_wr_data_28,
	ociram_wr_data_8,
	ociram_wr_data_10,
	ociram_wr_data_5,
	ociram_wr_data_13,
	ociram_wr_data_29,
	ociram_wr_data_7,
	ociram_wr_data_23,
	ociram_wr_data_15,
	ociram_wr_data_31,
	ociram_wr_data_11,
	ociram_wr_data_9,
	ociram_wr_data_6,
	ociram_wr_data_22,
	ociram_wr_data_14,
	ociram_wr_data_30,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_16;
output 	q_a_20;
output 	q_a_19;
output 	q_a_24;
output 	q_a_4;
output 	q_a_26;
output 	q_a_27;
output 	q_a_25;
output 	q_a_17;
output 	q_a_21;
output 	q_a_18;
output 	q_a_12;
output 	q_a_28;
output 	q_a_8;
output 	q_a_10;
output 	q_a_5;
output 	q_a_13;
output 	q_a_29;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_9;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_3;
input 	ociram_wr_data_16;
input 	ociram_byteenable_2;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_26;
input 	ociram_wr_data_27;
input 	ociram_wr_data_25;
input 	ociram_wr_data_17;
input 	ociram_wr_data_21;
input 	ociram_wr_data_18;
input 	ociram_wr_data_12;
input 	ociram_byteenable_1;
input 	ociram_wr_data_28;
input 	ociram_wr_data_8;
input 	ociram_wr_data_10;
input 	ociram_wr_data_5;
input 	ociram_wr_data_13;
input 	ociram_wr_data_29;
input 	ociram_wr_data_7;
input 	ociram_wr_data_23;
input 	ociram_wr_data_15;
input 	ociram_wr_data_31;
input 	ociram_wr_data_11;
input 	ociram_wr_data_9;
input 	ociram_wr_data_6;
input 	ociram_wr_data_22;
input 	ociram_wr_data_14;
input 	ociram_wr_data_30;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_7 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_7 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_psf1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_psf1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "D2622080506BCF0D06D1F082E980277062912CB244CFD084FC8EC49C6B4F28A5";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "8B4466F9986418FBBDC2D79799D62A2EBCDE87554821870A4291446385CAE645";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "9291633A992C2A4C071E706E6722D5D1FDC707F573CF0D406D54B651FC97C911";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "E6414F950EEE46E51336E633C4C82AD564200DDC93F4E4FCFE0F10D3E8843064";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "7B21D3BF8815D6EA52ACA5D90182D0FEE54279153DC162279DA35E59C350C65A";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "CB2A4C0DBABA3E5B0DC65CF4DC015DC4B93CAC73E3F541C878BD0279B1FC525F";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "9A078BB0528D733F0CE7360DDF4DBED01AA957F9DF48CA69E672F9EEDAFEAC73";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "A3591611CFF2626AB6D5471DD74C4854A7C640358F5D02EF6605C204E43D4148";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "FA490C89DA0AC7212C6B79E89849B2238B9BB6E73FE43D9BC8C166A1F9C0F6BA";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "3BC6737C19A08111F0CD2B4C4C58C3FB8AF5BED936D1221A104CAA70AAD52763";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "D61C0B3AE958620CF874FB552A1D483607D3E50925BCD213C99CC386063369FA";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "0AA96047012728D997AD87894BF09AAB5618DC7D301FAFF1AB6CCC1AFF1791A2";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "935D90F92BF4047F2973C1F7B73EE93A06E9824DC9DAEC9FDFADDB2ACDCFC8DE";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "932DB0CD28E8539066BFB50B0604E542D1D67047F6548C867D78F987A48D04D1";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "1B469EDD4BC3F1041988DEF2B79C2B0A6D738AD7EB2EFDC138C31CA5C1478DB6";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "8E1C13F7E86ED8B5C2E0CAFE8146F9752B2065A8CED2B02561410CA1B76131DB";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "F76FD2FACB3874CB7F69A2230993CF91AB682BECD42F86F58035612579521761";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "C9E45E8E2CCA3F98B355B4D77C1E3C88B38DC941C69776E33B1C652A6C84E883";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "43A4ABBA72442BE0093687C0D5782816FE7CE5847E0EC072EE77BF6263BECDFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "575EB9B1E2FF67F9B8C056385C7763CD70C3C6A16547526E3BE75D897A6DE98A";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "81688105F14E5EEC9F1AD891C645AC0EC442B741340091FA518E10D334A5CC00";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "AEE59F4ED31DC21880DB480F616A1CF268494538501BEFD54167C5679AB69793";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "AFF69E4C1F6675D4244D809042A238CD1915199CC77B204E9890128E2108FD03";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "430E04BE6ABADBE8C2C2F2FF32884A75FB4E414BCC5ED0D90F02E051607E4586";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "C81F56BE0FCB022E30A1E454C43F0A08EDEA0EE78B116A19AFE6DB876AD24EC2";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "6C196508DD5113A38E018C39BEA8FC3C6D2B053FC6729A29ACA3A834D004F110";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "8871A8A81B1AAAD3D7D688E515FCA96491A7760B8047458582F91DAF2659A83C";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "C97E62A2C8A25E376C028612C41166A7972AFBFFC4A72AA1DEC34D8048511E87";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "5696F0BA9F8E9501E35ED88C8AC651B0172375610EAA646E019096C91D55B564";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "89205FF25143060CBCF9A3D3B17971E078A0354875B91E2AA9D03DE4032006CE";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "B789C6A4915740F2841D3E15CCDE46521E7FCEBD107E14CF06B37D5ED68D563B";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "Qsys_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_nios2_oci:the_Qsys_system_nios2_qsys_0_nios2_oci|Qsys_system_nios2_qsys_0_nios2_ocimem:the_Qsys_system_nios2_qsys_0_nios2_ocimem|Qsys_system_nios2_qsys_0_ociram_sp_ram_module:Qsys_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_psf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "39B5F5641D6C8836BF000D1DCE468A1830B27E519D02FAF7E48644C58296B6B8";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_register_bank_a_module (
	q_b_4,
	q_b_2,
	q_b_5,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_3,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_30,
	q_b_26,
	q_b_25,
	q_b_0,
	q_b_19,
	q_b_1,
	q_b_17,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_18,
	q_b_24,
	q_b_23,
	q_b_31,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_14,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_29,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_31,
	A_dst_regnum_from_M_4,
	A_wr_dst_reg_from_M,
	A_dst_regnum_from_M_0,
	A_dst_regnum_from_M_1,
	A_dst_regnum_from_M_2,
	A_dst_regnum_from_M_3,
	rf_a_rd_port_addr_0,
	rf_a_rd_port_addr_1,
	rf_a_rd_port_addr_2,
	rf_a_rd_port_addr_3,
	rf_a_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_2;
output 	q_b_5;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_3;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_30;
output 	q_b_26;
output 	q_b_25;
output 	q_b_0;
output 	q_b_19;
output 	q_b_1;
output 	q_b_17;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_18;
output 	q_b_24;
output 	q_b_23;
output 	q_b_31;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_14;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_29;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_31;
input 	A_dst_regnum_from_M_4;
input 	A_wr_dst_reg_from_M;
input 	A_dst_regnum_from_M_0;
input 	A_dst_regnum_from_M_1;
input 	A_dst_regnum_from_M_2;
input 	A_dst_regnum_from_M_3;
input 	rf_a_rd_port_addr_0;
input 	rf_a_rd_port_addr_1;
input 	rf_a_rd_port_addr_2;
input 	rf_a_rd_port_addr_3;
input 	rf_a_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_8 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dst_regnum_from_M_4,A_dst_regnum_from_M_3,A_dst_regnum_from_M_2,A_dst_regnum_from_M_1,A_dst_regnum_from_M_0}),
	.wren_a(A_wr_dst_reg_from_M),
	.address_b({gnd,gnd,gnd,gnd,gnd,rf_a_rd_port_addr_4,rf_a_rd_port_addr_3,rf_a_rd_port_addr_2,rf_a_rd_port_addr_1,rf_a_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_8 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	wren_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_fin1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_fin1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "Qsys_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_a_module:Qsys_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_fin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

endmodule

module Qsys_system_Qsys_system_nios2_qsys_0_register_bank_b_module (
	q_b_4,
	q_b_0,
	q_b_2,
	q_b_5,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_3,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_30,
	q_b_26,
	q_b_25,
	q_b_19,
	q_b_1,
	q_b_17,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_18,
	q_b_24,
	q_b_23,
	q_b_31,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_14,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_29,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_31,
	A_dst_regnum_from_M_4,
	A_wr_dst_reg_from_M,
	A_dst_regnum_from_M_0,
	A_dst_regnum_from_M_1,
	A_dst_regnum_from_M_2,
	A_dst_regnum_from_M_3,
	rf_b_rd_port_addr_0,
	rf_b_rd_port_addr_1,
	rf_b_rd_port_addr_2,
	rf_b_rd_port_addr_3,
	rf_b_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_0;
output 	q_b_2;
output 	q_b_5;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_3;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_30;
output 	q_b_26;
output 	q_b_25;
output 	q_b_19;
output 	q_b_1;
output 	q_b_17;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_18;
output 	q_b_24;
output 	q_b_23;
output 	q_b_31;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_14;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_29;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_31;
input 	A_dst_regnum_from_M_4;
input 	A_wr_dst_reg_from_M;
input 	A_dst_regnum_from_M_0;
input 	A_dst_regnum_from_M_1;
input 	A_dst_regnum_from_M_2;
input 	A_dst_regnum_from_M_3;
input 	rf_b_rd_port_addr_0;
input 	rf_b_rd_port_addr_1;
input 	rf_b_rd_port_addr_2;
input 	rf_b_rd_port_addr_3;
input 	rf_b_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_9 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dst_regnum_from_M_4,A_dst_regnum_from_M_3,A_dst_regnum_from_M_2,A_dst_regnum_from_M_1,A_dst_regnum_from_M_0}),
	.wren_a(A_wr_dst_reg_from_M),
	.address_b({gnd,gnd,gnd,gnd,gnd,rf_b_rd_port_addr_4,rf_b_rd_port_addr_3,rf_b_rd_port_addr_2,rf_b_rd_port_addr_1,rf_b_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module Qsys_system_altsyncram_9 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	wren_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_gin1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_gin1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "Qsys_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "Qsys_system_nios2_qsys_0:nios2_qsys_0|Qsys_system_nios2_qsys_0_register_bank_b_module:Qsys_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_gin1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

endmodule

module Qsys_system_Qsys_system_onchip_ram (
	q_a_4,
	q_a_20,
	q_a_12,
	q_a_28,
	q_a_0,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_2,
	q_a_18,
	q_a_10,
	q_a_26,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_9,
	q_a_25,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	d_write,
	saved_grant_0,
	mem_used_1,
	src1_valid,
	src3_valid,
	saved_grant_1,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_data_33,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_4;
output 	q_a_20;
output 	q_a_12;
output 	q_a_28;
output 	q_a_0;
output 	q_a_16;
output 	q_a_8;
output 	q_a_24;
output 	q_a_2;
output 	q_a_18;
output 	q_a_10;
output 	q_a_26;
output 	q_a_5;
output 	q_a_21;
output 	q_a_13;
output 	q_a_29;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_27;
output 	q_a_9;
output 	q_a_25;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	q_a_3;
output 	q_a_19;
output 	q_a_1;
output 	q_a_17;
input 	d_write;
input 	saved_grant_0;
input 	mem_used_1;
input 	src1_valid;
input 	src3_valid;
input 	saved_grant_1;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_data_33;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


Qsys_system_altsyncram_10 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload19,src_payload27,src_payload15,src_payload3,src_payload21,src_payload11,src_payload23,src_payload7,src_payload17,src_payload25,src_payload13,src_payload1,src_payload29,src_payload9,src_payload31,src_payload5,src_payload18,src_payload26,src_payload14,src_payload2,
src_payload20,src_payload10,src_payload22,src_payload6,src_payload16,src_payload24,src_payload12,src_payload,src_payload28,src_payload8,src_payload30,src_payload4}),
	.address_a({src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!src1_valid),
	.datae(!src3_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \wren~0 .shared_arith = "off";

endmodule

module Qsys_system_altsyncram_10 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_l9n1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_l9n1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 5119;
defparam ram_block1a4.port_a_logical_ram_depth = 5120;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 5119;
defparam ram_block1a20.port_a_logical_ram_depth = 5120;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 5119;
defparam ram_block1a12.port_a_logical_ram_depth = 5120;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 5119;
defparam ram_block1a28.port_a_logical_ram_depth = 5120;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 5119;
defparam ram_block1a0.port_a_logical_ram_depth = 5120;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 5119;
defparam ram_block1a16.port_a_logical_ram_depth = 5120;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 5119;
defparam ram_block1a8.port_a_logical_ram_depth = 5120;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 5119;
defparam ram_block1a24.port_a_logical_ram_depth = 5120;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 5119;
defparam ram_block1a2.port_a_logical_ram_depth = 5120;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 5119;
defparam ram_block1a18.port_a_logical_ram_depth = 5120;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 5119;
defparam ram_block1a10.port_a_logical_ram_depth = 5120;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 5119;
defparam ram_block1a26.port_a_logical_ram_depth = 5120;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 5119;
defparam ram_block1a5.port_a_logical_ram_depth = 5120;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 5119;
defparam ram_block1a21.port_a_logical_ram_depth = 5120;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 5119;
defparam ram_block1a13.port_a_logical_ram_depth = 5120;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 5119;
defparam ram_block1a29.port_a_logical_ram_depth = 5120;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 5119;
defparam ram_block1a7.port_a_logical_ram_depth = 5120;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 5119;
defparam ram_block1a23.port_a_logical_ram_depth = 5120;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 5119;
defparam ram_block1a15.port_a_logical_ram_depth = 5120;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 5119;
defparam ram_block1a31.port_a_logical_ram_depth = 5120;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 5119;
defparam ram_block1a11.port_a_logical_ram_depth = 5120;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 5119;
defparam ram_block1a27.port_a_logical_ram_depth = 5120;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 5119;
defparam ram_block1a9.port_a_logical_ram_depth = 5120;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 5119;
defparam ram_block1a25.port_a_logical_ram_depth = 5120;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 5119;
defparam ram_block1a6.port_a_logical_ram_depth = 5120;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 5119;
defparam ram_block1a22.port_a_logical_ram_depth = 5120;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 5119;
defparam ram_block1a14.port_a_logical_ram_depth = 5120;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 5119;
defparam ram_block1a30.port_a_logical_ram_depth = 5120;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 5119;
defparam ram_block1a3.port_a_logical_ram_depth = 5120;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 5119;
defparam ram_block1a19.port_a_logical_ram_depth = 5120;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 5119;
defparam ram_block1a1.port_a_logical_ram_depth = 5120;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "Qsys_system_onchip_ram.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "Qsys_system_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_l9n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 5119;
defparam ram_block1a17.port_a_logical_ram_depth = 5120;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module Qsys_system_Qsys_system_onchip_rom (
	q_a_4,
	q_a_20,
	q_a_12,
	q_a_28,
	q_a_0,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_2,
	q_a_18,
	q_a_10,
	q_a_26,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_9,
	q_a_25,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	d_write,
	saved_grant_0,
	mem_used_1,
	src2_valid,
	src6_valid,
	saved_grant_1,
	hbreak_enabled,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_data_33,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_4;
output 	q_a_20;
output 	q_a_12;
output 	q_a_28;
output 	q_a_0;
output 	q_a_16;
output 	q_a_8;
output 	q_a_24;
output 	q_a_2;
output 	q_a_18;
output 	q_a_10;
output 	q_a_26;
output 	q_a_5;
output 	q_a_21;
output 	q_a_13;
output 	q_a_29;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_27;
output 	q_a_9;
output 	q_a_25;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	q_a_3;
output 	q_a_19;
output 	q_a_1;
output 	q_a_17;
input 	d_write;
input 	saved_grant_0;
input 	mem_used_1;
input 	src2_valid;
input 	src6_valid;
input 	saved_grant_1;
input 	hbreak_enabled;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_data_33;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;
wire \wren~1_combout ;


Qsys_system_altsyncram_11 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~1_combout ),
	.data_a({src_payload19,src_payload27,src_payload15,src_payload3,src_payload21,src_payload11,src_payload23,src_payload7,src_payload17,src_payload25,src_payload13,src_payload1,src_payload29,src_payload9,src_payload31,src_payload5,src_payload18,src_payload26,src_payload14,src_payload2,
src_payload20,src_payload10,src_payload22,src_payload6,src_payload16,src_payload24,src_payload12,src_payload,src_payload28,src_payload8,src_payload30,src_payload4}),
	.address_a({gnd,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!mem_used_1),
	.datac(!hbreak_enabled),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \wren~0 .shared_arith = "off";

cyclonev_lcell_comb \wren~1 (
	.dataa(!saved_grant_0),
	.datab(!src2_valid),
	.datac(!src6_valid),
	.datad(!saved_grant_1),
	.datae(!\wren~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~1 .extended_lut = "off";
defparam \wren~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \wren~1 .shared_arith = "off";

endmodule

module Qsys_system_altsyncram_11 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Qsys_system_altsyncram_can1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module Qsys_system_altsyncram_can1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[11:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 12;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 2559;
defparam ram_block1a4.port_a_logical_ram_depth = 2560;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 12;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 2559;
defparam ram_block1a20.port_a_logical_ram_depth = 2560;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 12;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 2559;
defparam ram_block1a12.port_a_logical_ram_depth = 2560;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 12;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 2559;
defparam ram_block1a28.port_a_logical_ram_depth = 2560;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 12;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 2559;
defparam ram_block1a0.port_a_logical_ram_depth = 2560;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 12;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 2559;
defparam ram_block1a16.port_a_logical_ram_depth = 2560;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 12;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 2559;
defparam ram_block1a8.port_a_logical_ram_depth = 2560;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 12;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 2559;
defparam ram_block1a24.port_a_logical_ram_depth = 2560;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 12;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 2559;
defparam ram_block1a2.port_a_logical_ram_depth = 2560;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 12;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 2559;
defparam ram_block1a18.port_a_logical_ram_depth = 2560;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 12;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 2559;
defparam ram_block1a10.port_a_logical_ram_depth = 2560;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 12;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 2559;
defparam ram_block1a26.port_a_logical_ram_depth = 2560;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 12;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 2559;
defparam ram_block1a5.port_a_logical_ram_depth = 2560;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 12;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 2559;
defparam ram_block1a21.port_a_logical_ram_depth = 2560;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 12;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 2559;
defparam ram_block1a13.port_a_logical_ram_depth = 2560;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 12;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 2559;
defparam ram_block1a29.port_a_logical_ram_depth = 2560;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 12;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 2559;
defparam ram_block1a7.port_a_logical_ram_depth = 2560;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 12;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 2559;
defparam ram_block1a23.port_a_logical_ram_depth = 2560;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 12;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 2559;
defparam ram_block1a15.port_a_logical_ram_depth = 2560;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 12;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 2559;
defparam ram_block1a31.port_a_logical_ram_depth = 2560;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 12;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 2559;
defparam ram_block1a11.port_a_logical_ram_depth = 2560;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 12;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 2559;
defparam ram_block1a27.port_a_logical_ram_depth = 2560;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 12;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 2559;
defparam ram_block1a9.port_a_logical_ram_depth = 2560;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 12;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 2559;
defparam ram_block1a25.port_a_logical_ram_depth = 2560;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 12;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 2559;
defparam ram_block1a6.port_a_logical_ram_depth = 2560;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 12;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 2559;
defparam ram_block1a22.port_a_logical_ram_depth = 2560;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 12;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 2559;
defparam ram_block1a14.port_a_logical_ram_depth = 2560;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 12;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 2559;
defparam ram_block1a30.port_a_logical_ram_depth = 2560;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 12;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 2559;
defparam ram_block1a3.port_a_logical_ram_depth = 2560;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 12;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 2559;
defparam ram_block1a19.port_a_logical_ram_depth = 2560;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 12;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 2559;
defparam ram_block1a1.port_a_logical_ram_depth = 2560;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "Qsys_system_onchip_rom.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "Qsys_system_onchip_rom:onchip_rom|altsyncram:the_altsyncram|altsyncram_can1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 12;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 2559;
defparam ram_block1a17.port_a_logical_ram_depth = 2560;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module Qsys_system_Qsys_system_pio_key (
	d_writedata_0,
	d_address_offset_field_0,
	rst1,
	d_write,
	d_address_offset_field_1,
	reset_n,
	Equal4,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	irq_mask1,
	edge_capture1,
	readdata_0,
	clk,
	in_port)/* synthesis synthesis_greybox=1 */;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	rst1;
input 	d_write;
input 	d_address_offset_field_1;
input 	reset_n;
input 	Equal4;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	irq_mask1;
output 	edge_capture1;
output 	readdata_0;
input 	clk;
input 	in_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always1~0_combout ;
wire \irq_mask~0_combout ;
wire \d1_data_in~q ;
wire \d2_data_in~q ;
wire \always2~0_combout ;
wire \edge_capture~0_combout ;
wire \read_mux_out~0_combout ;


dffeas irq_mask(
	.clk(clk),
	.d(\irq_mask~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(irq_mask1),
	.prn(vcc));
defparam irq_mask.is_wysiwyg = "true";
defparam irq_mask.power_up = "low";

dffeas edge_capture(
	.clk(clk),
	.d(\edge_capture~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(edge_capture1),
	.prn(vcc));
defparam edge_capture.is_wysiwyg = "true";
defparam edge_capture.power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\read_mux_out~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

cyclonev_lcell_comb \always1~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!Equal4),
	.datad(!mem_used_1),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \irq_mask~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_writedata_0),
	.datac(!d_address_offset_field_0),
	.datad(!irq_mask1),
	.datae(!\always1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\irq_mask~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \irq_mask~0 .extended_lut = "off";
defparam \irq_mask~0 .lut_mask = 64'hB7FF7BFFB7FF7BFF;
defparam \irq_mask~0 .shared_arith = "off";

dffeas d1_data_in(
	.clk(clk),
	.d(in_port),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d1_data_in~q ),
	.prn(vcc));
defparam d1_data_in.is_wysiwyg = "true";
defparam d1_data_in.power_up = "low";

dffeas d2_data_in(
	.clk(clk),
	.d(\d1_data_in~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d2_data_in~q ),
	.prn(vcc));
defparam d2_data_in.is_wysiwyg = "true";
defparam d2_data_in.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_writedata_0),
	.datac(!d_address_offset_field_0),
	.datad(!\always1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \edge_capture~0 (
	.dataa(!edge_capture1),
	.datab(!\d2_data_in~q ),
	.datac(!\d1_data_in~q ),
	.datad(!\always2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\edge_capture~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \edge_capture~0 .extended_lut = "off";
defparam \edge_capture~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \edge_capture~0 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_0),
	.datac(!irq_mask1),
	.datad(!edge_capture1),
	.datae(!in_port),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out~0 .extended_lut = "off";
defparam \read_mux_out~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \read_mux_out~0 .shared_arith = "off";

endmodule

module Qsys_system_Qsys_system_pio_led (
	data_out1,
	d_address_offset_field_2,
	d_writedata_0,
	d_address_offset_field_0,
	m0_write,
	d_address_offset_field_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	readdata_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out1;
input 	d_address_offset_field_2;
input 	d_writedata_0;
input 	d_address_offset_field_0;
input 	m0_write;
input 	d_address_offset_field_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out~0_combout ;
wire \data_out~1_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out1),
	.datab(!d_address_offset_field_1),
	.datac(!d_address_offset_field_2),
	.datad(!d_address_offset_field_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!d_address_offset_field_1),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \data_out~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~1 (
	.dataa(!data_out1),
	.datab(!d_address_offset_field_2),
	.datac(!d_writedata_0),
	.datad(!d_address_offset_field_0),
	.datae(!m0_write),
	.dataf(!\data_out~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~1 .extended_lut = "off";
defparam \data_out~1 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \data_out~1 .shared_arith = "off";

endmodule
