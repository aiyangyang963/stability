-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
obeTP/FeO75/+8l2xVDI983XfQn/RY7S0LRu0liLwrt97vJADERu1aKGOT00jIO5fUQayRjTkReF
x+JoHOhvKEr5t1M77irEUKx8rIo9S2+Kq6Z9KVsQqjfglg5KibBtaY4j0ebWZ+U3zxJdeDpJCh7O
tI3D7Rk+yoxRl815aTlwfTBayH5WZ5QZjL/n98kGioFFpbnXwwSBKJcXrOISTBIIzBCrnHtqkva+
0O700IUq1HXVOUp/areOatL0J5+cx48ouzyFBfIeW0Wd/M/nnPfFzV5a1869nSZVVl6lDaMsrPI/
OOIqd+eOD6Eh64u0yB6VPc/y3yIIziqF557MrQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11968)
`protect data_block
OkOpKN59fmWSdg6rXxOBjQH962O4Upv5R2XMQb0lvbw/REAtRG/Fnrm/Wy0YaeN4ekzM7hE9iZn0
xg5NDRXbZXwfKgLVxbhxctyc3REZcVpyrDuja9sAVCriDtVp/HYGM3cRuwlO9J345T3FUFJyWTBd
tap/m9zgclwJMRXAkX6TSqBSPgGjxdyEXfmk915DL8DlRWmY/z3BQ4Ve7m/MWrRc9uHFdnRkCHLY
a/CM2TZmOuSjSp7rBJmzuLiK7WOzQjPn6xNtlpFRCTrh3xeHxSCdcIcunEEwjphrcuhm7KvNQqoS
QaM4UP+MgDv95zcVhOr0F1hdW0dZpzaSsohz21pi1AXsrLoLD79DpwAb5sVCexWZK6nziKXfjvRY
QnFK37iHXXf4N18Up6k1ZB4DB1lHEaZGdxLUVmKPjewBK9SQAiY43DmTaGbu1EqVB+8/iAvhrYTp
dB2IAAlgUy9SlaMamNlN4oW9tTz1JyZc6dIDiaoKILaSbC0wE6fRj2hYJX8j4RiJCym4VbFjUyxM
pKt3I7mbGW/uJo0OUY15iKpoiYaDw4ZYojFE9TGVx0S/SdWRYkz1cyCSsxJ6qvVhxKka41v3+cQo
y1SH4h9JUJpsNYsYDXjdCumvKxc26ALkWUFb0cE6s3HXvb6h8TYUMqHLaetYy38EOz/z+Pm5S4rO
DUeepaNr1/+mb1x8eWsYM7D38GwsBX7jWAWj4ffO0b/T9+MFM8wLcni6YnDQf3D7wXTlBCI6Bcuk
4yJA9Jhagg7c88+pjVbyGqMkFUxMcMr13XbO1yyQi8I/AEX84LsYq2wXCV7J4yWDWUitMqPF39RM
S1M6OYHCkR3PTY5ITJCwxx1XBxn7LtX4L5zDY8DF1pjp6FDu8g4pCoEJdUtNF5LXy9lRGf8ksRnE
AlJAxTfPuriJlG+PxcqkOK9LbmsX2jHzdgIUvzF2dswB5l2/Btr/IpQVSQdlDFd6WnZCkOzszaRY
/yWpRjXeb0yE3makHJ0v9MVTHr9GcKCS+MgLddBBXDiFC8ku+cwgTv8bN7ikX5YMnS7h5VywRe6/
7StfaOtHO7Ua2bq/2kBNlmgtTMPSwsR0jz8ry376ufIhshEHuI/yVXI6MHNriA2T6lx6Jd/XYTd4
+Pq5H2T/W2QgdoiOBC/skU8FwLwoLaNDv1qvbZeJHHVgehCNFzpoygP3MoQp/LUrtSkVqvEu0OSi
w9rQquQhobIz09zEbwOoNJcR5W3au/LicH3j2UHND7+NGi4SLrsOVvC6KwO6L2SEAfdKa7cbxMBR
ENchzPiGe6YVM20FnaVB6R5lFyp1nh7OumHbLPVTyy2/Ela8wDG8bcrLBCtDBNc/YgCk7FNO27M2
fJmu3ZxazIXFtFFumDLwVCrUghzi8i+NzID8s/87+4Fb3qIsRr6UZGcjVRYjbmijmJmi5rxUz4+3
6F0k3KVXOxfIG1j5VbdpeXRaZAXepVF5uIk0KIcLP74ZR/l3dwh7bF3ImGWv7N+awftvvnWLL6Yl
9wWvCW9GzCkbinGXq6VlCBZk+Bhu3u3eOJ4Bme9RAnBz64en5BVByK2Ri6tSGgVNEbzDdSMXEz+D
OtxunuoCQPX+7jeRhQf9Ttcgoo9ek2jGhcA1ocL8jJiD5gTH7C69QCZ5wjaZRczcAuYEM7JyUgSn
MAiZfuHHwdh5xMfpUYAU0UTZMOSSgMY+GuFeAwEEW1L7ZxNODkilL+5tmRXq6Aw1do1YF94dkQQD
MCh+z5rZHMLFc8fyDZzoQJNe5BdwKGHTT7Wjhk425MAiKneMDUZVJn+LZ07oYAu5ZrObm5ey8IwD
QUA1SNv/M/r7iYprmLEKaWCSdFmGB+YNMXzItoGDQlzip/OPZ2B6xdpmYoyPFNUai8Oixkj5tPgf
cayfstNK22JZAzW3qfh8YSp3UVDSKJfgYbJMVbvkG79kMwtyhklqfahHLr3YKrbRMpBjV+ltojed
cRVLudhNp1SE9XWfUXn8SOTXvh+zmnKKntgY4v/PpMNrJnAg0ccuCtIxU9HnXcEiPgf2rIG+gNuh
o49zIQPdKRCUELhWtnf8jEk9AAgLPc8g7Dk4EZDczZ7hkc3X42HWzlSH2q15O65HqeISoXM9QlC/
r4mVh+tk3d4vwinUlsd63GPVrhBrtLzrymuc+Ogs2SkSm7z65/1rB35sSduhH6H8pwmriF3xRMyA
EihHIf4a0YZ9VPWHpC0ow/sEcV3KTCha0JU+4zjMuXJkS1zHqrv0aNIrQ/wyzB1/hEG7MQDBduTT
jvYIQyfTr9VDECQjTGJqQvPLLib9QU8mACPWnc5PYaJVeQgfyD5XXHnKsVLMz25TsLI5GivcyGVZ
VSRdTN3coacuwG0btMuptVBRHb4/IIf7nAYe+UG3qbnlbeL8xjb0rF070S0J5ajtm8MkuetZkGpV
PG00329UAs1vPUMJV/c2bBkYXrIrOjNn+hYmlqYIWST8imr7srgF2nuZk/gwJKqmqvOj1CGbML7D
/ABfwscmKk+VnsSNj+EjKNr7QOv960aMmT3pJi5BPXj5Hzle4jGrsQnLIcFXCccZmYrigq1F1wQt
dFLY2ew+5Wd/2I+OQpTLZCyBlbO4iPG5iyNvtuYiBoMqv1/NNX+bF6u7RIerzc8cpxjJHng+bXZl
sBHe5sqVR/286hGJ5iFPMbeK4RkYjwpnSMFbQ5PqEna0AV+MGKaEesH3K2ITKGK/3DecLKhtmmO1
teL8B0f8SznQlJKh6GSAYTk9WU+Avd+G6OyWg7ss4ivYd1Mkm0NKg5qU26Ok41hXtswcxo1wCXMP
TK4iE+HFRo+XvS7C/ZL4QhrY9KvQHize5F22fIY2nk0JYZc4pfUl+TL7ptiAq1kleG5ZvzW5mcdr
hYVY2ZiCVe1sl8IddQk2/K1GMDp8mXRX5LIdGGMjLqWwmPMY43STOWsVpcn9EAnpofHTMz6Z7/39
7teQEt3RLVatlBlfhqrGINHVDu/FJUPXMPH3cH3N3ZNJsvrljm4DL2kkKGpk1/cKyF8VXvDPJtXs
KVaFU/LzuAHdP7OhkP/h82oihbOWZwrpBR4hqTdg4OvCxYw1q1/CwurCpu+x7d0L/gf7o7ZU36RW
7O+n40SLghh/dOZKoncFvlpIGt4GOc2v206mfXIly8zcG6R1PpqysIzRsYjZfHs50qJuyJMDtpka
HMTNKDSUIiS65VQc3bIbNlC/Dk5yqzPg8vs/hMjAjXCOO1pkmp9siZoQYcqndr9++XoC7f8XW59q
t1T6G/0rVcZhFRth7mJHl9tlK0pl8L1IP3ECVG1DfC/D8CWMPU7XzpqXhZ21fAvOXAtNXrb0p3ru
WbkhiZNMA3iW6lFHqIrJ5N9yFx3EMl0aKJVU1wxk521rVpD3SqFmCmxWi2fVPWd9rlxsifUkdHn5
UzlwGTIrQBdZP0VXDcCWjiRbnBbG2XSBniAqH2xh9AglIuEDAcFQU7jPUHm6a4yUeJzoVbxzlk3Y
6ajCCY5WD3YY+y8MJ4dAgXggfCn2jYyF0lErvGNDMyO2BHWVfvKNQLzaVnnp9fWcL/bC0k0N/o1m
PBZPzMeYFLAcPtldNnKOhbYBU1Ezxt9lEhGRW1cDoHaN2eaI0km/RHUU2vqbg1KhN4uR83W2xNaa
6Oz1cKuMNzGSrKCQjHguaoKaRlwlmZatryGzVJSJj6kVD4wjihGt2B98++ltaj0/nVVndYFg0/7m
3HNEv/SatEiqe8jdOkNdEMZ7zkD/n7/IL1IEJIJCST/duj0Uipymuk8T9VHMmEwaTHIc2T5Ibfc/
fLPEli3UdwHT570Urd1aJl92xiuXJQApD2SSgIvCpQBUT5h1ucuch2f5cIzVT/xB7G08UrbmKp0I
boohsgXrPvqzzd6m7H4FnkidvGDGrvobuAyI7izGUbFQlFJWII54p6bNQq+gOqN2z5WgSQI4Gq3W
avSVuKDJLbKrKpXxgtpl/rqKoLqwMwebnFtfEF5+dMGXbeH6PyPMNZTi8GDw8JJJ9X5RZcnpeFTv
j6qJ42lAHRm484Y2yCb3CedwOrKeHXTfYJNnCNDGldQY/yG/OToNYZ67lfXEP7004JyNvKLTzujs
xSdXL4ZNvpRHrdH/CqnCyC2q/fdGajGVV7bxirQGQwJA8zdnDh86+9Jw5vWUq0AbPYDsYqXCl9np
73j9Gcf5akypHs/8n3oci6VpWu+b2EhI0i+lTlQpP0H4IC7sM1LjaEjuDsNcesJ2uvIAbSyTBbsg
SDww5ACVhHonkVnHBy1ViOC3WQUdc/3pGw7tRt5/hmyJixsZzd3JvaKVAGFkP5Xbdr9WsrK1Uglw
MgblSiOHzMqKUsKBdiIy0B+s9h4RmZL+doTrutIi5qsnVI+p+exBVAs6m/477yw2DwOEAT+ydVL4
RbME01iXg1xDQ4AxexwSEmw5jUrmSP7Fu1+io3N+4I+Ay6r+WaXPGX7fGXsMAh7UIGvORF8MSiq8
f+/YgicUZdSXKsN//wM5JgWF3LydqgoBvRuSs4mxLE42kf5mZbXMJUafyiNSXDZW8KNMGMv6bC1b
QqBmWgqhKCpBsA7qLJwkDu537NjTSL4URypx3pQt7VP49GPydiWtwqL2c7cuDaexzpjGg/wv5XK2
pF5hDzZp7LjEAcekluuGkDt7XOKzOd1Pn++9MegEJi/0Pu4zAA6SmibWD03lHyiLJQp1xEqm4oaG
QGVV8iH7ljF3qtC9eJ1XCubZSz1kwsl/S6xjggAqL3dyMFjGtU4xa0JjmkSXMOAfoUMTt0UglxOe
uE+5Cg/fORL24DUg6lsS74Csh44MYa4tjSv46L1P81kMOS8qdjHsV4J7cnkHs8QWVfgDcph3DGpY
CPSrOQx3FfgGl/boTeaG0FQO9EvSCl7mYJj+H3vSvZ9OhkUufJ8z7aLCdtu9KYTLcoUDCXU6x7ii
IhLj0zIAJmc9qD6/sziVU0g3HAYTghp4OJBSyATy/AEu4RthNDC8Qdn532m3PK85DQqv97R3qVc8
agmoLNyxxw7Z5E8lCJueBHXiHCFoB3SsMQQySdFLdikEdDxizX/bbSeogEfihFA0zIKIHU2ytAOz
7+bptWLXQLNRVpzZfGqwZmXbCnVe/hu0fZIL3096A/NlG4uvyRqsP2zPrNdeJpN9ZT+d4Cnty1GF
XZLP5ACxk+9UoBQujy8zsJDvB7suA5E4LuBsjNmXPxKNvdDceFTiz1jWmhMcQKNQVHDJfB//kANM
eDkkSFkPnpoI9jeZpso/QbReOr3NqXgy2n9HivColzoM94Uu6JamkcpZxBm9w5RV/NNYngHWPPU9
IC5e1AzioC7KtJu0ibJ57TrDBaI3shNdri76xNbbVIdMmRKeh5mMdJFtkqrRZ/qrV1VjAgvqC0bz
vkS3etrfUL9HHfwoHic/J8tXkHQlNWES6rMz8O0sDf83LgcLAGG561g//+wEro6BIZONjuCporkt
lZ9iqzrmxcFNrRaSrb2PNUfxiUQyg/sZRoFPcrR0fjE/iGhBSG6H3n5+dxyQ8nkOaKD0a5TphMcy
zmhB+wcWhC4xv96d9U5J0N57iFZGHO4rLEqUE63UFOddrgX8yyjdAAfdK/vunqeBTwL8C+AU2OOu
iE7P+ung9/NZg1+0Ccz/ebHaMClev+1h9GOCpAU6X3K0Umzt5AMW64u15u7s8yJPxIIwPUvm9Ect
OcIrbUiWlKu/TaNRwnfR4shaIeUUI69QeBY1GpfG7eYQak/Xzz6mfOYS+FyiEf7JvLqlBLr0Ye2u
JJwsEsDQL+IQZCW4/x8JUkif56jTJscUwRanhyOEyDnDLYCrCWfwXOfD0KrBWK5ZppvJkNKIF5Vs
W/JtHtyUEwTESsnv0cL+3GqACSrbx5KCM2eAfzjfHmF3UlQww/eKYFTdHsiI9QmLhqlycSk+7BAH
ngkKsW1BXGpRy+fs6Qxk5Ws+V3SDY5lxlmba2HWXXUu9e1KQ3rV6/T0oHdTpI3HMNCXe/IKXmb3O
rxTivvL7WaAInWnrp/5gSh0uDPOkAZkw6cyuVFFOTdP9EV5cvd5cJnNHIZgQGehact927ZPv+kBE
BGKpd0VSR+WIs9bmCt9aCNmFgHieM1cLQt/5jZmKddtRymoItyKGWWil9K8whZfT/bLVeU/VEeJr
1SN0fzN1FTyQHLJUg5DdTX9rpWDm4hHnh2DEqfVTR+3LJFQjiQ4eGENcRWPatlUtRfjGOkyCSRPH
p9zPJPIDNLg1t5wdMY7MpmAhKCF47MJbYP9hSF3sXamW84mZiWtiFcLbioJ67TuxBQTaiVXLlLf7
4XO8aWcqgie0hP4Zofg0P8XdbbAvu7iz0jrhCgWX+f/1x0z7BTpfkXlmUcUgDyeBcMn0z4OV/kbz
x5Uta46SRIqNYZKGfOiHQPWFBUa2F9pn04pxAgjdvOCqkmSddknMXuXgb1RC6KCoGDq0HAVp+XhP
2naAL4iCUxBL+FnP0VO0LferJiweOA52ZvCqNcCJWQntQEwY06uY/g0e1r2p6k7SpUUXSSTz7Sg1
/TJL74Az2UHvvbZmMNXTs+Lq4vbZ8J1Q5nAvIdCJ6fmuIlCPl/dB7ZCzlj2usvFzbv1Cy48X9+2B
bboEYlF7Ey5SSODgPBxsqWVQm/GSgGNyWgu+/UzBXqhIFD2XqJM+qkeJWEJSda3P+/xARKJ5iEuQ
bS6/CjC6qnNnJEwU7hGC6QGwABT/r/Aa9iP8jQ8RlSYj7oi+4p33PIHD6tr6lPvmqHyKLdmCL3Aw
K90N/Vf0yAEkpBuZSB2l56Sk1ZqL9AbWEE4wx7JJM51LeGkQRXQ68JVSw47/UmH/tFrzzGola0yi
U+mR7O694N0AbCTpuAlat59K/y1FawZZLkDeFrAhmSeurxEyTWySvfk/+XtqqtXTuK89z4PXWpTT
LIrX2r3YZbO/uz7Hdo1t8dUQrIH2LFNwqMouXiSzr8vo2KDUYTgYu2eHigan42R4iOocXZJU8P8/
Z0RBTVg9+nJnNHGAEryOodvHJUmZzg9hWX5FxmoDj62jweHaxlYPN/AD6g41vUgISmo3Kfqtrs6z
+UMe7NMO0cOmVtSGvlJZjFGcMsEeFOkCRcg3l7BKt9ik9+cnbjPc8yj0t1jrrLelyHC4OTNKJNB8
/GvkxPzac67EPGo6JTX0HJAeEQh58DY67Hpz53TYz7RDbi4Nl4Z56R9L2Yeyk84g62krHWGuyMx8
52CG7MY9ImjZ/314dkBdMwqc4NevsNKnXmCkW2XqNQAjhUJDkzY5EdI6pOqWkZpz7tKSgdZGMRWs
8AKBm7nVH7cS5+jaaf/Vl48oxuFgPFnnaOAmorN2pmoIA50NGC9A4lVD0mqjflEFWy12YS95uYVd
F2ui/n9lfsTIXYmMumGUTDO2Qi0rVXd3P2O2VFYdbxVXXtM8oTuiGMevQrSUFApFuUOCWs111Giq
X+ShM7JiUDL8iJYc8mEH+XJFir/drxC59p685ZBnp/aqDVzoIj5JPelVg/24Kgu4Ib9DFRuEc8Ar
xg048N6LeoOcn/vU3kCU+jLVq53Mg1QHZzfU8nT2NJG5HoHuKLZbkPZ/yExp9KdNnQtbCJVHfZHi
/NVYKEaN0eRdbfbYa42RGqe9OTsM6K+iM9uWwHCSYp/IAL19s2ho390PsSLd32pBW27Kmd8NT3hm
nqsRLGrmMIOLcEtKn0IJwSGpjBmpjeTQUtUest8hXF1k4+weZfd54lm/TPlkdY3HbWsHAH5sjyCD
GvX7TNxYqkfer633Hcxo5+6uNioDRf8QGFbsJzPa4rb7OxLp8Spfu4ctF+6x0IPMK3bmP6UEjS0c
GZWQGnemPmIdgaYmbA5j6dntnQiwmLRNKuHSUILt9VpU26+VkD9aWWvVH2UVeTYvd/Bi5NvhvQvN
D1B+fb/lsHOFN7JtmW0xRQvDK8K62sxFSQ8R/mLmWaQesDPSnYqqJvVK1eGBTWTPADUxs1RDv/Qq
nLhbb/IREu/vf7n4fJKWp331WEAODoUNIklnkkjkC+emMF9FzCgi9kRdXL97dtwatczGkd6TOCZ+
6bfDw80MustsekzT2FgtpzKgbdBfC+OSQQdKaih2uBr2usfALzUm0ebGY1ez/tIzO0zOEo4MmwBT
G9EQtjoyU31U478RdpCdVnpnsAlqcjYLmIo0pNTptSykkw+a0EL1E5fP+VphhAN01jHFq47a29AW
ndYkGxU1IGKK38JEG6NegKMsnlzW3vyJLozaXMb7tFRvXUfEGZGkhBIcBas5rYo35AxEggkNpCS3
H+efWScgTVKOwesF6dG3LfR0p63QnxecWMskoczd7/y5/AYl25XHhEE3QvLVx5ycjCRcd3HhJXGc
N31Iru2W/eoaYIP/qHbQ00kfyZXyZjoHhj/s6CYquN1ZM23QYWui/1bie8K30gFA2FQJSRLqgc9r
C1RMeMpnkK8PvLCF/0RKw7bWSZ00OQ4hfZfjn6db+izjvp3HNnwCMe8ff+jgoBMRjLHesHF2QV3F
AM2XtfLRDdx+Hp6l364ey70RPMKxad2joZnci687C+Uq7XiARKqkYIAF2ZvHK9vaqEIsjGTLnsRR
eBqYhT2103JCDE1QYZz9Bvf415MzhUiQUz01ZT3u8vPgPAYU4JBDmWQX1iy/1qhgBtsk8xiP9IjD
+Q7Jkur0ddeNIBRT18AK+Fy0z4HoRSsus08g7FhgbIO0KQzBVq3JB/ZBxFsBlF43RpzRZc3aTe23
iO+eQ3Xg76nQYo40Z8Lxe88KED7igBLAjspPlJGKlC90A/bCw0lM5tB3p9k0F94XA3sz45GrG9m/
bhHKKEaZVD59EOHFih2V2/+A7d7cPdUxnPzZsD9pd0GOR/6YPGaBGCl5LK8H8oTUUUc/Q5nh1z+K
U8d6f3V3yG/lJ/xF8NFHpiX/lONeUSB8GE+2CYWhWUPZRMPPYwpsGiFDw/AJvpvFVAxN4f0xJlRg
Bhsna5Ui5M6hYwL+UaPPF45Ji4ISRaQr1iMhuLWYdRwlBlzNYmmBoHb5kLW41ogkL6vgq1O4zyqb
vlGcI5M3rtyqQ4HH3V/YExVEA+j0UkDsIlwSLyE0U0XNkqbPAsI7GpZ722TfNRkeH6KS/T7kpi05
f2enJxta0JmioBKyVmFqdQ7keB9REfiY8H5FDODRqQDZK3TRVKEbvH4CZZJE3rqWiiHGrav/buLU
Z7aqlj5bmg7eMJ9K7DfQO9WJGa+jzs/IFaLnClPCzKxODd5NRHZbB/CmJjitKiCvabEi4jzUpiez
vZY+49RybcL4fbJ/WsceomBV6Hn/dHobsUnXPUC9GVr7B7sg50QMDYwYY45hbMnSEOIqvRSOBH4p
0FhWSXb3G5TjACCeREKhAuUk+yA4lF+A8ZeqSStkxO+T0TZrimp/E0j961IDqZbSOf/cAuoRveHE
ouf1XLFiTwAgq5Zlb5eJWjDwPnuML+sMrk44bnANB7tRsCWbDI/nnastBJvHJsvm1yaRzw1BqPpp
+mGWooShw1vvl2ySdG7O+qfv4lxVbaqRadjV9zTcFQDblXWd/GkLTsWmVppicgXyMO6LbHYxfnaE
PeL+4SDmhePmgCO3mjM6LMhksvT6Y4sLlKIMiCmPuJwwf6wRMik2tSNCl0lYCs4P/UcSlLmhzV+Z
Uq45XEH992mvmE8AzRsnGLnzlFaxh0LNnmLlbL5fTCG7gvnuAAJ8btwxTnE1nStL9WBxI0H7CuNj
Cw4GMmnd9YEcUaLJUJ7uvU3UidLHW+SfRNulu+U2l5Rki5SRKVAkQXWq2H/W21VUZyG3399T6Owy
oQaM8TJUki0kSDfDKOURqbL1cPz0a6DDkbfwTuByEPrJWojLuXstZjYi6lZ22Led0G5CVy6wJpY4
VmiQE8PuPP+CGYAJPC21xhwdiAQVzRpslOrty9e/LE2c4HTMFzqNfID/sADt6/8H36Fr3FD+hgeg
CehUz/Q/XzZhuST8+jfWzATb3Ok1bBb6zXq9FSzvXAl0CaKdu5eSppFey/pgt9aQGZXPpBi//q60
AkthFFeIX+ogasYBCCkn4PA4mgiCM2WZiNW9GXLiuLFpOLmt9DEpPauHA+APjgdeWcBh/zOOXmIy
DPsLebIG1If3rlHFyQ6eLXMZzXTcyjs2LpdOxPZ80iyN9vGxsTllGozilPgfK5bi3WmGHBi25Hfp
7UPf9jB58qQ6FSqzDgkxttm7AoBvtLDuk6C5/fpEbmr/oMEONMEf/wyRxQjOxWqMEsgMkA40o65A
snUA6w5EaTwrSPAPzvhil7lecymwIGdpDv8eDqTdqf5RQRDHa9xY0lyt411ObvNxbp3ToTfcQk2Q
jGWKVCnnXzE9Wy2RKTE0ghKsimJSCGwRMoY/oYt+k2q3eB5Iq91d2Ly28GJyZvp8TnPlqc5VPyjp
cB1RoHQInUClMl0WaAY0GTD7lqBQwqhuOBDvjCiBOCayur9apJH5XyHOeAlcIGxf8Jj8gaVEDeZK
oVWtqRNmLnWjMtGizkLdA67QgMUSzO2OXRMsBu/PQjE4F3w4owAnLSCDJn2BQCwpZBbfnwqrV5vf
F5Sy4y6Kti+8U0h3MHB3ZEZ6w3vOm1IWNeT4yiv/7qTvXDwLpEpnR20aYdOuONH5Vg65LEYiaajz
+vyXISHFv91gq7CdHrbYtbtzY7NmcBys8W6YCVYtvQ4lygffQXoe0XbgYFemlCB7wPLDjjdRnQEo
j5c/uQnfErFx3Yy/8sneIKBHozznpahd5X1WNvQ8HOlFP47uz61lOfN/FWx943gNooZdUNZGqZUp
GFmPBr0hHMH6jzWS+aStcnw/FXgrmtx+OXzQHdAxWpKRy1x9M/Ix1VbZ2GWewQlJncAptxj/iLYV
uJ4W3H+EF2OqQStbX1C/v4phV5vgRou0eorKJQ1LhecA9zOuz5eq1IrWiLeCW7BQYy1jfdIHQSpr
J7A8VNzw3U/5HtdsiqPc9qoZJEgi1ejp2FPyr+6Xs6nYepZ3RIO95ssBi8K29Opmvf+rTk1dy1cg
jecZNTufKlWja66UwkxMiHO6B0GnSkOqc2OkyBoNONJO5cGucPUC2sWzo0Zlx0C56AhXu+mrs+JN
0actYTSPFYvjiIzPUQfOAAmr3Bk7KfKqV6xd3Df+BWLz6L/U16DTDQGpcrfJtsI2kBEb/5XsAgPO
ptxTyW1d18y4b1Hkws9Lso0CwGS26LCdpDv5APfr1sr+G4t7iLoj4qXW41j2htvmfZazTctpIBUs
nxCel6WuNUbiS+IwNeq6+U+q28fN7t6qzejUdvjskzA4InBaRLC4wb6fRE1Xs4J7cjeinpqLkX2q
imszbdFpuUfEeWSUkhev30joRovQPOs03SB8q+TzXC8r2JriH/NVBC+fzjRsvbMpO1JuP3T7M3qr
MK7b+Furi6bG/924qgsKJg/m3Ui2vwLOeKp+eVXQbQmTSXHvASZfBOtnFTJ4J5bqhQvr8zfZuQjL
TusntH33L0KvBPpk4D/xAJblr2R3OknkrGf2KFwdWt+PUIUjn3cuRpasjxFLC6BFv4h5B1HKbPul
DDpSvgqnOIY4mzHVs3NyOw6S6nJdsXZY64nA7iLiP6f9Pog9b7gxW0p/a6s+z941F6r1aXIPvaBY
9GmFF9kxgJkUG3WxOb2EOvNR6XtTyMDZFO+SNFi/oE3c7EVMYsJmex53U6WVmmcIqRmN+zCB4p8D
EPmqcXCemejhjs4J2vauZeW7mOcYqQUZSvHGBTHIIFstIzke71BC5FUEb5yjHmmi2OZmztRGEdzl
FZKTmM1NC4jTT/YaLlI+FrWXWVPiCdDenOrD6mm+ewC9xDlndKyJsRqd5OCEEw7BXEPOKjKwuNVI
Eb54Ed3II15dzJzRTK1rNOSqJ/IyVkBMfBj1wQH+LC5o4Njy+pmbkUDrAEbhXSUD6LHuVMNwZ6Dj
tolZ3m0ig9fU/VlGqArwRCI47zQoNk4UlcG2Xnd5hYeTbVuzarmxRWENtPFuPeL33obIchpo9MrP
06ghqBDpBHoDp20iatYOLxETGuYz5DG5dgONuX/sJ7mJcUnMnJcQOBcBm2hWoEOO6Z4MP5vKxnAG
9n1/9csu5H0yNsyawlNdjr35XyFF3umafOUHClSqmV50UbMpEARXP7WkoUDZcQ6ENL/ETxlCtqt9
lFvYQsgddPFqDQhWAyZqM+CyZliePenewXX8ComhtGguZkBZ+f917vAQyAqQaxZvtN2c3FSu5OL+
iRs/bIkSVXBhecc9x2LfUzNa/Ao/LS6/hgsaGYLZ+5urYXDvGX4QutTpaePPlEIRx0Seub4+yvcT
Dv557biFpPRLBWVJNv1RuvywDqGr1k5Jp+q25TP18TdHuim0hidxqbcT1X/3VZz5pLBLcQ4s2kR9
K5DIc93vBOKW9jbZnOvC0/hBBYxHpqRAvelaODIgAdAbN6A4OESW16mB4Gxg6mmZb+Ks3jkAsl55
hz7X5p2j0eIfFTm9wT7bmA/jovd0BKt/tao9q5Y2egcoD+VzJ3FrKFwNTFJA6OQDaEIFmaxM1Xfi
073C+8eCkskD0m+vJyo2uSM3O9Tz3fJ49Lf3LZJ/xMajdwrnXE+pSU4OQxTz64DBdKJFh/+4wa5p
MiqOIrsgEL88R2Wn4plPwo9Cfvtpk9+SL9zytUy1bwZJZPnXJFIUbSG41Ulg2C++BgvaqsEawqw1
jir3SLAkzpQNI3dzeUvyond5cdem6aiI9vqTvakD0+L3ls6U/SszOPkJhFtZw66rkbKAi1wBFlGr
jTrh7GiZ2g9OqMvM3Zr3Macsj3Q0iEpGMG+VMNzxxcsAYeuMjDrj+ASTulvn+MRV6gyQVlvTmERE
J9UQW0FekNvhO75K4g7GmZECm/AFBFrNj8LN8gxgG1BoX3+CdcMSHTDOsejCgu8wynWUtC1vAZkt
XnuB4u1WJIzycTP+ylJB90tIzSZK7ulNJdT05MpxHUR2gHCQFGoBhOZ/HkGZrZawPOzmnUQVmxis
Rtg7wJrt6L24lg257zH9GFZDuh2ikAz90OLoPYZ2XMcmhvXCq+9iZkpxd7afqp0goioPKJzD0kuO
iSVr/8oqTnBaXeMqXV8BP0nq2Twfjx/u5WTeKuEgNStTXelUbFGdIiAuK8OzHfM9OaTliKpimfhb
r9mHGxSiDdEcmrGE8cW+Cyqu8AEHkQYeuHUQir16RGx4iJFiUwRhnVWXrjam5k9OZz1oe3934ouk
8p2gRnJ7dOORZI+dVu9vg1xcyvqv9aK69iByT+J9RB48BqsL5zjQlOjTCQGslSS5R06nw4QECy0N
zHvunS6VaxAkTopJ/RQPlXIaEV+/epxD8WuT8zpjYnbLX7vUBGQN+rZCjDUVqgHxS5MZeUQS9QZm
SFmZKSBlIgtxexJ2xIyl5tC36n7auopiQwUgqCRqGGpYusqa0eGkWkAxNc4UaJIvyK+a09U+JRbf
Akz1ukywpQyxm0p36d1F6H+CICCADHDTBe/+MdDD8GEC4ngMaDItKVMLSTHS3J/mQbScMpCGXodv
AO4OPUAw5/MNMURa2fpJs2JEet6nrdgCcgtdpdmBM8U7ZtfbYnJnPsXeeXAJpvq4odYijR7TFtna
A5Wdwq6WmEVWs40DnkjE3xlr6ETk+oSNpLACM34dbusS+zX9mLfr+5ohBwqTAnUdo1wLQBrXBQOk
bueCiBEDM/oR+6r+uwjyuFDjX+vmlx8k8hxUnNI5GYFdEgr6MUGPxbKmcuudcG1Buty6pjGorSwy
kUEVhqvneURvUyghlHVcNIbie6xq2zAGv2om3BU05nie0QCuMiUjM4r4Kawbid798opR5r43sghM
1n0i8mwLg/AigGoLR+sonZvlC1xTVGeAZF5WTtLaFY0EvUY5bRwGcN9aYkuUBnKzFcV/gIF+gEiS
fuSM2MSSpNoccI78HiYxXataYeXQDG0UHePTvz48SVA7e1F/x0DjkkYCcr/odEkoZu85lo4gCLyu
kZn2R7wmBZfE4Y7eikzZbST4scyYLqZnIz5EaVCdEnpRSjr3DIF5YTm+No+nk86TVEZmbk2AUssh
i1AaYcCVfn3w8aCHYjrFuxuKq7J7I+Yn+Fu/8GK6ZtQjvmJHr9weJ6ZDBvelhuzKy8+oTVFc6QEA
kvSRmYbLQZRqz+qW4/0Z8ee6T5fhQkIYu7IStSLxvBuYKrSDJa7akbP6rCs+9bTLVLwsr2EZ4TlW
Lc9tm+gx04ktkSVUkLB4dRos8trYS+ohrIsdx69a62Qw6qSvzm0vw62DiArygIwYaO1x0VADZ323
+CMWDm1hTud6QnmvZdbyQieDMchXW3wg/dxy2CLBOO/O9GuB4nvKIT30ACjEWSdTg8HvaseERpYe
v9SW/rMQXgFQoMM8rCcV/0bobEdf4FntPHkugVYJbVG8LcUb2uTdUSIyXesm7UZswRPXcOwdRCgL
n8//29OE381a71rksRImu/G5yKUuoP8/DFMMb0X6OhubpToHlrNXLhZwxZzmc2qEa5bhiO6F7ELA
slLiSeKHdTcqicpkw2bkQX+5AaT5U9FfCP5wPJR3wtabSA952EaCzQPSIDcluPRoie6h/XEgyoAr
X2vQ4V7ebdrCCQh9kRMV5yqqOFUR3ty9ydTjMOOqL/Oj+DvuemwxO9VcG6L6ZYvkAkRHciARjb8+
lp7Ob9dfijLcob/pBrnO/qjwxnLXSHl/ojh+EXcrdUWwhVAu1OqJ/oSi2/zt7f1821QpH3WxpdL6
E/Vceqg+GD8f/JCHnLKzzY57zdUXC44rafBSQrPaJiyRbaW0aQVu0lxvUVgPXeAyJdo6sFiu3JQp
sad8Igsa7z5Im4+4jJPaLTHLf/YxnyHuDBDSQjygXZUrTGfu8IbaxLkn3DCRdL8f5FlK708jwyda
8vt1+cYWgxd9StiiTbe+JIAMnHN+EqIzGt0+KJjRYRZfwSfPWVJxhBaZztpysYfCBO2ARNAvTx/d
fpEsmuxxKHk2FroeJh5zkWHcbWV8lEi4Qe5lAz+SXdUATdQ4uzqPHkxy4U54Lxvwdy3pM/wLb1aY
CjlAMK7mO0AQG+0MfA+qWDQu4AypujOgKuemQZBSEDon4xpwWN4T/E1SU/KhGL8p5GPT+dUKqXoX
25FjX0iJz2bHgySX1DPzDLROexz3R0iwNjvH23N4VEE29N1l8clNV+3HdQe2bDJ1xlZJOqfMtnEv
JmWHHUthJaB61hle1+xgQ3bvt3qN50rDPptaqTCCtOSr0Z1/g+OSNJ46bK+pZ3I42gz9ycwHlQqD
b21DQ5yrjA6kb+L04tzpl0SA/PVWCbF9j8SgyUPXEqqfl1q5eLOVsfoEjHeVwCUjBFuqIq6cosaM
ip2VG6IxO0hoK+pdFodKXkagUs2EIBX/i/KuyDX8hGf/wdNZHEBnIYRL2UcWdCgd1rdnhzrSJ456
u2hfk0yRaIUUvNxsV6itDtjBMv9jJgYLGUChUTFdVNGGhkhIL/dFqr2f3MdM9BM9jz4DHZN5F94N
MWrtkltb7K/noDfbZj9EOiBRlqr5v6SKjLj+O0U1BxUrul5JC6sJ/AcROIMM7Tu9BLo9BCp/edtM
3Yr8+HXp6XKWtRG6CkvwNfSvnjVwP/Tdfq3uNYwmyurGHvml2IinKFwivpzoaEa4AL2wlNkuc4iQ
L53NMMkoBWB0c0tiazdm4CPwqEmLzhPdAsvLwHYErxpc8vUIG3HkD9PPbIbqNkTflCk8Qj4ufJ1F
xE56mIdKqM+HFmS3jkF9+ZL4SroIaWd/QRx291vwA6BeekKRn7QPVSDqJixlBr1Z+6wXm4m6In02
kAEpaIOZDeOlVb4DYLM4Vu43dEhVYpTuYOfAcIZJ2rdfYDmDSysxgchplj3sZ8pDbZ/+yUOm3l6X
INiQAyxfTYXh9/NMDvvd8IaFdUobOkQSSAAt1NZzoWWpfm3VF7x1ZjJrC5DoYpXMoi5xzq3HZQ==
`protect end_protected
