-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
n0DpdlwesPP/gyEGGs25z2uIzkxU4tQq0lDNmrfl5WzncogfD5gV8kOiS+QoHPJtfh8BglGgR5xR
gLcCH7VSAbYq+/1EIXBqImFM/7FzDnlHbxCyoN1u2yY345Vq3kU4qjmxL85rLi1J+8PCBANfI8Ph
+YAA8HV5hhkncjqnN509NEpazBjKtu79r3Env/EmGrpIBwIcKqil8Vo1IUVRWAoMvDUYMNLSFatb
17utWbMknTwod9PQ20hEwI0l/0Rh3uZGPdeVTAQxgiIqspEb2a6QR0mUq16FSPUhkNBA80Xg04Fv
ziX0j8Xtz5jhlbYIUza+ZFcODkM4gAIg9kisHQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2960)
`protect data_block
qxWqgi6Bdt1BOC+6iI758nPoEjQeNw6n24xERR8qGf/QW8LqRgg+QSaY1m0Q99PntjDwx8pUh1Kw
BMTX4dCwooREAsgERR0h3PpuzNlCDU3+h676/tSin9XloFI9wnuiJG/zgnq1HdzKQq7WiWW6+UqJ
5EBkFMuKP34j2TA4/4k144wECfxLiIjg6H/FNq4EM9k1EQ2jcrPTOgaP6mdlpXMIhm0X1lsaIg8p
jVUK2EEENRhcCwLRzSn3KY+t5m/tDAizf7ikRdmqmtzJoi0qSGwEgEgLZvdZ3KqX0u5rj4ZiWFw6
Lb89p3wWdtuZvRkB4TW1np6s0PCFTevKZpY2a0YXEGjqb7op0SNB/HEwunggAv+u58PJ63Q1hj12
0sPuFtzypLcCZUjNEckjUyvuf8iMO0RwBycj2PUrgMCmlV7cSF2vApqrqdPtLRop0WNozk5EaQJJ
hoG5yUmeDpna2MRD3ZXSVGcYPPcE8kBwGm6JUeQ/7Tn/+Jr7ChoMQPMS/SBosHk33uUhrXNa90JH
heDvwG8U/4gY9lA9wH5Tb8CITDoNvIgFVEyjg3H6Q89vPCow4b89z/dhtCxiQ6FfPk37x4RjCcr0
tYDokzCZTmchCSK4po/4U+/4DbEHhjJvVOSD7lGFQqhDEoDZUXHrwSdxa2c0RkWjTtvYgPWDeouK
JYSDd0cMmgcPrrrrTsaQiruG/RQ7lPtB0OLteZtU1GvILFNoUYS/HCbUP32VcKH35IvNfPxHoAJV
uKILtdiD8CZ3Ofa9v6mgcMq8n3Woqk7xmcOhURHOzFPM6tzN7Xyj6YRAyuVBnzVMQUfUlWZ7+R9R
rNWAl2SRbQ3UGDVyRkIl7oBPPpB79aLNVvWcdWBlDiESSXoKJSy6Adx8uc+oAYTdgeKYzbjJrhIX
Bl2XTfaBMbBZP14QYpcFgZ45Jij1nIwjVz6rUcOZBzI4T61XE6W1zwYFn4XzYJKRQBOk3KaSdEuQ
r8yS52KPGuLUIU6Uh1B4GR4ansq9Xl7E4DYw2Rsqy0zPEXPxAo+1gpLYjg2fnpT9PytpSeIiMwZg
JZj+VZvPzf6HnbSQzJwb47UXkCi2XqBlJezxeKiTCsNiF3mZaOuX9cQhJrKfpU8ap0bBdrT94tJa
TPzqJPRL1/MTdCCeni3xRDv8lTGduJv17wY48cqXwfneeguWufOWKXIBaUY5MlDOTwpuwoo2sKr6
6cfhhFoosA38JZFhfBwA0n6B0/XqFqibq2xASvtfT7rY6fzyjIEsmLko6fJuaKU8yT7z5mat+nuR
8ACjtWRhPLP/IYHndX8ZZmFuZjoedgbILLNgU+V6TjqcAt73qzZI+SBncS95lq5+OeT8bRf8IGhj
FDt9KNle4OAF35ew0eeHWGETOWMKnKRzH6N58qi8X+cF1cUrneDxLKx9IF3h5tEbm2IPTNLGCJmU
qFWU8dEYqC4zsC87zEXI1kDHbj5OyEpa9rRVmZG/4UdGOFPsoBWOG5dAzArzXso6NRz3dx3l+hiB
7e06BMXV1cgP5ngSVmFOPGod7y/Ikk+ELZKqbSkf0WfifXdqKPnskQAsDU/74Zo2k1oALF2U8psf
SXFmzCyy7FX6iExUYItBBHqo2FNKf/j9Dh+tIta1g7/ud2iUgdTIY67Vq+yuXbRP1FyeEEl1saXW
KQLhU5yog7kfF9z3AfJT6hBi3s1/Uzss1Sjs3/Qfj3pYC5ms8FOgKHz6XzwfkbFuQJR5gTc47tTA
bhjKpbbH18ESWEPW7z6FXNRnlaYfGmLMim/E/HUn7WHyzDlgole7q5ezDjCDx1wjS/TJB7CBKS4f
iUn8HLcBmuo/f2XE4lkVT8cJU4lSbQJZzm+iFtLzE8kWcBLPl2BOO9F1DvfM0uIiLWD/FXdEc0XM
5T9ufLPu0BlgCMetQEMXTWZSTuT/qS2JCFMheAT8UYNEZP7j3zRir3FpAgxjlGbpbHbFsdnEETmD
iyTJGfNGYj8T5nmquGaqLkkM2on5qBxON/svnIOqupJ9MZD4gHt5f1RKMOtoIsrGSOU4U5gT4nqv
zliS/iuXl15TqtpHhZPOU/IVQGjFjNq5IlcguuzKCE8/10oiXWh4fIUmHWxAFPfjaGFNqOPAriFX
PJ2wHXI3mdKoj+rVVs+QN6IJN2XOqrc07goSHJuORkS2039x+6caFQSO/xN/4PHZqGhF400guOUA
1yQ9qRY/PwQ5mbFvgCvvaX2qA4jrCzI35CxZW36oj0E5bNsL0NlBYB8PDn4ZS6tRzf8VU6Mp1nKH
x+AxbKcNsYdAyh+0TA402LKkUw0+uCGOyd9BMrSWe55VTAwTUV32KsmRYbZL/H2l+0pGn5sdUseg
zEtoDd8yRVbxHI+N5Ss3DBXXoWfhNXr9K8Y/krqbft2bGsLQPS6RrAGYG2RfTWWNhxRpQnbTiRS/
ll7tfmExQRKuunDUtguyKmAnCt0sg7hyWKKkuse3DYM3v2TgWL8qSI5TQJeuGjgBYe9pLDJ/eYO0
g/OTpHExYTuf1aaJfZ3+QVvy+gvJi4FCSzQoqY1xjTpo23G7I+Vqee655kBcS44wUAH6omhTFe3d
R63lV2XDyUdgBWqSqkAtE6RxV4M/oHto6KM1FZu++K1DDlXsKRXG3/NAHxLaPvdjLjFHW7K2k7tw
tCo5atOOLUbcT0wTwtGETWikGq4tfeE2DDJt5NddVmW6IkbspsoumQ9RNbg6ZcSm4vlSKjrkbDpw
jeUDdThMAxS+DSs6cvPdTHi3bVLORsopcfvW+rXo0HQLVAdiWtVwOad6qCcevBnnnpHm9URubTUR
BFmunW/HN6Ckl755+5mhyQ30in6WooMciWKB+1XJO+3yUIue/OrhOb+NDXCadhelENGZOhk5Ugov
siyFjuYZzWTRnTqz5hoIhlSknmdZftuvTOkf4g1N8/D8f2t1lqqFLzSgrSu9pKy/s0OYLjT/FWtz
H63V9xRNG4ksTN3KuNJwmnCDvPscPucud0HE23KRewupKEBlvk26aD3bkb21VfHSakth7V2NTP/B
MXrAeeo/bJj+lV/IlhvoyWpSeJSPUW5n7BJBL66wzzZItyxNhalfZY5TFmF5O0FASD2XNt3wrk+b
sZibnrVE3LgxO9ZGuBmAII+tQpRivWO4ilv2rynYnVLAUR3G5kd05WPHvlNjC9hNt05fAdAtEHNW
oHKjyh8roLYawKD2BzSrwhuzHrXceHz40Xtp8Sh1YsLmTHELX2z9RjGy5bgp6yfH3EiKJmEuscY/
XFxm3YieUp94TF/AaC3xoeA8TsxIh8E9khKW+5zChuaBUomutaB1I3mzp1sk/7ixuCzyXT8oov7j
etV4cq7iF6iNWRdvTTQRPhnV2EH6du89VVTYHnIDn4VnTA/HzdeRGp29jin0v9CBeRyJocHubpEE
Ia+mMDHDeTlUqqwdGSRSCYmfTNmXcckNjFDffTvwsLzTQjmtzpIL5JM5OI1R9dG/CVztmZdJRbcR
OkSA0dbLDo4lszzfwsueunRLQ9VqKrj2ghy2KxTyCmHhKLK+xj3XsQLcV5wTHDMyjSLORqNC7DsN
FGHRdWFxnXo0gyg0Ao6FMz9+kLM1p/u6OEHvkYl1sIOEAkWps94norP2WwrZNLQX8YhLmmLcwZqZ
e7ZaFFbzxvuwgA/Jtmj0bEkNTv0SaNuTDsz14gC8CxE9IYn6K0OLU/C4DV6jU24sMl7CGsjWiFFs
GV6PjfAvO5jwqShkCEULNHXY5MP/t4FnCAcnGW/zvH6unQx0dbO0oF/c6bpcdSVX4wYnjDrONKx7
G1fpl9eL33SCLeDJbuM50EQ2+30BxyaR7HwxItRQ5cV/FTIOsxDG81N+nkZfc8ZmiMlvAAND8jlR
vZ4zp4XihtF3xKD1gyr7U3ZoBdBeRVHecaQk+vOH2kDF/5/7w+immBlrCHoZFnb2JeJNFD4=
`protect end_protected
