-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jb6cc8YoghPUiIE++wKn9L62YSgkD1dtzi1DVBe6dJS/cKMs04uxMIWVtCpzQueEW4UUsv1qcJEL
rKCkl1Vexzrk6YY5l2Sk2kzo2eZCQuG1jpKwfq/Oita+dToPuEFixpPAo2/kKfsTpo96K3r4JSm/
IMzL9afYb1OpnKtwT0v1c8CDioZ00oZ0CZg9Y1gdoCRhhOO74TLnS6eoHFFCb51bGwA5jHSU0/fk
qP0quI6oQ4XPU2gEpcP4nUy87R2bk5VyNdaEdZg5MyiThT3YaeTLyO2V7WmPV9DwOzBhwUKQTCVx
JBjqW8e+WeyS2YMfQDDb4EEmgS+fi/peTNHeTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4688)
`protect data_block
ygqNe5lVdtbE92V32t7tDLJJgKPNa3TYCqAI1fum+tmlTRyU0YldVNSH7TSgVRS6ou4DF6cs6yqv
MBZBtgDpsVmqcZyLnv3KtGQdbKcLNrMNaMc2Fu+5lMnALf05i1+y6coAK/Fm/MkbX2w2OoToGIXR
KFZ8S4s52R2ZRh2E4VTlWGsdsx+HbliT+cGshPOjl1v+/TuBwNnLMzrfv3U+bIrFjj8NZFXRBnsv
WDWzJ5/dOn3iAYDd8vgbYNasGU11PhAYoRfs7dS4lkUeaqGgqTLvDkxmzkiBsBFsakBad9CU1+G6
GzovPvnCFUxA3diErX6qFzInEG3Go/x8K4GlKptB7n2DsT4VszCaHz0kn32JIZ4MMK41P1bPqkr1
+rL8ba4uHJmJvFVzpTID0ojFhSaswtaUiMmelKAHWKAgZjlQJ79FQSDCIkVXwXMzoeHephNYxloK
ANoOogtPECyve+kv3Zpg0Hgp9KG36T/5Zv01PBqAqYdYo4fD/qIsn0Wl2yTvuNy9vjWGJVu9A5Xu
jRmdelzLaJU7+0bm27yajT3fYjmKPWpXmImo4dRtvEJ8fCO9JN23AsnrEMAMVaclz1LNq4zvTGqa
3Af03ZwI3q/qY6l16fucBqy/Ygt4+0XIjvhuKym2gL7fwQyySNpl4kJQnQ27YsJmtjfv4BNakUTN
OhrzUXpJGalKed9baAKLwGVOBh02I4qfaa7iahbHmDsUjU34u7GhCknzlyQ3QFzd5mTeqHccYeFU
4Q8DIZcwPIBygTs2StY6JNHo0vL4Gx/X4mP9q2c/sDlR7dgP19aO4iPENsB1FZ2HdpPD+Np0QJHa
1rR+AE0H8xT7aNXWg8f0TiQWfS6Ty7X8ScygN/jl61jmZnIVCbwgxBGt0OGDuDqCARD2+GraG9GV
QCV1hmB9jglDVT5gg0+aiqtQUU9WtG0zScRnxtc2dT6s6eFAXqsfx9+S6dgxtB29x/sogi76WrZE
N2lFVur+k1s5cUJcab0diynSc1d/XXNpzwfz2lbL41O4DfFSSf5ses604rhYGsP1p0TZ4S4gyVNv
JJQzDpVwdbcJJA9A+sRUs5MTO4dhlUhFM0L/etpxOzahKZaCTFWy8opfLiGJsF1I8bDzFRt2AkMq
R/b8bk3rgbBxDMZfRxZJH+NFw41bHfgGdZwLutXoqswwvzpCc+HddNJMT3AQpwY+fMZmIfugpQoi
7GXRwIVN8I+9zJxykVNDfxWHTiO9Xn4eQcGdtJD0ZY33VTqrrNxd32EYtllULE32g5eMfWmkweC7
MijDVVajHfw9mFNfO0bylmcmRHV3LsPAe3167nRQidDmzvXPD7EwlXTfsWVaFTchdOgJtar0e4Dx
wtE9IFJZQkZVeiiLyYubyzvZgPU31DeTWyjwKLEADmIuGTPtGa42Do+mi2mserPZGnCOwpL8xsF/
+ZPH6VNpqiHyuz85vtHwzN93oTkssOAc5nSEmtsRtt8kSQa2ASKTSHDMe6LGY5P3y2+7pk1oLm2X
L+0Bua1koHjo9+4OjW1c4LMeHfkYgZgNoQqaOD2uFgQgXtLCBHhmLIWWOGzxcrtOaRKWrX7ztgKo
iSSonOdzbzkhxcGjQ6ewJaz4xNgzlwGGKFhU7mxnSHww3A8W3XPshksDJy1T+uhAYfaA+hLb5SVq
rVvvXVw+CW9DlguqQea+OUGwXyYj+0kOMld86QQUzWMBpvMCfBoYq8LqJ7gOiCdVl/bAZTtTiAhQ
9gpFEI65+CE/sJyNDf0Fu3TdPZYcCQOptFgGgxEnbGG9ZUs/9nq74SLKfPTNZn5iyjvZFtxJvnjI
qjcUI3MabiUi0Ph0eumhQB0JtdjFFJ32r32qNtxFVkaP/2iWCToUtsk96W68k0rORa9nmOFlkI6h
+G6Yka+3m0kv/4BnQ2bzmpCFSv1GqsL5e94dOuul/59MTD74ujPvKhqX+a5Ovr1EwA+/tGG12wCB
gAjcLcSuqhd16d44EmXMxxWYuNXe+N4+UZlf59tUbzVw0nrdQfSW3vKVA4YIV00gDs9i+UJnofFd
LbILDcwg7+aPXvEGbVbgWiFr171LplITxDxnnrexo0SfMTn4mgFwrCHhBMo1jwFcOVmAnZxoKjLd
30lm1CF01KgQLWJnWXcUl16d7BE2V0WDDm/Hha/F8RdLAoKlU3vD5sZ8HcCVplc1ooaKSTpQElYS
sqBAS+FnISRyHai3IU/LA4QVQAAM/DjSoJxVSaZlJNI3oqu7OtRRcmBKUYjYtajUtOBODQEuJd+Z
N5zD3v0RrIP7KI2TSwerPITh65PdAxGPDacLNfwc31JPg2w+krix+URbHHMCckBaj3ih3LwL6lUQ
67jFqacL+xf1NoJSCKo8UZ2lkR1RGLM2QzQC437wVsnOwidnxrE3pRore3mqUo8SZbfZu1gETCNd
r5jel8VXeQ1V/n+34FESt+aJdKJ+l+JaBcq0ybIyCB9yUW93IS8DqtPm66sCbRrZQmq8d/7Tiwj/
/fOgNAikUybvHM00bP7a9eJO63psp6/uW2qCvjhqYLqQgyyjpn1CHCEpwIbJH+k6I0ArF6lb15lM
f0UDnqLxriXEWgkqp9sAQOOpL0vccGjokwNGwEScUwNtaXZDw+6SiRMVzust49A0Lx89RH0d64FB
ePycIY9TlfO8RaH6TDpO4QX4xhaa3ga4y+pwgLqaFM7gnmtmxv1ZPVlzC6A76dnB+YTOGIhdJayM
4zYFkvFFG5gDYLx1kE6udVHzkFD73Mvt5fAM3IqLPevDzHSxw98/GQyaBUyK3PmBySnc2RzCVjwq
uFfWfC7U4ehXx8ge2Fa3wG4FN2S+S1Xkjv3hTqVBpRwfnMelDpfBn9WpCSdmNl01lbngwXAO3M3v
ymZC04rN3zbbsm2x5grdABI4gD4luX37Dx6f9s7QW6ENRUCpuHAxLddkdDWCagd3UEAPRIZHcEl8
3JvfxlYCulw9a56GMgIEHQY9gTKAEBYSef2th7aFZSyIlzy+U4lC4NWULK6m5mxrL1D5nt/BRgIB
5PiFAh3WlhLy9BaVgsRTbCkOPG1McPrKx109mTyDn8ZOpRixdESJKlca3dt8hIslszsYZbhzCosU
LjhyPFeRjiiBRYgjQZ3TWE/1RWvRbQXgpNkIASG/MRfuX5VOjBvNBI9DgvMOPA6Qn/LzfDa2DbTJ
R/mlhR+efsyGzNkxMxMyWRP/InW51f1Mdy2nF2nFWDYQP1opPePJtUjWLKNEeRVYhweuybLvklIo
yV1Q8RSWRUaG0Puqk0d2EAeBSsZQXQvvaJqQZ3prQVxKEhE6C00XGniWnTRxHbBJtkzSV0NzFspg
MQEd0qQ4inR6rYs8CXBjaaWRXN+9QllVWC/O/zoQyyxvGAmzKUwOkR8pe/LvSk7u+SUCIubGkC7x
IM7JZknEBG+FfxZ3xgz1S9xKkduhRAmB22tNeF10tvWbd1lvuH2KejPo4T8Un2PrsZzBg2dh94Km
w7/CqIkPh8ah1cO06S6mVNe3G8MlQwwzpvg+cAn5G5ks3b+lpuWbhkNl5gmT+1U+FT1icz/Prx6D
Mmp1zz6EUk+0tGRD2uclDzaiJB0tmjO7m+JkaPBmEA9EZ/evnfymZhQxOjA1UnzSNH0eUW82DBR9
uH+5WDIWdLtay43GMUf/zYyDPexdZlMen3lAYI7L+idFGn4pQro9WwGx+DNtY9Ze9JOZcuET2i7s
6FvarWR054F55RDbqGilExm5wWQYY4E2pBajraRqnqXlW54+kCPXLceDC0JfDRZ/YjiTo4p3f+KP
TDY+4ikTNjj7Cbwu76wmxjfohVF1Qre3vO7K7Li7XDGuZflSPtnBscE5pB/s4M49sHXd68NCfmuD
ttQ37r6A2QTj4cb84Ms5Ws6BLl52PRspV4iBBx7sla3YbA/PiXA4FFpBvcdobrST/SOfgbewy/NQ
EjzAEGv6Lu06Xv24c++wCut/MUpT46/uh+pTyqfQPAB7XNG7cj3cbqJdwqKl4FSlHsraJdbbU3lc
0xaB+oHpPcnvzCqLCq9kjAKudnl8rsH7+sy2+ATaaDGqRoL1/KAxpz/UukDdthpIIsqN7bGdlZX6
hUhrTj8S/OD//sIwJTG2NeBJWb/UnlOv2lbnykDqtJt9zFhJIpLthdkdWCKt4qkLk1ft/ztBUFLu
RgCWwJaQanC4vCzb9CUC8oo8LAdvxfJNSTMh9rOg2I1Y8swAXJyfu1GcFzbNQljmzUDU4N8Vmk7s
za7lxV4FOilkyckPOg/Q6W7+WABIzxTvpXwfePt4XXs9NpMO6PhETfi4Y86WpagO8hyUzibVWgzD
1mZqeN68aSXm7UtgMDhDt8d0sfmhgqv0ysAjbqqi5LzgGS7tfXixXA4oG2Mj+yUjYzGsuffngInL
5VPbA+pIKnwGTT00qa8cB138VcD69QkpG6gcR70xznhYW7KK0pGijXaqLg29MJ5sfIVTi5mdz/J4
Pf1361d8tj4UzrFge49uJpegJ2+gMCbbajXVgquNZ6ERCimAbWjsEBsyVm542QVpklMGLsKWUvIa
l7ojt5LNoaB2Owqw5AOrk/d+0cpXkmi1ikdTQYDlwMI8jtE+szjjv2txchor4lXyeGpvGeEuVjqv
GBdHX1NlHzeOtPMzvEiqOCMGsItVEr2rCVVvLe+L9Zrwis79WdlSqxpIBzD4afj32sQ0ZeXqpdO1
vdWOf6pNdiSn0OSNCwWrB4nA402mO7WPiJLLCWJYcd4hQUruFz3iy541YR0OGL4hBP0JVUYiRCou
mhe/20MvBz38GUIzfm7DYgAIvKOhpoEFMMXcSvFYCXsKHzGs1/QiFORA5EmXDVT7yWDYEInJT1Nl
iPBsmELvArSXrwdUdd6tZmwtsgQAi0wIG++tvrUf3/nDfClExhJCjx5SWm8rx5rsdkToOWvnAUV/
LLhZhPP/b7zNfBam1o5RDvRiko5LFSRskpc89V8haAqTAF3o9ubBqmJcoCQcEwqdrsrLZ8fOFqWs
E1Gx16Yg5EWW245KfojColk61hI7HrQjg5GOCx/KmkT/LfJLN4TUx7LkeOLbPjGZW1pZH48KhhZN
bQpyRk4tKkxP/pSvPXwg6PG4PRBy1DMCL9AkYRSqqiVWoAd+CL7FFEz4sRD0uDt430GNuShAiMUX
Lyjwj172aUCq+guuB6oXZKoi5Yys4SXj2tBFrbuthdhlh+XDQpRW+TGsjFhaLCP+AGwdKGaBhcKD
b6B91FLCJqRKPTJ5Jg+fn4rkFoxxf7G6i8YDilPxrkczw0O5G8cKuQnbjzjoq2ceLp7RD/NwGOLV
WkU+JiE/nJSrIHMXSpTQ0eCFPf+V7/tCZkwftzEiD4fCQu5zucGlftYs2dXije8pE3kwDMcmdNYn
5oby5pd/kmywPToqaf7ljuRPCkIl8Wqn/RjA8teGep/h59VaIIpexSsdyApknI027jOETRDMdiaF
7nusYAoeN9TnIzu7fR72TM6ADLCvk//iNOHkVhothUEAhn8QIDjnk2BYOxqdbdNRSixLPeSy8TJS
7D9Mqda/oPumJ2fU+wtkYzkrnUE4VmnCEK7NkryX4b2VHqGvUbzfVJrwclobdmAE8WbjwXpxjZDu
K6F4iVmxN+buNM7onWy9QFJ88jfE896pGNELro+R+R7ZrOGYOzpSL/PgFCxxE5m/+3H4WTQBLlyI
qplfiFmzItr3/DrerJ/c+dVLIJX8L0vC93WcTvbMcbRSGrlpAcqJVY5IchHpBrCVIfu+1Gca3s31
P0G43g2a9k0/koVvR2zCdF9pTnrUKEI1KeA+JeXg9SAeCiu8rCM5EY24xBtzE4julZNqgXiwbPOZ
Sysd+wHhg2wdyawDcSm/r5PZnDwLB8/ZU69bpmzqu/L3/7F304IfG49+wjLusfk03OpHdwfZJvXQ
gJnDM6Dgs7D9dDVNpzJczVlmdKjzlUCkiyhNWvaziTiVh3Xa0159EH8nH72CSJlSpC2l/7dhs23E
jcZRGVlmgeS8U+CEBqphOJ8LL//w6L8G1yZFpTW/ZWPAZINhmgQJAIa2GMLfjpishzJPrUQ5uM/y
4VICMUShCfD62ThlGizQe0rtw+RWFKWu6KTn1H2zwWqMbVO8QWYNXENZ9hkZ6LLCpS5JqMfj9OjG
HNi/Onn0ZmsiAD0SCRmT3IvaIeEnpv9ZO3IXAfRI6VlsMgfxnpzIiyKH7rPnAOKPhRpa41uIy7uA
RVfopSS7/oEOuGh0UjE=
`protect end_protected
