-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sM+Zpd9iWd+FkYFnZGmiIPvefpNZVbNCEiBct7sQsn8vLhVT4MpEByi38YNGmdJht7AUEmR6MlUi
KGbNeK0apOgIms8sLml1J6wj2xsQo/ZIG23rxj4iTROpAtFxt9wz8hmMdsKCTMA/ExWjq7bEvqEL
27ZjduiPWRzemNDLr1gqlzW8m4lK98rwz3i0VmyLbYZL8sZtIMaj9kEMzL/EswrHR6Bt7dNe3FDs
3MrbHUnIQCq6mSnzaoLZGzZQrUME1LxE95sQGDcCtSbErlAxFkrDOPmX7rvsr772I7n/j/ksZtVh
b5GsPcvNoKQ/8b3Jtvk1ZKv2b9izv7Vrql/Lpg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
ZbqVJ4MArnzhsoLXg2M/V+X03GAnIyvGQViZ8OLymc+wE2pplI7vVgv9UbpeaEKkbQ2VJd79tx6o
EgAp89i1xdDdSqgNPAOwwNyL2a8JbPfzEgi5dQmMWepfDSK9eLkvxGNuX/dFrZAnhhySwCg284Sv
GxP8i093iWrZ5AihyUpY99pv50lenYwULNvcm31kT96P7pdNALybvT2XC55XBeQhnz9/vuyhiumj
J/T+yYpihZlSLP9NUqZe1tMBRZY91NPpPVOm0nUH9kWY2K+7t1J7R5oQI9+BrIs2zfhgpR1K8+GA
KU1Ngs74ZECuQizHCxucwIXdJKGiKUVCgA9lPAybHjTC0dBRJSPX3bcwlEMmWx4pFgjU36W3dzQg
JSFQLz4FfoVoFmiM7eA0/FDUQAFAzJDYjBgjtSBytH1keRcJO9EimsR6r3ucaulS7kYf4WScRZmY
JzS7XCEQfNqHxuSBEAFkN/vSLXIzmEXQBoWFKMa2Rhjb4FsePC279QH3V0Jf2JCH+p1wTMsPkd1z
vjERooBj81cjxJc0irZEc1XtjFqyUt90GqHw8tYQ7FK8G1hZO5uIrlKbH4BBNQ5OD584Z7b/RQjR
iiZd02bC+v/DLKkMWUz3Q/3Zhbqb2v8eBbwQRGqyX5fW4w9tpKiGjrBKWbrJ8bXwXXxslsJ5Gz1X
CUV90+SRfh3JnRQMFVRdAZi1iiVLAeNJkn+p4wGCUJAn/VUxOfNfpRKu1uwPFuQguPH8Wsdyx5Pw
o5iG+HGyr9Gebbc8lzC6KE8o46+VvR9tQH7TrcyQLnPpIopRkG8ig+b7JYsG3RwEJYRXmfMDkMbU
ryqXfnqJBe388lj68XY1DPUCOp9Z7SnXmQYG7I3lu6Ki0eiUOywllfe9/XAffVU1jnEU6xGfmF9h
RIE7aNBOnbwDY4iuh4jP09Dek3hD/0VEXWrR7UzoJ4MAEBm13G7ZD1ptwxhxoR3AI2YXlyT/DA6L
r4ETVlil/S87SWdAgsYnpKXAocMpZnEzXMgDYmycbW+14tYAMG5BTdSVl7uzuyY1eH+RkraNh3/q
XekdIkHgIosI/dz//N5tG4/gKCMZv+ZJObzC6BvpM2fzot6IddS2a8yItDSyQEY4INIuHAU6G/bG
Z3dP39p4YDrWrsXQjNjsIKwzmpKf1gf8FVdO54V62xIeXoeuo8d5QNE9tc4Z5wKvULAGvRV1zd9Z
uuFWCwQ+GtqcKPXbfRjEQzwnmiVR3+JqPxyDOzi87t4K9t1N2j0PSs/LVwbp1DttYFaABsrGmNJ0
jHgwSkuXza7j/I/wHHVaCog2hltHewcXDoJvhlkoncC5xL8PMohG6Kj65GpFdsCgNhqsqZQB3dh4
/CvY7IBRLdmyCiWi7/xOe2O6SlsKGJpcnVP3ttUwrFPviRu4FGXIoCwu1eelZs2CzC+H5KhwTAvF
hkVouabnRN6RIpJCFXXlYh4poADpchIhy8RmT0MFhwvP/49ayd53SisRGNZLszUIOeAcw0F8jP5i
uOJirNmLVdPiRXaLgW/cY4Z+XrRwvucHxflrduRbPGT8QCiPC7cn/jqGY27sdfGzg9X3xmDtQ7EP
Dn+3YSRtt9WSTkodA5qPda12NYinDbS+7vyN4mQo/fy+KI4YSe/3cmHkcf9+3cbU68OXreHbZytx
NPDB2MyOeqBsfh3it+P5V4YL5YJzbOSXWFLYRt+MLMZ43RTZIp3nT/f/rS9iyp4XUOu+FfRtv0QB
UhVCn0rOlHKV55skL+h2hDrAzWF8v6k24YkjopyRPKrTWrNAUqAjkJC+KUYElh1+u+AAgr+Ka15Z
yN57uMDG+O2Q0VfiOdJ7bYZqcyPUfk7CLB3vwVfG8DJckMf7FqK/11Igt22emdq4jVEqZjz8m67C
hP8bQEyPe4Xin8PO8auZSzXpFoRFsSS9V+GVtIYwWQfaGNkqNcse+6zuqVphVkmZcDtteoIxGaLb
6WikP48/XzYIaXTuvBw6bQsy5eZyY5jMLQXYER42Uh1wx/LZ3OhePIP7FstMPHycgIJ8tO8OSrgG
v9YoFhCwkY4EepKcxb2rV293L2ERCLLWJkGZKl+r0Ij6rWIIKzXkAaYIGFVy4fI2U8ElgWf4YqMu
axkd/fdsjYsNcdXyGmSei7nvNZKdytz72B+ojVGESv3lfqVdTrONG9rKHiVAdvoZZHDGUibW13Iv
30X45/oRmJVtTJZ1KWmGsW0TPd78ICJyDrVUiXtG6DthBGs0ZPMz0uWkbCId2XkRoCctdl24tmVu
zv+oJl4qTVUpyh0Qm4pjZfiwUEIyYAzN0ehc4k8hEowtbnjskvkKRMxF1yMzn+s0TFKf4LfSaFYJ
MpMrEeQSp6KIYqE1yKHlpO1gM12idawqs2ltYozb+NiDic9bfDaZYKjDxLyNNXXJF3bkXp4YROd9
uda9d6IyKkeOMDCkizOH8/+l+8DZ68RmdS92BlV3NjrPoyD9OUQu2LqkvHwL6ZVZjPTcjU3+ioUp
uSugTiYzI2p5ij0oNq2/0V2/SnB2wm8BC9XAuNJ9RhxjUfiohDFfeAgXcAQ7Z7e3G6DNwU07xXea
+GCs9+XAr44ydzQ9Mj9VLujFDEY447vypa8I1FNomN18pHHV9FEorUDM3goMnuTiwj6x6Ojv1+sT
ZQ/RR2krTQR6nibvphQBsnEM0jzKM9x4KdL+cuqNF4w8hOglt3dtUkQhSX8AqzEm2scQ0ndkSbD/
zk37cI0xgn7nX/QGcMbCo1i4EjxRREBFUNg4Bv97irMfTkzskOckBnKsJJL2luJrpvmh4TeQK1OJ
L7aXjBfwzLsQiGZHgdYfdxObt123+wpxNj5M6c2/OnCG3tVhl+Qw+Fzj89Wvkrtj8fPpCtGOf6KK
u/GPb3/igDkET9l3/GEp9QQQotHrRi7NOTLsj5uDVvpJt2J3gRh/VPI226gPi6cf5WZmKeN7YYp7
sxseYeY50NCCq8DX61fFcDoz49v21n5+haMQMp4mgsQgBqJh22fXav46DQ6U+c3q/vsc9+j3Czte
Ou8psfls3CeEIxkefdO13MooLMft5Y/S2DwcCaEmGsKgifGL5qimVac1uDKWO8SdkxrgcYhcWoiq
6svarnNbgBKX1SypjjH5/XmouztLQB9AMPDnZOisSICYtBztH6fH0fw7gOSGBSueiHMcfS9d2QUF
ERicVscLsdF4htpthvJReE8jfoOMkmEmHOGoTpQf5bXOz/+duNvYIkPBbcvKpg/b0ylaInUuyTRc
CBIN0wSIak/QAJQ1kE7LnVRAioTUD1uJTTczJ6g3eevtSnBCk7Ib0LfBCm9MMr3TcFd2iCBsZ9L/
JTvvWMKBkZ5Mjv/wrNrFQeuFBHSmdP5hvuLdVSVZ3cHxRwekR+WisNYhQ4FCZkoAxjki8PdOZ9bm
lXMJ+NpZsj15kNPpdbuCXEhg3tqZCd57LKQyi9NurYcC+S0Rlv0huA1rskK/MUSSPbBRTwKYEYgP
Mvzik4QmD7lxSZN5+EWizbOLkilmCCQvgWzxmKJEup7qNT7t+ZKXC85+tlaHTZYW2JzikAeLf9MV
pi0HieWniOtHrbQz+qpFFLzhiB4i4Ql6gBRW4MulJFlPNVDnmBbpzg+yL5bo1TyppMyCTTvGQ58R
JIiIIsTVbFm2ZoInvQnzuSF6q7HysS4xVLyX/DlIgffZqi+KYuSk87RQxuxUeHD91xKXM9Y40iFN
yKK/7zyQ1jthBOBfiqxJIxI47kBY1aE87jtCnhniR8frkedTBL2vAwgOu++ZzvdIafyL+ILcUIU/
aIGfDB4tVjD5jmEUTpY6lDAoG1EkxwroTm7X3Yt7Hmxio4O9qrFCOlQVN/t1qgY+mSfIGWhi4Alf
+Kb+K9oevUCyuDMxH3o4tsNCI2hYaKP74sVDEG2eiCRfaGcmxKIIDgozqK4zxx6uZGQ0iDT3/MQ6
mwF7k53bEnW45tgDNAbPwdX7bV3laNL/31i/bnoj7l5LZRbcAjNALQes/oNfWWLipHQr4IxCJnFV
eaNHZsijIpQRX5jgsxnbnaPBGqmMSraMfcUuf8KBFWTaV5DLIzqIW4TVaimLQiVsMVXuvC6snZ8p
bJsDbieuhV0Fvo+g9uQZCHReEldWgBwcmUh/zj3wazagVIfvK/2I2vuPky9DmIpu+l0dNNN+L0Qs
yAjNeoF1uxFLVcwhDjf9cvIYKsO9MKhBMqBz70E7DhOy8QR+Xo0lg4o02TI8flTpg/IhPggh4Tq8
clxm33A5d5J9yvTiG7hMaVMSdNHfqasWipthIov3REGMQZmG6B1RksOr9x89Yi5t1MVy0hhn1ssB
qCKI5UKzufI5ad2zFUS0mg7DtxhuPRXPXYAC/P6X+ARShyVh5tPHljYhNSXmzWZ/hVxFJNb5zIgs
KPAU6HPERDs4s3JP1orNwFJfnI+uRATdPL9vWoDwSnA+ndQS8bfj0p96XOIpv49oBxmMqT0Ug2Y8
5SKkT5s9ZwR4OMJu11MWbx43LBKXGDD+Z9rk1NIuy3QVjpW4LNObI0xvF+K6F5MwTVgJHd0gWOvI
vSQmCz8cHVbSgqwtCEpmFUWidLe/MbdzpgYJ75c2G67WcumsjpbPnvbYstJZvwQCmRi2c9xOFpfl
WFazZL39JmXM1n3BZ8K9j/j+MkxOkzM9TqZNSo7/P1NG+5t89icu+1kBWyr9t21mqiUXajVOPx7q
1sRCBQ2gigzZBf+arLbT8txEFdZS6W25f7WLgMkovq4Ft3ANNmygaylmxDDC7wdIiBm3Yt8KXOkd
8nvEwsZw/2qZ2g2/bKgml6V1Pp9u2EfsuS6+iLfwtwFu03Km6R0Y2kkZcspswfDsSQpbHu6Avoe1
Rt/PSqifcF6ql8DTBLtUfkzKCErNy8+Z51Ojwo2Z8cD58D3WhcidlDu9XjTFjXS05yllOmdUXsCT
fIsOyydHuQK4ZxltzV0wvOtw/wetQmZJ3+840tT+AsLWD5qgV6ipKHFMh0O5RgOhpYFs3+ckQOgS
RbzWtc29lNLqUWg8UV9SRWL9x7ODDRih5IgbgZXqp7SFEjVV0S7ArKXqJRNAaQqZjYZbA0WWouWS
xlML/RRuTmF+smRroMSLaeCUDeVB98Ou4eCdDlpB564tVRv7N+iHUnL+NQaD0nJMk0JrSeXdF5iz
11fjXMZzJAd7nSv6cDeWKmcykHG03wJ/quhLOErUoKifKJEIsebD5kuB/M24yP5095uOvcz0Vdx7
5noh2w/vktE9LCD4Bgp1oLW2oYo88oliAW1pfq37cTnjX4j5id0YGPb5Hixz1K4M3HObjNtpVwXg
iSnzQ/BqXgoRlt/ZlexgGuCUjhcA/N3IkZoQU7YpSNd9tcDUh0aKbOiIV+fUluBU0ecvbFEfH5ws
mKvp/bSbvRWsB/lr/IYDv8ZCnJ4D8J0kbFVQDc8R6Tk5D8h8oAHtBq4AeYYHYqgb2sPchKsmpKtm
ZwhMpjzpbMeYGQlh3rWn4Bktgk4iprjczt67ygb5bcXAoLHrzaJiCvmv8RItC/vm6bA9seCnQJ6J
MOINd3Ua8KgsjTI9fKmIN1xDdJtYIyHwaD+Ku7V4O36AVLn2Y2vVNHO1f6n98eXdMDqxGnuTPPq1
1OL7CflxuBy8LtsKOAIriUeZCv5GrjTjVzxltVPggSfJL78ffPcvwpnA4m3ZxbNrPLceQGH1onjK
f9DP5LzuToqgxHgEB46zvmrVaBmgYKPwBFRPw9ZisoC05FJ3mUVn0d1w8k811yXGSHBxyOhW6IdS
ZyR1pfx5vRv+CwB876t4jM5/IAIdiONVAuh4BF2G/Tu8uYujulqstuG2F9ZyixPan47FbH57/YIj
XizLfz8DdPrrWPT//y4p7fXLRi6B4rcNTtLoI3FmNeo4VmPGIMQsHBMp0qmHRSzPyedNYrRjT0me
B9ZcV/BR6iu3UCdRkOTjE+7QT67hJ5mS0NQCxJn5TXLOOfR43PGDGMoNsRISLuRylL3SBz1FKL6U
6qmVEB5T84SNEoVm9+ejFnRZGVOJn6dD+xsxL6mMu4aAi8NTGJE4SMg29UTLF6uSB29n9m6q3ByW
nlSrscvhVn23gWb+VPj7gut9yXNpuHZsFR56m6YoHkBaENE2TR9O5zWx1SVKLNLwv9vG6KZQPyH3
TAMaR8zbS7TBUdLOjewR6HOPIYmXt3Hz2S8dJZf4M1GBD9OSecuIqKEcHzgdYbsUiViEKGpWgEMd
obBb5kuCo+vjrasQeja5EKJ4cC6toxq8CabsDXVAK7MYwG+evNaQq1uGyGx44xiFoK8getZyxaAB
2yUYT58erWMpVBWzru0YpKegqSpKOxOYPHsiOW6tiOz6h4V5go7KoS8Tf4cucjyKdL4SD9grh9iy
zrDSPr7VjR5q+yAysIGlrPy3QUpp9zYNL4oH78uH29G+LT4mYLMl7qIZ18OU+5derGDFla6aB8r/
y8RzZrl/VCxMHD3YvGURjqfBiVudJdTreu3ZbazoxwkHL3Mq87pybQjY3+BBU6olvQVo7Nooq0ia
6aB3b+aA1CozpKXU0DiT/sevGpfrzyTx664zAunEYd4q9izqFWzCjnaX2ZRICm9xTvcZo4+oKznS
gptFOTztpPZeYy2SWVLbRW5LTq1Ryn8q9s53qX09xmkGSIPUjd0hvJWQAJ0QaLoXaukG8kJTPlRp
wZslWei+rGtb09VcR/xSllSJPLdU31kIrycxcqzkUIXsz7ZX8JF9jnLItNJWNsFSXefmH5toeabJ
Dhq73zrj+LcwlZV8+T0PKKOEmPWiWn/nFcS3vG3zjDkRF6Ju+n++HZRuq3Z/bE0GVX9DXQgl88SG
Odj9fpSdtVRBmubW5V9mKV4zTs5j2QwFy61Ytll71xWXEwMMH6cslXbLhC14gB6nTGkAAjkkjxy2
91fy0RZBl8uA9RdNjVVohxd/WdDhSUTj8q4xR17Yc8rgdA8IMK/+DgBL4zZ5NvrzIZxxAa4Rb0wA
vdNMuyFGzJ4Q5W3MpGmbtUnLomkQmhmsD6e05WTMeZGMfxZrEftQTmLQEzav1RzmKol8dVeHxYT4
yuG+oPRVMl8dh6ZwvZH98UUdxyup9jHL3fiZppGUzwX8x1ZexgrPyM5/FO47bNgCJBInv/SpMrgX
kx+oh2ly/Yx8gYpTLrnIvS9FRkNOBvP3aj/vkEQ17ALWTvgC7y6Cjoq4YGsh3GsYG/88lkHDdoqP
XsQ7/9wbmIXYnDJD1Ml1na7kNoGdmPoCKtix1y8s29ZXqryARkTA3gsuN1KSDJKH7XxlkjPQThRD
aevEK2zjiZTIGCfFtCwFMKAD1CyDMwdERVoqRqyUR4Hi//gXDutj+oHZxh7kOnrK9fQBBB1baegU
tt822SEnjZck+VtAQagraGbM0E6WzvRVEUSSHStBM5MvuqtXIMbZedtBOQmAmoyUwG/F1qFhQvzk
W0GE9xRAT9kmw6DzxnSAxH8FU6Ow0kJoawowwpnpMr+BBgSobGpfn4govoWcQcl4gCv8U4FIbfT5
GFZhzqAsQjVcpYQOZetp7n2foLNrEVGs7ODhSDYHeeqrGbwYK42HHBCkJiAHb0v7MslJd0fMCFAG
Ecd3poSOsU3zPrYezRrBbcg0CZtRuVeU2hvquLpCIvt3Ej1Z9L8i14KXwTfGbgQUbAwyymW2tNCD
q33AjrGvGYTCwS8b3MuocfOo0DMb0ktr0/iEnfNSTmaoqOxm6kw0poAj1EmtlHC7SU1h4poZ8tM1
d06d8TyDhFdTLwT4E/zIbAvd6/GBO3x9GxmugZNOD6hnc54HJ7kdKbDIYS08RJfx83wdy6iM3ssM
Y9pPpgM+egobmbcr/aYgudDvy6fuc3v//PnFkAhZ+4ydRY01MXotYE74wxHTaHH/94vNPbesz2gR
QoCXuw1ovSV1Py5v5Bdjjce6YSnfhr2OMLN1AcnatqB1JDPUQw1F6n9HrvqR++7H7rEfCt9zIkci
PlDFykGTAHi+ctkB23yPBjJbdvHUDAbJ4ntPR81z861agOFJcsy/w/+zmsPtdDp/hahCUSg/fc2B
Bs/3Y2tgZwfNST709392fsKJ/U2XItL7ngUrmRB97KHEcf/BmJh4K5CwJfB9KeWGf25cp6sVtac2
HTlSneNzBXgrxp5yK3+O24lPuVZZre8fSrwovgWAc6ZxDWOLuq+dcQNcYLpLo8JEcuqdSTF734hI
Qygb310YRwpz6vqrQxj8fGPB5CrXb6x0glosNrryLFredEQ4CPdO1jNdmyjGvZo3NXP1HVS0wlrV
ElX69aCa2l56au1jGIBMo2QrjIsFZjhOibpGIGXzjNA+QSjLUUsxS18/3bW5qbAghUHkcijGZaFi
KZP2r9iKp70pRmJybHT+bjyXmKtbgXkLLwMgne3oJfjzn1fmCn+Fqlnvurb4vrRsjdAjmRuFUKwT
4k1zHkpYxk91wv18j3bqgH+L38X6e/BHgJAorX549jLw3MZ/spUJKoE1VwBkqo9jBfPK7UuKCwxP
3tJ/UOk9yKRVvZosLzUKvRWxiFS5AuDNPCxEUpQzFI3CaWbnxrsZxqqfoG4uaXYrpoT8LdR7gcgz
EOs1qrapCyXE1zn4b1xEerR2keldpi3XGFdaUbgDiXcefzE5+eZnY3aD+cmtSNt+a5bbHmo7dsQF
+rihWAnDCObj7sRSBqkyrQkUNHzYL0/67jZDMRK9LlkjQS/4KaV06+eb7ddzJf1/VPI60ia0BCCp
RTJPQFRh3n8xd5z/VyQT1i9aykXPZK3+O7gfFPWsaTV+elqkXKKejXn7nTwnAvEYFGEu6RA+Ijxk
ruIiwkVF14J9MykL3orhmuqh6tlTDg5VAIxdOzS2v8Wj3ABIIMi0WlUxshVFHmrs3dEl2xlctJU9
rOMqDx9zV8UgP7oMKPnnXWiwNi/f4p8UxdKdIfnVe0hxZEioZZJ9qUdzVv4V2jxKD+HtwGiKZNcA
NaDyZm8cs57bhSAJ25Ewp/ALn1FjiP/H5GheCFic94ASgP7mZM357BW1sIdHMjS7wphEQdlV8Ran
sdquAGQlsM4SlLrlOfxmSEAh7q8TSKe0qFjklTXas0Agb7on9ydoiRA/r0WHN8+KFWKxYp1sWDs7
/2pf7Kf6lw1YblFTbwoHRVVd6g8PmrL46YoNzhFCNuaoR2ynF4q6ki5etaUSLS/PHgOasLKZpdLT
hk6EsXHEqCtLaeCNP9axfKA1IHn5g7BCO0C9YNnkUqs1ixq2KWDsk7+xqgCyeHINaC54s+OEvj4d
NAbylj9Y8IYyBaBhxLD8DlkEi4bh/lg86I1iTT+Mh55Dl6V5n12WXM1W99CY/4XqlGSetefl33QC
1VmwrELKxmgOaoJ6fjeyhl6OfwWTcH28XU19m85bifwMjn/qyrknGc14B7aVwigYLhasM19bAf0M
jh84rHblEwO/n9tt9wbYVKfNda+bIx3tiz3gZXIrlLT5fHHfTPk2yztM2sS3pavM7peIwMp7Ds/F
JKu2cWdfRLnWUprWvlWJ14qn8ZWBUqiB0bfPT67kwyBVnpgr9vkvwiGTpGPJ0eqF8NrxyF/YW2X8
2C5YNq/dCnKg/9Dax87mbPhFOxeyKoWTV5jms4dW4EfmAqZHPZZRVrAZmh111kzzHArEJurPUGG5
omzSus/3FHd5NjIxbX1W6dPuZLECf0mpS/wFpDhsC7djC1z81nkA6KKIPGKk7WaihcGmmcwA+3gb
xDV01jjwYy10qpdDg5R8ScM3Guu3jwDi9vFo7l5N3kHBbM/ZGlaz+wW83lxY9d4zhbWAJ7hzfu4m
Hz4Ryx0ak+2y9H0o2N9qrgFtPDmWOzAipXWTIG/xtHja2Cq4QuJcq0Jkj+2H36rvt0S7MY6NCF9r
Vnxzd6QYMiJLmKLFySsaabaQQzWVCVGAIobRqUx7q7rp+cGFJlXsCsm6vuQ6nC0HF/wkmmG4odFo
0VymcrWmIPdYIofXmLn9/oaJZMUJK42x+K6n6KdLFHp/X5gghJAa9sOb2LQbcgEo8LzRsJWvvid2
1QF/EtSvvmxnVw9vZx2dqHh6cjPy2YqyFF/CZPPcIQUh4fo7+0vsZLKxQjQz85HbV5pWzCm02zTl
aa8ASsad30N3laC2/SWpe9bKDerOp7gxDtjWbQqW2JUcOjAGKwvuJPsGjhV/Ay7UZnUdZYFtXn36
cU6jaR/DJO0vgia75KkfUpH/70FOqWVcK+R+MMUu92FRJXioqYZH1z7yEe/sQhtK+of+GthEQ1Jm
ERhjPxKSoNDU+R5Fz9sOqMlSgnbJHdDOsR8lQb1E7HctyAilCAJNgH9UhfrO0q0NJ6H60imYQTSC
Bycwvlpmtd5/fVyZZcl7jxu2jhMv1xmME0fhMiy9qonSSjn8I1RiCKjSuG1FQT8NzcBFHYUFLZNl
qHaBVh0j9Lxd8RFYCbE2KlGPfstshS4Tx7wdP3/5lCS5lHvXyX520uIAAlmcFHQpo+qpUmIskQ5q
8/pWzDaRrqMkV6fflOO7LtHLDj2BX4pMj+266cc/IzaPvqhYpqpm9EPCcl44/hGXaV+bhMc8PYuP
oUYTK16xaEo8sDhh+LKVWukThovXe91LfNTW/RCmnn+leLIul28ZHc/Lis7ZvWDQ/PQXaNWmhI3Y
Y9z8uGL6MIQ4O8/dZNB82DlG3VsKGfldNIOkHASKUoIotq9UeK03HpedRgEScPUkHgqoIqhfk0OW
gWOTdFbo1g0PiH8XoQrSqm8HqazrXfpkaDZpWcdRUfv5dv0+LOhNqtXhcTDxNfTnptwRleyOxXnE
dsNBgB/7VbGnb05JHl2f/kVWMUW+mN7AaJ7pxxr41KH7K6Uo2CjnsWVGwtkBL8psEji6h9AGk9OY
6uX4lrBXoa7edHNwxIgmkhSK20Zh4gsdSX0Wp9G7/q+jzZhcmbWHJEYNmyDZBIj11kZykMFaV8uM
2P+lgnK1dcpPsM7BhEV5jDDBYdjob8JUMUhoNPautlpFTUUwUxhjG8SnefB3uMh2sWjQHYcobcfo
E7w61rxmbVFQDYlwt5b1RTz6panlS9z3qyByewqztDNuvgT8DVN2+9/Y4GfGhKe0VviZd1QfnTbw
bDLjj1cFeJ7cAVP3qT3E6rVEpXUFoewYxd9q6clk
`protect end_protected
