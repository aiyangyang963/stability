-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sYI6Fdq2T25nOEScigFMNAL0xs1/DcpxzM9SEZ/1ZPR7V52qBpDh1ASVMV5OVqib5UidIF2Kq4Te
UYChmmHXppWIOVtcJOoop6Z4ryh+rkjpeGLuj5fi++XQ8O4HpATZ+zouLoDwQymPGV/c9TLnNE09
zwqzfJT/BRE3Lk/OxOxmFawQjBAsev7oD69hmNVE0mL67lroT9Rt/C4cTKeDq5eqE61CVDV7wLbv
brkQZ2yMQin01hCY2juy07o7HW5C9HWuhpomgfg+XkkFBXHoBEZ56A9G+9D+3G+dhXj767PtxOQW
JCLaasrVPdFzSeqJGxsQh4kdbovB2FqgDBkYFg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
94TpAPFTDRQqquSRn+H20HP56wt2cHOWqKUPg0bMH4NC5QLPc4uOcw8uWwamvt4N8PljrLgwKR3h
pH3SZ8jeOngUIEMyziZ7l0O55KEMmcVghOn6P3v9/Nl4NBMTqFa2r99gLZnHa581XAYdvH2dfl0B
4XME/t+3LT4ZL4jlfuvwXJ+qhrLLExohQ0wdQVrrHxnS9G9h+jMNOQcThXsyysX/wOUj0QLzwpyC
DZdWh/uXlB7NnlDFplMyfIQzt/ZaUHRVwwNL6heHEGB3+udBdCm8uuyuRptwpZ/Dszicjsx4y92+
blSwzoTHjNBT5eg/ctiR/Rjkg9Nl+rtMuRE0VrkLaDWmqAlXcUisS4jnp9IOh+l87uVM/HzBfX8P
daaHqMDnepzBUaBmQYPbNNX88UqvbxryOyflY8issHYmbUDqn2/uNpnY6QxAZ5xAiizaNtma7HOY
u3VmSEvz4+yyulJKpJQX+Jqf7VsLiJe5qGeGRgN/GsApyjzFHugUeZep+3+EGrPISvQgV67ec7is
SBkv4SC0z6cG5kGhuFceTEb6ytzT2cW3tAuN7uPrjGKStC/3tH/uSmS8mZEt3BhNz5707nb5vDJ7
Fa6M2/mPVEvsxx1nvBkRM8yfmY6UnC9OgUvq36v3HwUj5aMOIzc216roPGxtqvPMLIbPbI77bDnu
09Gr2yCfgRGqbRVbAH5KHzIsqldiNr8g58mJHeGHeM0YPFvbS/VH2SXwitUtB/mo+lzMiJQoynmP
IyjCNcbN6pSoyis5QXdUYMyXCLsDpkJhSVO1SQKNtVGQoxPHRA4nc0Kn3eTI2Rrsn7TDuzOcBvxX
7s1wTREs5zl8OVFrhpx/oI6phyhbSdJXXquleAijR9WOBDT696C558AhdKc59UPcD4rf2D5DyLDP
bioMz1GHMHUiKJDEdR9ABgZX6gGV+FPVbw5p/Z6JlhCLrFwJ5R3rNCoNbPRtEmbdaYQHgeQtViYT
eCyqKKYHw5F5JhAQnXvOu28RPjYdupota6djwv/E1vKge82ymlNgrHrRo8u13/Z7MdTx/NGkT5/C
1aUq1ppjRVfoQfdh8JugLc1f7x1GxVnRWtqReaUSNuiiXzWFoceIxgrVRXmPGFc8xbwpZJkFzxpG
Mjn7gra/AhDVD9shwCs2frdBXKgw1kdB9FForeDUDPrzh1244gP2xfaO9rDw2XXp9jkjY9YTFUyQ
dspUD5PjTH1SDURsPJ/zovZdM8u/RC2766o6S+i6+bEH/w2IkujUeEBwNIXWNbmQ4dEYx/vBGgzQ
oEaxK8I69kvwBG95icUM4a3qKt3t9O+b8STG7QlJQW5opXFV4Dt6Q/HHVp7Dcw5oEq9GqljJuzs8
KVBrjKdhdJcsn/Rc4rzdMOlL4gTcraunky9GS/wAf5R/YwDwP4MS/9PnxGGnpRQOiym74AuytniL
Mw1KQka9bqLdR3mIY6AXIjXiRvYQ+qacOAs473Tl8FJzYJ2OE5B/r7YTtofKmY0jgblXsc5M0Awu
hCKEUfuVQ5EJghIoi0GlzkqHXNCw266JlOJVecjXGgPCIIrSDKvzV0aNUzqZ5n6ThsVEBTkwSgl+
D99PJYKhB97YJdI4hbpaei38ttvVYsYH2O4TjBMlQPZwUq8+D/h+krru3xtS+8SwBxeb/dJQOzzN
H45RKCYfmgcqIM9N4ARjCmnKSD3Uge2vFJPKf/wIqXLgrlH3M4oljcRO5gIN1U4fK4u6divaLQ4q
o3alPswqst/uBdHUYNg0EM0UBHpnSVFQv3eeORWur0ZWXU71Fb7r8xPgKvgXhEwktxeUC6I3j8so
iOsp/irOLX0tIonGuT+VBC3Rc3PW6xGZn5KQbQhCOdr8k2/PslrCC6Sg0uGNZt+6cixyVMjgaNgf
2DOACkVOjvDVvojA6I4EcvbK/FMMrM4lTkkOuhD5njSOFWxUzWeDDlosb2zF2NP/M1e/iW0t2/aq
rejE+rPqggWul6Fg0JRPkroqBzc44r0HuZh7AhvmcUl0cr7oShHKjPAAboKouwycYytrzFJTHovi
OXYQ3FiWnRBU/GbApgUMpo65b4Ikr+ALxQYvvlb5X2TBdRV2IIPEZzQAXxqQeGH/F5mJTRfFdEdp
4Wji8oBXhErxRe3RrkoOYFxjGYXE7HGGDmt2PbA6nT2G22ylBuKeGQtKHWb8zAAXdlwhaknFmAaS
LpgXJXntxIHAZWPszBft/bWrlrz8HguTvd6fbQsqhW0kK9Ke5DvGD+83YHxLTnPVDlAlYKFHJ0sq
hAQnyyCijD1klptwUOs4cFksvu5oGHAAqAF861psSmRXs4rNTbpjakPm8cK8+42XFg29XCHoLSJ8
sKzD9IuhCDEtNhxGJrph4Cp2JA4j1AdGbhL4c5VzPloM5tp2TPkoBcuikzAa/hzpB1zfpKVDppnW
wE53RPN16go0OyIgYS6QbGrUVxC6R6fZr1o674gsojxY9gpmZfHlT29zOqgKjIwMoP6aVISIuh0Y
pJyUOCbK/aMwkQ2Cy/rct9JoQiWCF0eZbUhAUPHdH5Y7p8bt4hrhSV2UY4kT5wfA1I7REOEOEXao
14gRUWaC2U9KDwiSxMvO0eFJKekQQaxJxrYz3HKDumxB01/H8tJN/n6XXdN2z3BE9F0NjxaVqhqd
G4uoAdiVrHgt7m8TtwRtRMVLyPLtJbduMRyqGmxh/rTJExQ1QN2gVwMO9ednFuFCsa9MGY36hsUP
lJzHPNeWRmdD7U1FlSbIBev73naapfL/1b/uT96Ty7zUzyRJKfrh/3OumyC8D5V1mp7/xcooLlWs
VxeXi9QYSwSb71oI8t/sV1Gz+aD1D6a3ezj0qDchtgDAh0HK25oniIoPhnrjqmCJ/sjWKI6dBgO7
mXp1daIoGZEM3F6DRyPuv8TAyfoCUNx9tSUFiboynDYRaoWu6jg3A1AGUtDAxXW6MuCU3Vjn2zFf
oap5myvoaShmoWg7SjCJa4Iu4pNZBv9EFG8l2dhNQiaOnF0sX1reEIVcNgc+oPxC2JriF20wYpcH
8AcHJu2KnzVJLMLsGtuYFg7qPQNjp4CLQSmpNV0l5gjVBy4QGVYjXW2UkXddApxjq7XZwUUfv7Ov
E9Rx0j3/oPbt+UTvVAKKbwh3AnY2JNEuFaoUnadxjRi0j+fVzMjx5kKwoMWW9yICW/bWuQyEE8Ma
+jYagXV0cJruBLD8s6UttsqxYUfcBFd9rbVRGNag5Z9X6jhY3Alm9Vq93wUM6B+nTWhsJKyiRY7B
5GjPV4bIaq7c3BKbI2K11W/mjb6QimHNTvf8hVAU71kVWuLoeqnwL7/gWjwtMziB505Zexc8kwM3
HZVz9ovx9I7N/9GD9xjWMv/vtNrfKx5sMU17Yuzj2noOUvLyyq7OTP4Jlsx3pOg/OFnl9A+zZG8C
Ghr0qlmeaaoSSxz5HKBLxA+Hmr5vgSURYjB8YVJUOizPrb3cDsGOdC8rVARw3vUTiuvRGdllLYKz
72/QSAeiV0rTcGgIODIHIMESCpLVNWuE7OyxodujW0dsrGeJuoJgO4K3Bjfc+BXmsjGircXz+kbz
qTHJDuvRl6fkoEglYydkMwSKbsILw9TIOk2bjyR8rwlRTG28316rPxNSHMLjbLW+rwuaM6FJRXZM
qm7yqoM4KnoF1eWI0wLrWgRllwhwp97T7WelImGqxylDbC82YftzHbkZwGsKBxe3sJXsDLRYbrsg
0PlxLQTw6tkAd1480R399Iy6fdxy51dDmwHSgovqu3zmuB8Z/HUBO8UBPYF7LRDeFM9r2VXqIWi2
nn4GSQmnmzSNXhYC4YJ0JIgQ2kskqLTO2/UuQzuM7Lbuc86CmSEfiTZEWvFz27l1Aww060jnA+B5
OIX3VvLc09+dFcGVJblIZ2OJDEJAI0ZCZ7ZH8mGW33EPSoNePzOdjn5qn6ZsLZqDIsCM2tG7FlL2
Al1mHuqrNVMHdzQzIatZoa6YJGCy/tyesFrXC61afyBNBlcc3x/0g5Nq2np779JqDyCoMzrgDx4p
qOaly4unufvWNqxNl0aSA5QmUyVot1Scy7go07aZZDvpIhjLO2Z0ScKYKD7Dv1WruRY4McAQojQ6
hsz5pyXf0nXg2wzqQUnpTpsrnoHLWAvmlGFK+izdfNRS0DguPo67TEdbIarpjvUQS53xpaqHTUID
Syn3kcG0OIYzfyKFoL5jFrJPkJpu+ym+TxZ+bkokFpSBm9NyWHTZnzHVGDkPYy6yu3oKWlcO7TQt
4UNa06c6zbSrTku4BpQbwVXlf0/0Sm14Bvmrpjbe7XbpswIIhps4QBzDl9qyBTANazLwXBY1Xd/Z
OWhFXdNlmgInm9u+68qscpeVhQAoz+uOQIwcpbWh9GUjT2wVohT8mS5kb4ZITwJR12eJCi5JhIym
0m5TzpRPaBbSpvddvrGwYK3xIGnTM1E0IdepTsQya2FoVO+ST9CMICjt0qhn3UbgzgDeIHhytdcb
fbJWrAOZeuo/IJ4Ye7ABedIQbZFnZ7hPtKHnGfCm7J9E5ZqCtRCMgeqS7R90hTJ0qMFbhFKyOX1p
iZwtcUS5MIZKuWhnoHl61EfLeFux5rZ2rqyOxOM0Gvl9w0lY3Y4J8i0Djlz7DQuA7iuK9DxbcWu7
AM3jGU9oafDZFVfEzCEX+37rnrnp6NfK62VczxMq7oETXVYYB4X8gcPGLFPCPem+D/KH6LjlT6xI
wgKcn4qkpMdNoTJV4ndlJ2Z1T6OQY7IMf8LvgbJ0GnMBp0ehm6VJ0p3PmxT61GOlpl3Z9nWXQvas
Vknq0x5vqMEMlatoMaoWGX7ZtOhNReGSqV6KBygUhtglQ9gnjOdFyR3wMCYMirs8Tmg/NAjNtioA
qAnglsdr/EW4/ne5p9HCzUmIF3OX31ZBu36jEdKUqq9reBlW2y3N1vBbO0qVaSQy/EDsDG+2GJoD
gM/Tfgttx9qZUtHYcmzTjS8YjYfqXGIpL9W9bAwTQuDIe7bmXD9bEUBS2juPtP/Jm19MkG14YY9k
I4PTZf8OgxzuT+UcT/3sNVdkB/kMN2hI0wKyOqWHYggo41tntfHvJNdpPQUsRQzj5lQRnoXmn48+
S7e2lKiT30zBAcX1dk85k/GPgIW/O53JrXNEW7Bwwin4nrkPHVBaq3qHmF/WJ6hn8uTUYKz/lZiX
AtV+TVX9ZWkQS9tSyC19he6cC+K8rXY1SbToTAh+PrFrF9tJdglWZk/vrqRBtQ/cZF1AT0isAKfE
0YO6sWMkyzwAdPZeJhoQMRdXnNq4xx7Fsh6/Pg/14ztHZa26F4YkFYNn2u4k9C2s/bCXPKdlE+L+
u1jDOc/vVW9TYnUjdrK26iUze4L/uyaNravoSeS2j1CEKdY3r9oCJhVEl5HjTQ+AxeNUKZ1LcWnp
XImtHcV30IhMQdrzYUjGvyretfmPpsWGOKzzmcLVtsdaStd5DGR4MHO3ejSBL51vRDOjdS6qefAw
CfdFXh0ttqjhBFbfq9zMfMG6AzQ4V76tgvKwHnFfZjcm9KMdS2SH2gOcyFVNMP1PX0s1Oz2aWNPt
jKR4IdHZGlHNJ/Wpk0y/Bp0ZmyLPOc+ixrraFGLddK4plEeiTC/8hn5ORUzhYABclSe8It5Zpp65
qF73+4MRAZez9jbb6pvGW14B4sitZXFkgJxXIppIuKSHj7twpuRqMWxDy/VblXeadFUC6YZgTUjC
I3UOxUSjzmAhuJLlahAvJDi6uYJGYBUMZxsVcNZuB0/GIna4yUnU/NPieCNS+kWDu7gffXsnstUO
U5Et2WXC3f368mRyLzF6ueeyWAnUXuZUxKhXU6V5BQANIEX8wYmlg0ALIJfWA3uCxNQM9ge2aphZ
WP7sl0PGDOfelTzRxJK7j5w1+RIxWSd+6REStgdQlxUG7785rf+62Kn3Q9j88+T98FkZmyhs4l3e
8YAe5izivS8upychpF+BVZJqqDJNYS8WLwkhvvjfjJ8z3mZYUxvDF0yIAfjun0HRe4HFjlbeInwF
WAvbsQJDckoDTVxQWeX/D5xTMabyt7aHAW9rsQIy/IwWogEEa0/Ytz1vjpYQOnTxj3MHeOD9u2ru
nE7ifUiWPemUE7oMBTXDWVhvwkpzyDnusJHRMu+pOIF1QZNotezN8dU1qSOVE516oBSkNDlh5iGX
0eJzjFJupdDNNXmUhHyPjv0/XmkDvr/VlVLupe/VMXnjVIEzZL0CEhtoWGekEdQzcrSj1aqiEr6i
7pTbpNfuJYkDVBY4tWISuEwvjtoQb3ZandD4+7fiqoCSkWI5/qq8eaRdKWW5pLfHihS3NPJbtz5g
VgVBM2ygtVJBkD5p7ckRmUUaOB/F8wuKpLbJzFxVYCbDZkUvX1wa3W9Hb7O2YQ5B4yIyQvuWpiSg
agZchYTLPjEG0yRNOx9rnfsBCq1UnU361GBkbHvDo9H31b63ahyROMAW7Z8Vxyg827GB3EfanD/e
8O3pp0fE7q1SfFnU33/KiwRDzrBrLs44bJAF9R+/G30//BpYzsrPMoVcdNDVV48c5oHdZjsx8c/p
7HgmgZpD5QqrG+hgLSkydSr6nu44ttkgR0iK38VgATte3In3BnSkag+RskgpTPQx1i1lFtJcCgs7
LryIe8yCV/7+iInvDC61ysCUebVjcko7vXmK5m+FBhN41Yc6Eeq2cEdgF6GqEQd6MA7Amw7fL+8l
JJIjoOKeyQJEa+qlvf8+asWpTCMsG5bLM7lfVfxnM9P3Ud8giG2DHaQj4ecMRdKXw/+pnXiOHSEO
IijAFM9KEYGmoJGV6n1yuBFhOt62LUjBVhNUczNvXYH/W+vf6eJKsi7c5/DUUHgTyFGzfIaaes7P
SFP39QL+eEQYJZ229jJKZdzcKTwV2vQ6wEfrG4f7QtAj/R1shrZO3zmUYdkVkC31RAsa7G5huhwM
LEJ3DltYKPYD7NqhXffh7DO7PfxnurgpEdj87Oqj8Bs4+OKQI7l2a8cszYkZfTIjUEqkgyENDQTz
QCdMJMB27vpI2oauyqhpRGAsx3S253pElcl2GXXkM6gW7f65FLepTqYb1uYyNKos0z9TiefXFuC/
8udYpVNRUT6VtDvgYhrLLdxz4eN5Qpx4RNSheO7zYir1JsMTJTPsywom+oN0HnR+Z7/KrGtf/cwO
ccebmzhsmWW+IrCvDLvPA0t9rlwXn7yY9Vngd3oH6EJxIf6vM0NvJeenHfjrE/LvHZC7teRubH99
ogUqatii3kITRpprQXXNHPCrGuTXZEKVny9bVUCtFg5LqEQpljcRDuEzwS/hpxYFCDUwO82a46my
HhU+WQflRb3Q1uh7A0Ft/5hrpdQ3XXx68T2XYwByNX7gxCVbHQjpBQpwtYfHjI56KAw1dJbdeA+M
juEMg2HPKp9NcnWvmpGbyl/jRzjfxNQzupso+qzuXbmoZ4ummTTILIa7qJsItk2qrOyuDSZt/VRV
kb3YGM35NVkMJVSMHxUlfyCIBhyW2UvoeZJY/E4wGr9lAmwRinBvJvJny+sqDQ7pWXDkZNNgSgYR
8X6hC2rYQBiCH1qA2UZyALHU1lFAQOyhJPv137FOpi09KxLejPsNBttI40D/KbcjY5NNa/RAfxi6
IF0lEtaFzAbmeVEub8UQJcwMY79kJ8i3KajEF+2Y9D/iQP7w3A2hIU9sRLXgm1OJ0Pf9niuPz7BK
InjWjT3BI1Plj90puK8MYX3I1GHtf4+0CjXilJkD0m4JUYuriK4AA6sRSL5B7vDHMvXIY8LRYtRe
pYOd5FbZznpzAOQipA5FyrgFsb0IVs6F4ZBvHYfQ0QcU5EwEme0XZQkypvE9k4o7r6+ufftcgt9x
YsCwlmM/Gzcjz+nI3f9E9GymwMy3N4MKpY2ZEFI/5pFKnXGL9JhZ7Rryc7YyhxLG1/ljpKt9+3OX
UkTTaZP/bW1XtRKn3gvIVf2HHHvAWNQM2bbXfcrN1sbbr25rU8gTkLyKBz6SPLj5NUdNhhIIsLPj
bU667fdojccqu1xub/nUNrOSgqjv3JS6Ac4m4CLxBUiPo6LRhOi/JBr2ji/Jxt2bta1+1eKnRgBk
B/eAQ0CoXB3lknWw4FXQyckrJTeBoACq8L8h327dkPlyybQjb2m+WT8gx8M+O7u50HSUVNaAR8nD
WGQtk3/P2m6x13q64q1keDmYraLNTIuWVVLsNH2knCH5yMJXO9FeIXEA2q/ZqotCm/CtVGCy+3mX
aslVaap5TbpIZgFETyFDJJWboIWtTPSQrMyublJQ0KEQG5orojJUxw01LmO5RN3uiQmEoefcHnJ5
SkT7b2fGk1X1UMqiY0HruusshJZEs/0uFT0jGnYK+hhwWEUFD45gz6WNGzKHk9i+s6m5mpsbwsZ/
2MGRbCcVfzBRCfA2OQZWsFhbWkRxrIRUDcdzJ6JRMI84g79oKrsL8mCVkFTW+dGBRVn4Wti8cf1C
8R5tuEgaiYFqrG4ysQXpzyCbTE8mgTNEXDH95eQoxbuSbh1am7EsVTt58/1ECuTffpIVjx1IGf9T
sfDLSWFg9gNTQKliRNPT4oAFpfb4J02+vxDi+Ya0+or2niM0AMhOf44f8wT2/94krH+hShnfPEJ3
CLWpp0SLuxWCVSud2VJ3MGJHIw9WwkXSTmC/qz2nIz3MobrkHZZ4Z3DpIHixGcMxed7de2nROe2p
bcMV5ChEllBjQ6eQggMd3vVTjSKVgJ/EQyFiGJRAM+02atflj8AEKbN/ZXOa96nchm+JdDo6A5Nh
e0F2SniRkyp5zih2mJTDnY68M9vqUref426NQLzrdxVTwfPcZcBbT5iIPBK9vOBCr6/3yCo0a0TE
FdoeQ5X5HS7QlPp5lne9eIxhnbHINrLXQ7k7EYwwCnpWTyCt0tQJbKaj+q/SAVXbXYG+dLfHgkor
JOIvjPNeLGKrIjR5+iuPrwU9px3KKzX8jp/oVbc+X1JMh6IX/oEW68+lO5GCPihEZB47ILn0SGWb
N2h2OaGG5dNMuvynpdq0c9jXOuTnD2s23JiHqtA5HywfchqIg8pDsv9ZCnh16nmkkeGVaRFr1dR4
TjLIs474kRHERHNc5lTdvDhSL3m8kXnLY9YlEGelRLkJrxoP64MY+vHLPfz7Jj3SZZp5G0+7J4ah
GdbAf+XuihrxPCI5U6O6QlXNXESzKCZsNCEdFtFiBtJJVySEkvKn9v0BjfmgP2x5ZmKnBAugIarG
3vVhjrH/lk8JmQ7EPAGASzc0VFKaR+tmvbalkUumYiVP/cnXKdFEyY8C8yWfyy8UA4/B2tzlBt+A
WQ9EKvIgwqaN1DbSpI7AN2GyeZe3KvEdxGH4cIMPVv0y1VmIUf/iHmsyCRO/46CM3/KPNpkGWR8z
8iZSQRpwiUtsuBzYzmzUCWC/LvWHxellghM1UmHGRyyRGqNCVN5QrXhNEtspWsi+RvAKiZWcRZfV
+iOJ3tniPuXoOBu+YI83RmEeMI0mqJGSmhykvx90JSNYV/u4r52NxI5IWLaIte4iH2ZVfwqhjyuR
NuZ/Dsx/BkjK9+1iD+yas76J2BWE16JCQ2hwLJ3q9X6curblvlsPn/IpAjYfr0dn/4M3V8h+sXC5
zqm+TZZcxhvK3s8I5UgwZEOfDIv2Aa8zZ+mPl9USfF5DtacmIFHq+571hDj/WHTkBwt8s2XCV9Q0
B+1YlknFZ5nzeMjBNaOc4gX8lTXRztN3opH1YaYUUxyvfPRQ5HGCq1vBbX/XIIi+Z9ekJXNvB2J1
kUjhD3sEHLhIHK85bVk70tEpIugB5BsDLTl9W6jpojnaN5RldE4d5SLt8o2aIbCL8uSBA8LXm7vF
ZzAtCHPC1+Yuz1yyTAxheN+q5SNKmwuFjpnTwITGQR92byJzeR++t5YILNjZZ31BqEt0t02B/Zt+
kTSd6xuBJifBzgtcCE5OXNN/se056DUHdKvrpJI6SENuWitJz6gfsNmQq0AxN3CSD8tovaL71oao
HOejQbYnBmwiqFmiNS81fuZTUTt6WFAn5GF1yBkSpQK0gybw4Q2KDgNxjX/LqRdv21cHt5RrMKv6
+Yor64s/DEzvtzYtPjmoyjjL/HacD2jRN6mgn6Jbo7Xd6zdJKfXM8HxnR2UWVeKXeiocUvUzTOP/
UllJg3AAguZRE7voNzI45y8BXK2uh+rTQGsZaEOXV5LVX9t2lA4jS81/6uir8hm7oZWiMtfDZ5hW
HoktaAfAdAnZAHJDTSbpo47j2vJ8nqGDhqAppxZY3sd49gc2VzqFD+xNVsrycgZPmhDc2+r8lepK
aAGtz+emk94lOeOHkD8catKV9d+HCouPb8em8mffMO/IZXHDlkl9zuZfuocEiENLreUP9aBF3qm2
XZLTPnFH27uFQzrY7QO3H9n4fbnYfrdj68GsCpljwjqTXhMpS/UUu2/ZI0rxsARNA9NPj/iTiZRH
QbW7OCdEyObJuhY0Igo0aUp01H0kF/TzjBHsAT5nZRXm0OE27K8Hn9z8HJLgZ9+TphlTNHd5nNLi
q5VgtY4en+i13fsCnuHEr+upskbITmHLZFB6xiEsb8zT44OG19ZUvkjbud6nJQ8+yITksC3VpQfo
/xW6rW25xP7tALI9g7DbvPhr+JOxOyaUqqnJa8Pq1Knuuz6QtM8wBgZuN0pHqYRAfAU2tgIW1pKp
/ZwrQXRQJT1SKL1XXMMZVZ5ZA6t/t/VfT+QZCD7aYndlbMZMyBxY+9xg5O3ukeXzZ70o2cSi1Rt2
FRE73FOoMa06qQiLC/WBUgXX5wu8OtDL3Q4GNA73v9+gjnDrV7SsjRHJ02Sudgj4RZ2c80a41c2G
XiploxX8/KsV8179wocQtwq65NeaLtYgmPLX57zigU+SDEmdIOliuVbXn7KnzPsW4Z6VOsAevv2Q
kadXDG60LQfdeUbH58D+Uq2Y5v4775e/v9iVyPnCu/mEbL6gMUInOSmVPbuAbQWG2TluCGD5vWIw
yUl7XzJDx57fT1A+yJpf8TiWsYrY3DJnmVE51AEPHO0f94ecddgpUR8D2n0CkC1sfcGhuH6B2GYe
JHY56QAYeBRVYPcueIqljuAAFhQU+0YbEOX4Gdz8SYf76iiVdInuD6efXy0NsvprIv4kdCHT3Q4S
6d9/OCoTnTrzK5ZYU7q7HfpKRZ8Nn1pW8/5fffX8jZDFLCKd0W30qm9nVIpUKQoX68XyUnZoAo7H
HYMJB5PxrY9qmKqaAEoBptX6Lo19THekVMZkS9nVAoNLq9ilJWcWJgwQLmnhnhSvrGWaieVA6mOt
1/jgjiP4dH4QpJZwq0PbQ6F94IcyNW6wU54vXANCdGzR2oTY3/QhRTxN7PDNb77em6414q775FB1
GZrhTAnLU/W+hr1wsoovMlwKQkD5al/nGTmpl3bNoXSgLElmI/7cUp5FaGq4An/PoaLv5qNMUjZf
NTo9ffHX+TkU/WM30jInO96f2EzyoAMt8vbL2b/0JJNeMPPeRgFaluHQ6jPGJ7+COam2oRKGV007
TA75crtVFB4ISzaioYuDAS9jjhpvPqvClA4lIII1MHtl3Y/IyEqT0PBSOa7OW+UA8hSiM7JwY35v
LGGnLcVBpq68rtZpqiKQL3KYFQQpi3a5xEdRFw1Q5Xx4E3k1toyvqiVNaHjIt32oTKUZKU74ylwi
vDDdlmSR7Sf/r+gfCZgIAZVBDWsaHRAsx9kLc51ew3JReqsNPYPluiG3lWpH40Vdhfl6YKaSNFEv
G+SIHWiixSCOisd5U1F9Qo6IOSTrQKH1NTKlt82UPbEGUV6m9+Ubg8bKhe1VNdICA80FnaIwB4SG
XFnHclXD4JI2doh+O0L8cczqXR01QM0A/QA/pEg6SOUWG6EFx1LJri1rnznrUS1ODopEmTAqOrhY
XA7eeAh4wZTf8BAtPzXCe5R1cqJtvkhdFypKRnKk08/0JYYdurpx6cnAblGeGh4O3YVhxUL5gACR
5PG54ura1U9s3KzS6UAYkoGnaOh+Ml1jHJzr6xAMdRzUPeqwxwtzhM+cqLjfr7hPxZRDtxgdz1Po
6isA7YTO9ZaM69vguv7F1Rid6GJ3pNRTeuBhTnF1HRZs99+Q7ZmC30Gxl9CwtX3K0MQf6dxC1j4M
AliV8fKie79BUvQj4/WbfE6Xsz84nIfbH6Nd2LuIWLa+d6pCefN2B//EEane9Fjib1jCD6kvQao3
HDDU6wwNqKtlMxW8931MJiySH85lMdc6Yqj/m2LuvaD1/Mon20WG24ZAes9gvpsTLInt2egC7Mr3
sZKHqt6akKKG1JayyMapJ2emVXhu+CvrDOXPnmfvR+7Y47I3yYLAZawSPGOtihkSdWrnGVISuPk1
ZW7++uZxk32YZzsZ9Euk7q5KgfoCxaPrt6d9ZCSRpsIbUj9+vejunG4lu0y+yayvDbavEs7zlegX
qh2Nbndtin0LQ74S4VXk1hIeVQolPDoHmAe9ILMwxgy00unRU4gl8Z7oVvcVpDtxaSKlikf7/yAU
qcn3nXZzWT+mq1Guhu+v3nrUbubP5ytXPBxHOHiORtO8g0nBzXaEd6cahm4uCADqBQf91r3sTnbD
gZNTpSQNsRznCZH28fO+wdx0K36E7BOfFTirvL8LuQEdcaOyK+uasf0TraIdClgulCUwnEMbLFkc
ki426N4xm3iEJ0QjrZvSG1na0d7DUY3PSACChs1/paATH9CXgP40ub0g6E9TF8l9K1qaCjvvbLcQ
keyzw4+mnQYVL97dN5r/32QqFxemw5lmPAGLOh/gCXgT6SBIqeoMLcNAm2VyGTz4SZ9yzwUdtlPg
OKYqH/3z8zc5mCyWhTnlS1i/1lr/8v5qm+skzZyBSWhr0E60mZWalCWg3Y6ggWWFPjX4UEQ4DNQs
qBNwbjxbzXHULbX9LaVeQOhvKDbXnvCWkPzaXo0j2J9Ve+rBcCSsnEuuz8Dm68LU9CmzEXxP6fKs
bI8PfNh/I2ETMxtFxWnwO2C/nSeJmte5orpFPJOq4rs92mM2Gk/Lg+gRc/1Q18sThAg86/N83Yon
Nkbr7xEKjsXVQYYXetwyBJhuIJc1M+wwTZAFAu1nMPSClWg2QLaoFKIxSCQR0YnlMKZ40YwfUV+S
gCM8AaO5kZf46aKBf/xEzPVOcFHft0pf2sl4RZ0RbiLxlZ61b8URY70a3KzP2K/7mH5b+XxE6veW
Y3/xIkkNqFMlOSwu8iSmxHD02ilwEAM9LpXRSUOdznAZ2eJl+h7xFSpFf7a0NFgj1Jo0Fe4Ny3yS
nl7e6yAgwNLw68CEFnp2E2SBLNTimEOPqcdJ6WDEOTO56JAls+rnJqz6jAsckWybz7UgZJsP8u6t
0HduMIXUVuAxWwsM3PgT3jwWcCNKaIGmU8lw2gWFVAN50cfxOlcAVajIRq2frJlXHxI9L/MwyqYt
GSN97iCgYpmlKOGre3A61LCjaUimTw22sXlcKUlLy9lTuhtaAmhZnQA43T6kSCPCNue3GG85VHth
3O3kOODTn95oEpHm24awmV9q+n8wLh0nMFNlh5w1/EsyKJtZ6GbAsQGJANUeIxxCpYjftJXx66tA
s8KJjXawFVKIVuq1QdosBRzf6nRPJN2QEvjB0gOVy1bA+jdomGZBwwXX6t1AUoCuDvckDhybEzz4
fwOlWL/EDvmNpUHOtJf+r2ZoW4gJ8amqFGjYjxfcIWahp9fXxDbZ+gvRlQJ6Oc6Hr3HaSEw5j2Kh
F945B9ZY2J1zk2zOo0mTaHhGnInJO74Lb+aHC+PfkbLGK3oPpu1bGfLNZ9/uXdpCiolJx/hwfTkU
3bA5qMpOjPrKI6P7WlXtSQBeSjKdgs6HnzYpetR4O1aZkjsIWxsoRrEH4z9Jf2e0RetAJ+k5wRix
ldi8ct13y/+qEJC+7chOlbpNbgCsVRZxy6LYpKbm4SljhAolCVfQvsIJCh0xqzMUo6ivvSEyoCD7
O8uqqD3j+05tH3yW6DBXmAGEYkFud4nL0Pnjsi+acDNSsHXlKdANDOnrnL6oS+gIa2y5FzwBTvVJ
2eDXig9PPHq0PfN+XHDv/8bqMQycJVUkky6VvuLBGqH43hj9YowmG+OuMIazJibLyooLAdUZ1Hbz
rX1xtsro8WbD8X5S3Pt9Ormr2RI1r65eBbNZv/2C1hgeJZNzOCV0h4xyffgz4lrx5KwPPOVisbJa
5OotDWt4zvxLIStYyLI0jPTI64HnFZCxdzHK0vdHO03GqlEN6GvO++I+wpJO/ZBpMBsYj4saru1+
o/WkKWj1cKIqFm+qTY1jj+lNckFENGF8SSNLgboPmB1wAuIS2PPIefYq0DQ0QHowUha2iElX0HWD
b6CAz5v8akBpJUbqzP6Z/lt/rChrhFaMZKofLugCa508iUXRoYkf4YnCtCfdKH72H5MPHD+xiTmj
6bEQU3YwI/wO/oTlLfEMN2xB52RlQi3p08NpCMYivriLIuo0DTsCgajrnn/FY5qCyqnUr7fUuG9k
v1effy9riiCmOoI3WmvG70ZJyKeyG3/nRoanQ5NhnGCtSDbJNakqyC+aKLLWp4tdlDsWkH48qE/m
tXcnEhe9CyJLxQ71yamD8znRGNRJKbJ4p+sVS/tvmJWoTQyCfqPpFvZ5Y3r37XvR7wm1eJVxDXNW
BhmUz68FMBp9GobFu3z+NAJXy8wEZdShf9Suko05MN3foMNQJwOpVZJmMfDfPFpuHsd1GWJjblMd
dWrph9Agb+mjX8M3mtS4cheBULme4XTfXqH5QKJJsO+3RIRDPadC/XZdBf9ItDD1rs4udjfw+GsJ
rWZmBieATu5DviqBiDRAXTScPZvk17aoNHF1GZNpD21yVN1YNzIIyj/P9F+ttVfWs2+4sbiqo3/D
Xn7m013uLHyG5/uREZnFZ0gUDsUIYrgJfcdnZygaOZGR5Wwygo9+IO80XR5btezrPknea7o2aWfK
iudky2asieqsUFeMP5l3KJYb7jsMOb/Wi+e39ykgE568TyuGgDAKYReJUox20AFlX3p+tMuxyMXs
a9xYvNVNxC2K1TbwrgslLrtP6nvZwIWEJpmFHTpQrIheDIBFbmuvRi9E55d6MMm2vF3z0s2eXvvz
8RPaU1RhhJt3hzdERyWMlVUYmK4LUwYOCUZR2uoNjh7lUDQVaEF8WC3E7cXab4/uQODJvGtGNz8y
PVaWwx5YW5OoIf8Qxr5YSTqHdSyvJuDlLJb4arp4z6BetDPJKTebmnfsl6VaSKL1rIGo664u4pTD
Grbrj88hIQOkHXpB0C+hZeA5fTAR0WsMENC1xieSS7PKyoO5iGtUF3qeEhWjL+9rd/ieZJPaF0Wp
M8Kfr8xy5NtS5qQUZD97yf5XnjRqCVnm2EzxOjanMKHy4lOiGnkgZjbBAg81A2ZRQuMxckdC5YTS
ejIXzdUhoSw/Anvo+5k2xY0318Q/lDCJymO/vkzlR8Uks2AohH5wp22zQuEYCP8gQpAmyHzb5n8e
PSUYgirb0HLStJvwKBsNayYlOkB50xv2mtqRcmL670e+NPZf2VcyAJNvyq+2h8qhGvGxbLRuShKI
pVTD6mPh0AEKaleB8Ibjp1qHzOO0aItS9c68u4E2K/XA2d6Q7ejaTPAetxx+CB72EDZF0in5I0E0
BNsL19uVh25BZcEp7gv3fH5ryDaf4gF1rY5+UVtrDn2nDhzF3sf87iBgZQrYwUeD75eHaCdBtpCW
ktKRj5lCONDvhSFHTojWXAe46tSBIzOr4Ptq7/mkWNK59N8TlQWS6vswGNg4LKMWs1G2UoZmq4Gy
k3zXxeID6I6rzdDWfoftNBbGdl9oSE3oCbzLX24DbewKNLUYgEYFithgqe3CVH8okvboVEwMLgsm
1aIcH8IH51HNTiYtSnOigc1TjOV5I4hSUbLa2mM6dtlB8srIfH18m8LUNZFAPQBicHhXn+A4wOFu
lccZV1VKXnkx/dvGi5acZZoEvCoy2qLAPm2E+oDUsW9MOXwUQXXSmu5p/03LLlKzk4jdkHFPxtOc
QdyOiBpPI4xFhe2kq5Sa4CjviaamVdOb8zAFHz1jJoNvGyMuHG1dFSFWfH6lu7qyGA39XrPHjsX0
Hmeha+Ea8E/oU0Sv4SazpKoHf2spE2ExLXOTUl15/SybDXsXlkglMqE66uiLghT9Km7foSTXPgSn
mDp9zlTpLx+gepOM+9W2B0d3CMS8fudygruKU6Te4YJf/R3c3tAaKmooZtfwHjfaPPueBK/DXyD4
t+CIO5rLUY5kSy8xDk9X2Qql/qed6k7wDXe4XR0kn8cvgR2tsTbWvQyg/aQEBuVQwRUFkN5Iipbx
CTDy1QVMzxcbtcFQuK4C9RQHos/WryZJnAuLqZWC2z7hlMStzvKNlniMQoMP47xbLKXN+qT4380I
+sP2HPmRwXj5Fl7ODYn3vut4OiVdZsc3/JA0zcb24kC5i22N6nP9te42xOwS0PMfbahUzZsTRI3c
ZK+FAB7tvbfptDKD/FlGtWHxNYKOp6ooYrYSFlR7oVuTC0kK+pubJlNF759RO7RdxF3r1wAlAqpB
Ks7PVEi802b35qrTrH4dJAzbCWJ73uuVhA6Wzoj6KmtDD2A81V/vB4d1uzDg7GgL/j8vFTojRKWz
z3JLKHzMeZ8Xc2zTvGYxbODO+k9o12+aDlQn6W+NNo+skKfcbsl11+9d55czw1BEXSkotg7aOyZe
tNUXvD6sj65Jkbd+mg/u3OdB8NpINmShqKIH3kjD5BvDTffxEQARrpr0LPnboLfsmCZe7fQ+oQQK
3Ch7NtLZHc6mo11+dxhQPluf0nSAy7CHgQLWiqISjOGbr6zOlUvJcA3F23Qz0TQDWIoPR1HKWGW4
KcYaT9NSqELAVD88Mmwy4wkgPyA6mT1vvv+LTo3zGpEdeyIzn4zYOfpt4YY4SwwWW8AZAilvs5td
7aoRi9GaiDgAzlP7do2DxD5oR/5sxcAhv25lRfbvZKda7hOlIFPNXJbi9Z1kZ4x/As9WHaczl3xN
duklclDSW3KctUIlUKmUUojIJv6CnMlrwjslA14ZzsCw9TvJz7jYYMoINAylaUqEz/7YQMPK46ek
8MOFoJZXu9XjmXBRRinaxdKJE0zOnMLOUDV10suSETD5avcM/puwibL0MXYgpETHhgZCFt5Z+E97
A6QT9grNHuG8aK5m1plcjNQRODj0gcHmhEErZFNy6kzWVPczZ8iPPndxZCKljJUxezTNb5QMr4UC
PpAoDDajVI4CTQUUD4cWH2ZMUWnAax9LOF+DP+/TYi92kxi5Bn5o2GU1OPKhMmDKwx8HZ1ckJRAL
Fg3+SG627A2nM4nnmMLCgXxnXczMQv4k8E+tFq8mcf4/iS3DoycttQP378IhAvjWu3wZKmj8cid/
wqPGiYAbTgkc7KJhL0bNUSULL6JdGQaAlaW+HKc5fVLCXvd9a2haBiO/JnDMqeXegsbT7roJbSS7
u1xWINc0AkwJeipPLAB7wLIi1Mn6CAeluCh84/BzxKvYCOfz8UtmhKX/4KyqDKO5OlFUVGmwxNp+
F0l2I2C/MH2gNSYHO3X79q5KCw2zCBzxa5wy2471IqU45BGCXOPmbhlDk+3PSU03aTVLDgvAkw8A
3Se01qNfED0ybD0nU6SMY4pcwR+CsA46fp+qSKVZlnAZzb+15EJgfg+QNtrBZU3FAEtIt8OakqrC
UO4MjdLEtu2bqzFncH2L94Havl5Y9I3nkU0OcRo2/wTrMShXpnkeigPIZjNpXiMnCtgmFM9Gn8cp
DIxtR6V8iCL7Q/ERdSeDcWcHEiuCWJiPbD62WW2Fl78kVSzjAbUTMRw8LDo3OFa42l+tbDMdG9zM
oNhbjf4ZkEMOGMNffDd/o5Rb8y5oLfd+7v4MTSg3HrsdnTYtRKY1U/7D2vKQ1/Hbrrp0KRNgx0I0
1HOiVT/a6CcwfbXoApKfK2jJKVOG0Qraf4vNrvinyjNKLaJiTLKXmIVSocmn5zkBPiK/L0MQJd9s
rl7F0KFKesvQpcF+SnjxR6h78u4jsp0nE/Lh8J/eCNBrwCx6uW4JycR4QLnnJxQTSYVy7Z/uWmjM
p6iUtVKAZKSQSQfTMY0GQtfW1GeOTyePNBGfwAMXlrjdWdeCGK9Cvp5ciGe7aUzOrMZfCUykGyD8
OWoBn87Yj913HOg4dlSXotF46/b+phn5OP7BZQB0dpYgVjsSA1LcHEhTfwBGzRO/a5BgMtBKvFii
lXN879EOF7lxcGOWSrlY7h6Re0mJKC6wOwsqQo9A7rbBe1d652Mt9eruWVrl3NLWC3HJxU693iO2
T3+ViZheNFecqhaK3E5I063k2XmeY8sF+rLbvZJJEpGxc07bRwCBf9wMJK4Rg4CxPkQMqmkwM2uy
s5yNS9QhmVkc4ADFyfT6zE2c0jStaaNP/090osQFTTFk3UCO63KZcu7NSGF1O9DHN94roTfXdUs/
agwtRUuwBl8KarknzAPu4RllYKRFo2sSY+ISbjYiVFESlLFbQ3gp55jCFpo5MAdFw57owb692hy/
akvz3xsUwyZPtpNFBbn3mISlXFPfi+UDCtMf1PHjyU+oJY1TYpDcxKNGmkuHZXjWNB3zq01JFSRn
TM63KUS32w7NxwwdU+jPZjB8zGdYd1REF4W02ob1G/RIIZPMhrYo5PWd5+BqdPG19fwKdu9MK8L9
LCSvH9iH8bv1Io8tdU+vwpcus7YtxM5Uufg89MEDUvTGiCW8O8vwauOn7057gJKOeDN7oM/N3iVB
Q7/4ttH5X7fo5+rSY0JmZZgJfdJ0xp1d5UnwNNLEOiZ1waP04iLAsOAvV7AW6YSNxmVluM779plU
cXZUNS/cUxuolum+qqgEm2xw16c+XpaTavCYj4N5asn9QHU4qsMmOwoWn1pcPSrAAnlvOHzlUx9e
DXtjnHDzgTP1g+GsoSw1bgkce0iSCXQyndVig5SmfWJ4tNjbfrsVd6yWbZzoDGRvUbAedk1W4Br+
6b35UWfx3dfjgkv2uVjRbjsagQ0HEBprISrx1f4A8OGOOUf7mXkx6N2xvSfUbjpN9DhMrwQQ9dnh
HLNfCWRGPuqtebutankyOpws9v9NiK8tXMMRtjzrL7+aTU0KTc4cyQKw1tjigrnBT0TZ6tdGLdjV
GrhbM7R+J4mEQhCemb+HdnvOZDuc5zpbKrH38VJIMZAvFGJRHlskOCDQrq5zqo+BZGDVPAtAskxO
0ZRJTSBY8WydQTaSWvI7OgyBo2WlDxyzvALXg/HF/LtfYTIC7rpQ/GpjRpITMULjW/HwP/YSR7hF
g/S/2aDgFGq/AAdJ8bIGy/PhnKU8qQ7XEcebHk+2uwd5uA+OaXSCLtoT57hwXY7jNj+dEZ+/dUGH
amiFmCbtZx75bLDXWc3MRRz0403nq6QPKX5sh5EMPrXRMci1An8LX8uPe2rK4pHBwUK58BRKWG2n
h0arVwSj2z4FhKvY0rJoRS2r2FHExK2lRZZ2yNNCwAhy9z8Xm2xvg7o38JxPV2Utj7isc+1lGM2Q
b3H3ecruknWY8hW4pnaH3CemNs4tw+XeNbZRpXIVB5Fw2cragoZaxKtJZn/gGZutlotlTTAvnlJk
ZmVzNaDguyFU5Aktj66sk63Q+aXCMCQiBHXuz/jGtWKDCziCSYzkZAO0ptGpqy3yOQuTi0SNAnmU
9AiS0cA6qBrchNoPflilUEtt/JbldiTKA3NiuXOia2dTILedgJi/avPoa2u7gFw8K/6bqjz4Jes1
f1RcuFHWT+4bpU0vIvVMx1Ot0aWE5W00Era6pPdAJqK4Hwza7MXL4HHRhKCMUru5U/k2K9XeY8Pl
lL/fZuHSf8STBO/q92rwQMIxYUob0R0h2kKGuCxNejZiuaY6bqc3C061jn1LMRKHcV20W7ufqii3
3X2QzjgQRJfomIgphw2tHpdt7rBz4V++8dcTmv39YkVyHgJQdMMJZFUM4puplc/9UP8G4uglq8jX
FCEAvigohcXk9FTsFcCtOD2qJ0zg7NhnYY/QW+skZH4VkbrShobNQLsBTSLQ6zRHK14lwC/UIU0n
cKyKx0JwqZ+jOMA/xkB34rMnAKsIfT6XSxwb58aBFnanpXHrdb4GXpMfvd8YjkoosVIlNZePryky
MyQsxZbPoLpPFO0Nci9IQ6OiuhXOv5jWtQ5QR+pWO/EP9mtnt9R38rENMCTmn5QSQweg44w4qwxM
ymuSaBdmSQtQB+Wp7WUpeDWETkt7rT8oFwDaM8Qi22ekGqYo2izidpmrYNyCgcM66zs2EH8M8TRh
2JcOchR1SPqpneVjBIXMYSb5gy0EkkTxiRQpvlVMUis1xv8yix07HXv6IYiF/I0PDTS7Pv++v4LE
3YXzQBD5Xk+BIfZQzDPC6+MQP1+PzBvrCzRloLBXl5ea5pStsyoAn5HfxG/De1ZguI0YTou4KTOS
qHpaPwnLbAb91C93jMFFraXh7Za0opLhqhPzk5bLgjfHrNDWCJfFJz3sI7u34ZI3sULw57jL2OTj
wh+8qxbpCKjVXoC036/J52KOnIV4RLgsnnYHCKagqjxL9YVofbHfos7HfKt3UVtd2bk1F/vGw7KQ
MckIDyDCiPHy6u6nr/7I4U9zdetkIeZ9DCUpLn5Jacqiw5LJQsZjkLO5A8GERihKsNcN1BNyPD1t
mLLyKnxVK3AR0EgQWZ3qZdjZEaI8x4zy28krAECFRqCxLj8aO5DwVHMcYpKZJIyR8plWiSDoiXSw
UXzrCn+Jt1knhVHCcbq1GyL9s79e8sL7TzFz03CobJbjHLcO7gHSh9ZjhJh3jMPCzQsUaVX1gcCM
i3yst5q5nc2mY4V/Ycbt1tP9xmC66aIXf8GME4jUUZjxZ3Qew4NA7BsNw/fWdHllh+UnKOEfzFyp
OsPpFoRhppa4fPg8A7p9tVjpRimO2JaZ9esdkC55YWsqaBnTvgqrAyLK+e81voLfv1tF/3AA2Wh6
JfZiQeye8PpiIguQ3dZ5BOvTTt/nVUpZ5BEXD2lVIhxdpoQcFcCC/Z7imyG/4bQsXe5VDyp/esdt
DjKylqZRhExES6jGqc8BO1fL5HT82vf3SWDKIzwt0GwABrYzoXx+2Xrm6hl3ULDZkMtiMG4JaLs5
w3FHNWg+NLGXtb3E/zylSMDnxcJTuH+rVtQ2Xe9B5NmQyPQ1BAn14GWN3rJ18vUA+1/TNTwwx4XX
b8s2PttR7s2sroeU8jo2OeGowdl0APKzJ5R0nK8Sz1eoLio0PWxiKjDwhHHTVkD4a8V27WEW8Z4A
UD4F8TL879JObMW3KNjQY+5EI886qwAUUPws0Wm1NUaR06hnF3pme5TGtlaRlb8g1Tdr9IqkVmOQ
QE6Y9S54sD7pvh1kMnDlqGiH5zzq1k3qu7vV/NV6/Gb+avnYr32vY752QJCkbZs/yuZ9gEoZROFL
olmVGw9lRjcFq/tdl1BBGxr4464/14pL1xx8WMz9dOTQxZBWyNS0/MzNjqBHLxes8J9kiVplLEBs
rafMz1eIfoqr5uvz1t7gUvVrstA78SURKLzcZpZKOV2kVwsQaougHPmmoKuspfksZkxHA7Ee6vf/
lBVabfHErMZK8w/LHgGgo5lGsMC11ckpTmvxBLLUH64sNK7a39yE2bhpdm+EaFzmXUP+16MpTf0x
v5IugMx/uy5/ugEqQVg76rcE/1KbyI868xq4ASO/qE6RJRx9LKquKXY80WeKgR12LgaOwD2NnUnc
EtdHuxnEloRKg2NUHG0CIXaJUuoQGRupNcPQoJD6mvrjp2lCDQ7ElKBNVLq1MQSrjJPk2Ol+0kef
982bOcrWsUvOqslKipEtpHnkydE3Z3IB3HfcfeIEzxP29td5Xn2m6qCJUjd40hLkV7iKJpgqvqlo
gOvEM7q6pgdXUlk2HednrI+do44a4swK1khR3Pf66TPj1dek4Ed5Nb5BmxGNagLrD3+tHPD7bljB
gwNY33jM6dN/1h7CqG+uPeEb+BGW+mAEmpiWruKDMc2US87yhvUalHpwpONsNsLXv9Me4Z96oxzf
06xBEnXckWOgKJv5KF7vzT7rrCr3Et1Wnl0Vgeet2RIRuOafekbMcNEUufy3bOQ51h5x6I3rxwEf
tHPjINrx5yAHQHoUg36SjeA44DoZImwd/QjNTx7Zh3XyRiH7D/romqotg8EKvn4M1yXCVuS71A9t
WTsLgnnp95kZ99Mck5C57tqJsPsXjCzdnA96Gd9lr4dLgACIXoj4sfDJCbu1Wga0Dh3i1UAYNJ0F
S//4/tdIq0B3kEM4r9L4FkQyJZivjqCeCIXEIrIXE+HAun52xjy4HJVf5KI3gFV5b3h0JNRw0og4
5bLyQ1uLvGY8M3nVmG/w8M7ZqKiF3VOTub5Yl7u2qBFfFxdVyd3iVcQamNrOJW3bCDWckIflhHQ4
RSj8DDeQ/ShtNXC8aeqOvmlyaRV+6WvMNCOCcRpMeuUTpSk4dv7SEpdkZmjB+XlaOIfaTrDU7dye
htUp785mrOV4TLRHdmjDlA+d4CtnAszRxAKAMebydL5P2m3/QsVbHoXc1OKKDq5YFkhTmJzRaHcC
+4FvmEhKhPMBNIaSAYvDxH9CDQyHZXb7ZaG94ixIQSLy9UfUqLkJAXpH3BYZOQwXRBeZ/c3yIXGS
3w8pLc98QUKH4V+exAXXvspCzLPIK2FW6Y/EATQAgF9uNmHRAM7QDUXz80CAbyTjLmd35xkxiA8W
eJ2yzhdFcsf75dFH9AY7+VDC62ZTpaMtSMAEO8/WVGbyYvwUKbpinufvWwmFmCCSeb1GQ2DLQtcy
RmnVblyX2+zNK1JIJFW8E3+UFo0YkXS8p4Hyz7a3M5APZxDXX+q8PPE4K/JJgXvjsyiPVNLp+2wE
zntr07Z+eSkX7sYWqdz+UWovP6VC7NqW3Ng2nS8v0+NpXxIDqdHssdNXIJ6wW5IW7qR/ULB8b5D9
WpGkEUPIE3gZaW+GXjN7534UoK+5xPyjMd4DgZk/4DGNv+AM+3G+bcZ4Lztlt3yhNpMUm4E+ha2t
/xH8HfalQjuSyyraa1rKzfihQ+dau+zwKJNEE8ywQ2Yy2h0nyiY5l6Bn+5mJM2xLcZc4eW4l4XCr
koKM4WYrolJTaF9rq1NG87E3YuXavaDpkVEGTW+ltU7F5jhaF0vjhs8cdwxDwLIVF9OMl+VRpZGJ
QRlusk5fc2AKyAKM8fWGgQTpt/cBXlg9pcrB1Nxvc+jOsinwuenntTudTS2WDrIkyOfTxkSaK3vc
o/PCjOReQypAC4CI2Xcc/M264+WBmxQCo2Ernnkqm0TUOnbDQeiAm+ff8TGlHrO1P25svAnqJn9I
w4MQgFddcFEw5L+IIyDgqKoF/k/KtC6uBv08fxzUF442pGcqV4H258/+kbCQ9ULVDpnQcsYrIoEu
tojueElnjIaW6yFy+15e4x1b/01sSJeaP5lm102SXOfXrKkBVrOzH/2i10KwjifvMdT0nt7vsDjf
ydS3YPOp1Xh7xBbLEsSfO0qelbGEJ07Ij4DUyHxk/fCL84gCPX0bcJHlTeMnhIKFNMVTZ4b3K6lK
gAuFXpUmjuzXpgL0St6ePl/PzdEGE0ie1uSOuL/DGlNoViQorqYdturwFtsvvutUs3YJb63CXJJ7
cwt1KRQqlqHEW1onuUmkiXgqcEPravWkQIqrLbG6yAIPAv7dwKOQlW6ntFc8DJOSQTjUIVBYL/Ly
TDC9BSGKoRvDxSYi/dyS+OZAwetNKm3ZcSNB3Y1kHboqmMn+3jeIT7/V4dsl+/DlRXaOFhFOttAi
ECZ5nNPuwsz5TqdHL6ab9zs3PHXw1hf/s7De1M+gFCNyEuZQTL49pwgbH9j9Ke04Hz6e7PCLsMKk
iVnXgqYgtt6PqPOJLsDEXDLr6ir6GBpK8+DfDIzWEnBh0PYsNWHSb8aQOt4Cl5oSh8k7ECnHXjaG
ux+CVJ0GpYHqvK5/hMFdvXmXV29XRJT1ihS2O16jZh8zOETzFmp6UA3ilq0N6tNVq/ZlirnUqnow
wfvppxhiw/ebSXe4AlWfHbJ3f67GRIKM4EXcrIoF/R9g08l5upkeKDa8XQRnpvT+TSXAv4yiXr21
A+L26FRUrydibuy4y/Ko2TEMAdtabR9uwErj2u0Kt4ipitHPuswwajEUZM3TbasqgjITE8HVZNej
BN+Od/msbUwugdkT6MxFxA/4ncuSqQ1n5VrYgPHKg6xj2cpuOQ8z3TyxNOlh3Y2Ye9TkVpBEeJR5
eC4buNP/9pQVujiG7iJdd1wV4HkNxkiekpM2OrTUVNu31DNQopdQROVjuO85KFWUY7S9V9I1C9tr
7Jhi/ZF5oWmwvzcGyYlBjSEuhY3Ggbt/mu5yeFUO8TvsU8qfJxaSF9HHBPXa+Z+C9KNnuc1D2pNn
F1MvufB+8aFTTcW0bYmD+PW/YQ3OeLth8sNN9Tg6DCKp/3ZtjSQIh2YU7R9hV2KASW6iP5/RcC7y
AW5vwWrmCrkBSI0nvpY3mDhSE62MhkhGhyp4ZaZvZu1Dx7+66S3/3o0W5FoZWDXqNx9a24Xm4lwM
5voRoqUK7MLrivItGz2Ea7hcYCLGab1/P3/J27ryEQdp3Yc5BETm+5Xi2Dy74PDJ7vM8jY9nqwIz
+njxtIF/UyhMPucOcNliA3mBJhXCQDWDFXhAEQrHrvOK0bNBXyblOfrWIxXVD9u9pMW3iUxGnZsV
IX8pnr1zo4eC8Nv0duM9wTYxL9Q1h81w1HWQPuBD9/4sa+DML8brJHOs1n5xwVoXI/SoL//h+d9g
Jfz7jwn9iZruL0XmSDWAzUFbxJ232Lf8bkI8n03Rq/LEVQ//ZlAesmIjzDjjHt5cwwaHtr4ixYWq
I0/EFFPWNU8vUK8eYTv3JzR3c7b+tvedvCAtfXPlwunbAc4GwzIZCly1F92x39zAdk5b3keZv3EH
GPuhL7RuHysztjiLJTI1Idcc0wrFXRaFs/g8HMmxNCiAS5zdFFoFibH9elnH0RWNu/rz4HBw4/iz
x/39VH678Gxej6ppmFGljyBAglE35pIJts8wFINRAdg2XmUR2rVIQvIIZ+1IkLqPKZIoM4HbMq9B
X0kaQa8SWa08UmhSvsu8+WBJj7VBBfc+pIKef51g7uNrYOV53mLm/IkCld+MP/NOas1Ral2MpgMn
wfNSxkMyxASIW/K2TENGDuH7TUA3DDe/Z/pJfquqqaTRZyPO1IezNC9mvic1O6ABMmA7Btf1fz2Y
TKiOZgeTlP/7nFD9rZsgsqkVgPLsr3ucQMkTUMmFb+8gYvil22pj/enFKkgPFnXmn8ACVwgddaA6
LF5KIQ4c1kPp88VQ7n09z0ufcHN3HeOVvcBOs7xAB1AJCsX9jZiLduBnaPdcu8wbvavrCNKE41Gy
Y5Jrw9zxju4G7j2mFjin4tyFixeOdKwn2VXrmxo2fXyHrCB8XxwyGNP2IH4TrDiMG/OW6I5oVrxF
dUwQzAaNEtaMYSxh76p/FE01nLH1EJSjkt55zUCIkR5jhDsei86pe6KjKoIirFU6QbrK3qu6fXHr
+gmivgbFjkEOnkwKTQJsSCYSVBEyE45oH/oVHn2Ci/Ux3BIMzM3Vm4sKFrymB/S8LaI2+6aD/Tmo
eU+9kZiq5GbwmZFY60GGwJpzqdELOyG1ipfynls1JaDtSBYiL7IJL5S+HrPVDybyZw3c4wZCSAXL
a683oVVQSsYiK1jBiT0+u8SWEHC3EbmDtgt7YiVcUZ31FcP3ojGAcoirmP4y5tCjg5vwlJWFfRtk
RoblTC6PtkwKnCpCSApC4r5KwWEmqA0O5fCdamDPgljrC58IKfhkg5F/ro+K7qUw4OSU/seJUnu1
Ks0W7PprS6kLchkRumqgYVnyuSgyKmKD74XPbk7pwFdGs6AGtnbpuhqT7jmg29dr7Pl36QCxOwdQ
Y75hfQ2Jp/yMdESJW7j41spit4jFyv9q6i6x/q/abOWqbYTo5yu46Yu7IEPedwt0fD/AH0i/Hx9e
Wn5bmxHnNVG+qAZVtSfy2Lrzq5LzSt7usVIVp1wJGu23BdWfDjMEGHUS/AHdFVO2Prs5TysNHV5S
ODru1UjxBy/FOy5mrK3mXPhB+MuCGtMtjN1b+nezFX6tSjljHxoVc/aQXcFkhW0Wua4A1ajitLph
TO1mTmZpjTMIw5gQOpzFaSnjBMJJzR3FWOKMPMSfkcgw9A1YvRpB4XCEZs0BXMi0HswUA4z6zo6m
jbZe0zgYHAiOhmH0heo68IcVF0cayEGxlIpwUKU6Qbzab/aiWtY7ZzKmLXjc9lFalgzFYo8/+OPk
OBdkZJjNpy+kJAshX/sMeJzrAVMLspphIwKspNwGnOOjv2MonGx27ROtcEzkgoOpEo1GO2NoCt6q
yC60sSPyceuarigxMIL8ITZ7TtdUuVf9Lv9SoLtZtVUIxTi1R4+b+HEUnkCOqKBV9vW/8FRXNbqp
h9Amtk8bjhTXp8se7AtUzGXBbqCuoLXQfU4WQW8OSApcdsaDOyMTgRrguBOLob0cZdSYD8Rcva97
RsrTWt4BvCcSXWutZAz8cGnKwlH7IzU7GBMmWRiY3Fn1kVtYe8GGcf2mQIWWCMcEvik0enInSjQc
SXsU/lZZ/2Cw7s7hYuM8kNEYNRcVAYuQL6PDt6HsAKDL+CYPW7fvGRCnhV0o1HmONzomfKjU5JGc
jZ5xil11UIW3jzfDQ78ECbfH91XwsODNMtAK58B7EhVrpigYOg87VKIt/hABAeR6sSkoOawbP1sZ
aX/KCWUcDFqeN5LbgoWf6iHz8chGPNSb+RT2a59csV7SSRtf5Xu4vrxfRrrAb6979kskYEH1TnUV
xwzG55XuBjK8OydIajeTYI76hvy2eJUtNXnYuprW16+G+tFsT1ZEHDtg+npohm6Lu2/DZhJ8csad
OxOTe5jbiqVOOmiPdI8+ee2MB4VZRNFgdpMa6VwFfVfqpkycT0SGOdE8ldUE+lCwgf3v8BFgTorx
2/QxIWYGqHE9tHcPhzLyqGbrku0gtyCXUHBtSbhRZEab68gQgFFaxBhJ5NUQl9zaFzVWufw6Lq0M
MYLQC/4McQhxZ9hQqqBv0NZoJ2u5DWBIM/HjUJKwpeKWBDX1pWEJdeeftqjlGr0HftASjwFTWPvQ
qfoVKRhtwEDRGiGI4hEJrUag44np4wER5EXNrQDTxQlYtYFSLIvpFsitp8Tq3XqZ7h5UmwBcChUY
6PyKr91b/Aj81TF46OxC1ZM7VYpHwBHQDpXMVvRMLHzSq8SvobZKq/hZz7jS0ZaXzZIHtoXejW2T
s/92Lr8mZKaDLBFk19FaQWOII3yw8lvS1UuH59CKpF+JBRHoa/FGTTUv3ArIdFwT/zuu2ZEZAS2q
iDgLbrc2uygEitVrFM0UII6x3fjCPcT08dnARPqh553We9S8QBafuImiK1JCg8tISlVwwEOi3wIl
edFL0dqYzD3sEittxYStG+Tn8akLw8kgy6QGIzdzziGtuu22fleeOYSObES3q52v6N3KAvx9vPsL
E2Q5hogDKJ8Y56HKkcwnUnRHaasS8O8rVp6/sC/6YlUNcHj8Hcrawou4+rc9/C9JgAL9ipmLb+PY
agfdq25H/qZV/tom6DZ+YRAiegiqhWIU7Lxe4U6L3DE6gwEg+HYD7nPWHnieJTYRLdO7T/ApI7lF
Mm9eolila91Jt+ZoJ/TC9SsJsvCfpGPJzZ7ALa5uYnDeITKTOy4LzID2NbLjN4jE3MYdgR+60IyE
oE6l+TiY567ljun5FIPFdZ1Sdf+c49/oLmbAmgTc2+29ovO/P/FDsKAUno+qwd/Lnz8LJVrEH3pC
WO6s9enlCVVhefiKuVnkJ68lmVm/pVhihN79UFKdVDRXBIzUGsWL3u4tlqjsYAZVCdVzRpcNc8zp
XJmxnfX0avPDrV0Zjzyd8P13/T3Yao45PyT2Qu3xnUwQhSC+B3z0mscK7YmKZJNr1z7sCStf5EkT
BIYgbPrB+8kG5mm24eIbNqiLiIgli1LvUARXHYiw/bZZyjBxathFr8W7vmU/WjxlM0COrvDPlO+3
Js+3h2fqom+HSb96zj1gC58F7m7dI43FyUFaVEivr8L4aPedgT001IcKBCa25b5OAWH8r02bSoF4
IKSSYhrxdFz3Bn1wl0zBe2TJxMMuNPuqy3BJFov+EvHKUpB8Vshuk6KnMbxGEveslfq2OOpUKHs1
KdEdRxX/iQOXolhaop/orK2Bv3FPNttaNqhmJwI7bxqbN1pPhutcBZADajiDqGJ0GWOr5sOKZD/9
VEPckw7dbdXoiCvAzX7zMKgOpIrknp5iQAK2VvZ30pj9xDqdeE5P30dZvskPq8Kj57hJkuJWM8ii
RR9KmbGcoJRN/R8LzHdgfWpcyHpvDaltiM5ZKtQU03hIk90NqXFWVf0xOVONLuMdf13JR8PZ/AS+
RT7X9VP7mYWG5Fk8B1VP359go+jY8NLBbA9vnjyVyWnNFastEl9Yle0zr1IN7Fcm8GV5ToUf0K88
cc43Ovz4WxrNGqIrHsK8WMhhCO8kkMg+bkVDERVA3AcaED++2UjJNq12oSYN01nVSwKqV5mjo5uu
MBgovRXIHe+sL51pLZTGh1GYDkPITQQZ3yHJsqakcOrvZpbyxlyTWBt0x5ucWGSVVfZaFDwFk5Gp
f8Caa4ECLE6HqqXsiRFPZTcGx4pHaAzrCDaMrZhaXOuz6ZlrA26qqYa5yLWyc18scq4LluG1R2qo
M1yJW2PaEgBV7wVwjVQOlW9ZfKGZJyZxWCpuR/bLeVrYJOiuxoLjyLd3vdqEKzHDW6eN5mvbhahL
XYDw77FFSFoCnzbULWGFiJTC3xd2PTCgBlhmdOhvqc1t7TUzf76LyL6lISzeaGrA2K4SLWn4kl7m
uylXHRON7qMlfQcYClwEys415yhZIoMrIddRvpqeWvFffLMJMWHBtK4/A/2PDdfssy9LGBC/esAG
2ygEsMvIjikDhL927bSidEc3Iq3aneTYU8zp4IMrdH9HrlGQY6RSDuM4HWAmY83skCaXiLxUpDBF
eZa5CL4axufm4BVCkZfpn3Spe+cg76Hk6hN1Pm9bdLw0DdOflKs1gitNw6V04ycWSu2FHIRUB1e2
lEaG+n7/o35sH1gMcsknxjwBXTlwMaIBGVmHHE754H5qWsZHaY02dAgSNrHo1jlDe5klmF+EyPc3
RjgUohrvDhBOpRwUuqYcweCMZS9U/VxYe2FiZUxJAwtQTT96AD7yuYBKRTFAPHoEzPWeUeHOmGlB
Bd0ghewE53WEU7b0F1j524eV8PF3nj/wN/v/pcPh174fBZuLmEIuIBNm3Ef/ntQNLtR1P44ljZFO
3YauQZ3btH+byUAsmXDvkNzBzOT5qdiTZ0ueQu/dpqZnH+r/ajsRmv5BcMJxcfUhQksyum+JMPgd
NJOdPFtUq4LifX7df4WrI6Aq59LgGjS8qblWysPv9eCk48eCIIeac0ZojE2hJcPqyGIJiozt25h2
0ziI+hNcq1hfUDReBQLes/XjmNc4STFWxFLDgazLMu9MZqIAWu+BbwUJKfGjus7XyObyscpiLHwF
M9bxfFyEWKy4kz6ZXkmJiTOYPVN0dYiNL+9GaY4k0DeLbOEsrQdKGu84497L0OGQ8fYPGxpagvhL
1mV6tUsXdvNRYI7EJXhcBU75FlfJir0kcBZKncXgpeBH2YrX5nry5xiYw60xDC30+E+YT7yR5dlm
NHzn4q3Oa6kMDgqNzvbVRdKUe/dVLqTR0Mz+6riHA1c9JWE/DJrIk8m7m0b/4yoWZVEOhCFV0bVe
h9ir8ruYM0Uga2diZVZ/bbAnuIG4rWMMFvVaem9iH5at81sVKKfWVwnheo3j+atzPVoSem5CP3PD
qiTHPv69hadGJ+cileBwD98ji+j+DmpWAICgRmlb68LNBoIVdBO3kcI6CxgqN9i5vT77kJduYMvB
K6ByytWRHvV7mcvCOpdaOkuQxIlYJSe12Q4+h3TXNYFm5OuomPfH0+SJ2xZaKzgcrNcdUu9hlySw
rkEoapY3+x8TbeuV/UP8DFt130nVSzKbSdRrXHtWZP338Qy4vTiNuQZ51Cjki+CRnOdV0zl/asaA
xxf6tQiKXPuXMr9PQUO9AB9E5t/rSYjK8NDTWq19RrRyMqvRGGb1D82Yjy/nOlUX8qDmuPf6pOar
AC54GaBwx7wTlwPfAcZ55nqs9pM8ThFx7nfHA7xy4bYblELhD/7aCxVHkOoifaTfUoR5+rNd3ovr
aLbmPSjezshzXyMvVIaix91GSD+6szADvp+occuvJmA6p2YiwxmGSDa/tgE5YZFSj+Fx8yGOPsTD
KjNl4tGu5dnZdBL54j1KRS27nOVz/9mFi3w2PS8OcMTd9cVEBgivAENDcIwQJ79GJFuQXf7fUq9k
o2vHvKNmu52qxsy6tA+JsFMiec3vF8o0cdZ8V+V9Yv1IeXytRpwUe+njhTf7E6V+ljGhCa0O1ir6
g6BXm+dZPUh/k1JwS7P5sW2vDKYFKZBYXsXJDfnJZ7Rq3jo/jCqeqKEenb3zW6L5A5jy4U4dek+Q
drLypEZ0PlWgcctXlFWoaVXeLfrfEmLK68WnqKq9w9LQY6HnIIWvvV/7QAvQB4QLLSHamjE43vCg
SQ64TJSMxgTibJHeZthQFdwGjUWNA37t+s/ZEyhWVM4bzrsWApFv/HwodGyBjQzQyHhnuaRht1Fv
DvhgJtueHnbrUyJkkg2CzaMYB3QBqGGvIVcGxMMluAv0FL/JvBVj3spZiu+8SFzl9MVJf922foB3
8QhEO3lbb+DlUis/ygd40WTpTo74EqbJLgUGJ3Fj81Yy2SyjIZ6ozO4fy/qAOflPAieNsJPJhVDG
D6fqz/dkT050yjvcCq4lEo1nPhlvYmq4Tz8Qexb6Br1ueKQstHqlVDED/CoqOo1SKaMgNwdXzZwc
dk6HKWIPBKkt6PDl9rH39TIk5yAMDXe51zSWBMFYc2MOoAxm3Z+M3huTjbm8293N4IyCTSeP1b99
YPpeu+85MnXLkcAsqqFo6OOaL9IunyigEb7ptFnRoexFkpxy+vgRCYqntaPQ7PTfLjfeEnvO+q+/
VrbJrahSUISjHFyOVMHr8kD13j168Ur10FK1N2OQtZq+7Bps+n3LpLubEGoT9Q78mUxbTXJ3st2R
AkMmvMUsU40C2MILktjWRbcas0SF+v5BL27ic1sbObm+hTFHlI4N03hro6QMqO5zmfBajoo41fS4
Q2Nsa22Z0fyPCxEfqClGsYCOqGWuQakZbafxAKavocx+TF1YALUdfGIfUjyqkB1xxmHhHSjsqK7x
xhCdlL7cYZtSaWNHaKrHFYs6EwOV81TUafxZAm8mchJ5xg98PLcuPJhdw7BdT30rIY7L6e+4BJWk
swEVzeVdNB1tfMCudH5TuBXJPgPAMUzr1tCTmfZhRCJ9EAs4rhU4RioNzd+uk7yyQ/utxlP3M6om
66D87YdOK2o6aBTERj8uIyU0ZySx7ri69hkZ/6ZhetYzF8VrpdkdX9PvAdzMcRQiUyr911DTkmmG
SHzG5+A9vqkxe1SYCWc4uZFb9GzyCcx4jHhncEpIY2RasP3nNmxQBki9TFJVBAQ2cBnhmgm/nYU6
0ZrSz85RiwinCBei3pQ/iA73JCBPDL5aFeVvflLzo0g6YQ+aUx186Lfn6RFvzgrz9nTKsKEV/UTc
6VtxyvPRa2RfQMqn9ajhsMh27qBTmA1MfZUx6Pgnn3ojVGCLYTwroRy4czIcRLlhznhkDJ827PAB
w2YRszQK7YSA7l1EQ/yi0gBT9B06YLu/WFH1Yig8Bh4Q6K5ze261dSARUrnPvde0Q4ttx1LHjQmf
umVJEqqoiazt67RGcUVyOAqdpyReYNqoIZYamdLoRA1vEnFMC3J3dy1oAXcU9LHTwioONa5TVczw
SeWYC7Kef+QIqyyMrGSf0Lu3vIjj9KcDEdit9Y0jkhc94TKZDG8TNCHfPcV3F8JPI8oC16n2+FVn
FEBCWBatpJgfJA1BaEOj0mPXS5k22nI1A/QQwHIOcR+p49dreHHpahB693OoLL1zm1pCqbSc0N03
2lWO6nWyb2KQcBNNAQp7jyXfcWuKMCnu/my5rcDPgoc6XgQfGmeNVyQZz3I9PtcJY/T58q8amWGw
8AmErMhzozzmQNyfk8TIJ9HPRueN7g+f+6ygTMLMeXAX344mPW3v9dJmNyxzspObHZAblkaCa5JQ
u37b4RxCLlf6eQm3XeiQ+zvvrvJEtlR23rZlQPgJyw8Ct8uDszkBbKu0nCYMo0YoJhooTCvRyl+c
D4CNnLDGsvL4j2KI0bLmgGHpC9DgDJjmzZUufFL1vRS3Svhh9LVVGVW2nbHa/XPHMZH/dLnN6MfY
WY5IfIxJrNQpDvX2iOHCE7Z9Owowv06o3pSsDtccFrXl0SfirRW6absw8Q5eFFH2MYZGg9+ow+/w
0EXL/CGSXK6AKU5o5gwIDRkkrUkPbuf3TmE6eupWqfVdQc5gb+1rksZsNJN8HLivDRHV7kOfY+DL
LkkWRatd2bqIm3ymgF583iI+Uo4EciXxyxzXGGyjWUxr5xWYd1U6r59ZmjQZahBfmWgy7fTLhn9j
AytQi1K254zmQbN74KkO5LgSuqeyz4mLhvap79QYv8affbQkbH5+W2/j0e5gBvwIDOM8s5/lMNhI
y/GS0xAhdxw+IHBbl8HY5v+3McUdKWFuIIA03PlvoRxP4QY3hvVDmI4U5dzIqId83wEnMqwaeAh0
EKkgAY6XOeqZWdYiv0iQ/dLm/gai4oK+C1w43XamqohO4Jdtm8zUq5732RWc79ODjMeo4JmlGwv/
wfjRGpA3GkxGZM1u/upb+CVzHIXjh6WZjYh8Lh1uz7U46AtD1bZJXPUsa3N8swDM6uZk7SvhqSNJ
udggKbMpgYpmMHqWP4nCrlPmwjJUpSRTx3fWMoRmu8PGH4Xs7gH8YaIjJ9JYhxgq93D0PXiOk0Eb
vE7I1Ay4krBztWFN3Bftvy5f9cusfYbJU4FEtEnNV8VyyfBjSsZY/7QWiaDSraNaJmB4H2HvSkew
OmheGkgCuraeA69yS89pqqZRRHu24nr5Wms4628p21vmxatdNGFXXw3RFUlPjYWk/aHm7feN1c/M
ki8z5w7wMo4AHC5JQv9VLIN0ojw4PZIzDCw17XJEpuO2VUPsOD+l3l5w3LYZQ5g8/M+V0JStvcK+
3IGec3jMDSoVM+Q3OaxHiTjJEC15mGHnZDXgCXsgBLIMS5uS3MlHrL49Bm1kW+kdNaRwGvW9fRrC
GdOygUPMnyf0GLd3fw3sawLEkGQvn/SMFGsRo2vC9m85NeyYsLrVScLeIYZSIXW73XKR/+50CtpP
AK1IE7DQf1bXS7pq8RbiPzuGEuabPc6Cthp6QPwTiRmstXzqUIipRpTa3bg89kYzOnBFkZ5TAJ3U
wpdBhdm0WSp96Ou1k7a2B5/4odXvkCqhHPxM9CvF50eIjDCCxBCQzncukH/XFf7Fk057RlbXqIPp
Io1ok/5slqTs6Y9cGubhHqKskeax80Nkf9qk6GQGqVKm85gHvvUuqjXEKETQjgc/y2Ul1gib6DnY
+FrxP7ERyryNLU8ZAMoGG4qNJ7994zzb0WTN1TjdIbAOyTLnyYKaC+PIU0Rb3MrAPTuTcd6TLrwa
MIU+zmXLtvHUBJeunK4p6sWSKD94YDeXk8BXxC6ZZla1R3LYaC61yZyLal5SlnjGwldtfcMWSbb7
5NAcFysh31KAkrkmEoh/oI2zKZtxj+qsW1TmVU5LQMBqqXt6p0XH2yRu78g3edS+OrUD3YcXCE5H
4YepRzUIdNNeMtWQbPAXT9qQE+v/xz5ki1InfrWVKkSCxlWKY+TyhnGlFSMKHODcN4OdVVtab3+V
VNI9/Qy+MtoMpKCPW8iTaH0/L49Cqo8z6vU/UEWgTAl1JAo85rG8LBSQttomj/rRb44Bg+s8yF4H
QgBiY5Pc3kl8gMAcczC7E11b58EwWkoUaiwpMWs3vA19IzPMqRARgM/1MI6odzr025rB58G36Il7
Ht8U2cVSIgEWqNeA3S+67Q4aCR7OMYIEb84OhPQ7kblVuxUpfgmid7y53dL6vA1iThYlusZGqcVT
6q0qk6J8r/XzH7rWnrAGPL6V5UxbUf4Kwbp+x0YRG/E1N/RoXq92qWIfSC02yH7Acmjp+yQ3uE70
oQlHMKQwpM0HtuQt3TtQES5cU0xJbAZuidb8f+wTCmmyHkPKhOPEEqh6pmOWAm1txK80Qk1VeHxU
GoqY/zqaGC9u49Q5fNcbgI9FnZSKXFxtjLZu/gkMhoZHiG7LmUe4GSJB1JrLg3Hb6nAc8ZU74Be+
tjkLUwM0l2nzMFCusTdF7L8IgOt7ggPWS3RV/6Y7454Z57qole+6qsByFwClVnSoWpxk5XiEDlpM
9fBy6gO0zbwWuymdIaD85e1P6FaHmq+edpGRMH+eltvW7UqN4DB+mAg9441GlOxhldJcivtzjBoh
ggP7m2AKQel5ZchS18DdtzSS+bOxl5r6YGPFQOgTY+1zQhRebs4KDk4DiM6/9bD57CmMX5+u560M
G3BjTkzzQfWOc/IAGA/0wVSOV+tnmblMga1/mfNP9uvalbuPYsoIUBm8vO8w14r4sbCyLB6J1S9Z
YEcMU6rNFOQY6zQh2/Ym/cg+6vfHosSdfm6zgVq4c5bxClVCv4ChuoKh9sgOJVoj0LtbZA3AH22l
2+eaPqxXCknO30onCT3TMRN+sSfQUvnH9S9wimSF6m1Wxq0SbooLoy3XDJBUvsfS2dz4T7pAj8UP
CjXM3ujhU4FJIqTecHDwJstngFcL+sF8hD0sC5PbJaE8ffsKqMl30qI7tz+cvXuvDF2rd0Rx+RU2
PObzH/g1Ihsie5Vhl5h9KY0TZFVqf2XtJAzbRKemei/YpcycfjG62OBnQlSiyGN/eUrYQigBJm29
58RS9GgIb4U7SZRwUFDcNSNMHwz/Gc3Pr+JqXUkOGu5cMcbh2Qsz9n4O3QHwcOtON7FKX5kCztih
DmMX4JiQgqVkLkWWJXU+Yuu5iQrMN48BkTlfYEaUyZuY3hw/7srWFVZa45r+scca1W4t3CYewvss
/UelQzZSHPScKc9XDUVmp+U/nABy/mHtbCUH1tN9UPkPQSgbskTrPPhpHIXwc4QNsKd6xI/iHOBJ
JpfOtEl1WHXqKXFXK3IosMSZAazV+nF8p7uzY6nCesVwOR01BOq1iZPGrRu1RyeNtQsVEK1K3wUk
BD5xNWtn3ArmwIoFEBYnACD5QgmZh+utiFMteK2RO9pO96uyT/SnEjwgTChjUitURie+Q4a2Ohre
kHGc7gF1QU77GI880h6TxMRnKS0NXiS40VrJ4Ib2r5Sxz4nhJ560khAh3eQz36ptX7uWjwXMhVNZ
UaNVgMtG/u//VRlLQIkFUW/XBI5WmTWJ6lb9RbNU1Wmz7g1OhH6e1seMqmERxzXdfFEbg5OaYj7n
lh2Rmi26NpogJuziHToYeB5sRYlOAZV3HRWO6NCexrz2cnFNJ6eBnPxSdxcwAuG0//gfa04o2r91
FbYXfty5Meu5aHA24gqa0Ly/IqSa6nl7k+3JIG6Ly6eFp5zdrUQm8RJcky36GhehA1Vh+cCqjnNI
USjSiyDGHn2zG7B1bMK6ztTqmdpkeQ8pJda5q1uUXtvVbPIIx5m43d5eklnnOs5eZPMFwzkTYiaD
/DVqZXZWnFv97cXX+h7u4OLuNj5KG5u4AfC5G1V3jTdTFxRhIWe4rlGGInk57BZNAfuwbIZqS+yH
Zzy+n2DLPeIfYv4irm4jzSAs5TTNMY2b8vHfzUS+HpG3pmfpro9qulBS80qbOB65AURofkUC82Tp
Exti3auzfODKRYl/JYdXR0MU108nFN21inVPfoAXqnulnX+UsAcsHU+pG0Lpof26lRGY54HFqRW1
cZygU2BMhYzM/M4gTzkE++OaG1zTlXOXQ0JMUFBztHSizvOVHk/ZiQNR7MnjBCObdgVVHgJeNAJ2
MzzUXLaOwCt8a083NfJJFc9x6LTxky9XGX5vzRqG/nmXhPGFU1LqC1x6BethLWH3ms/b//xtQyMb
Ge6pHgO3LYMivnIf3odxDay1bTtx46Q0kpByp61UBGijEtyptn7Uhe7tXJFXTpxmXikWrMckxlUE
SOAvUpNUcnFGwwGDUGNIHh+1HhRtc9VqtwljakDR0XIHADE3f/Ljp1KgyrqlK0XJbozX6Z5XnoB3
f+5kxHznKILeY3mVDcz93uic/2PCk5fUxR5tY1Teh+caBa5ktC8mdMCT3XvES2a6udbDAglGQxXF
nmrIxHFFHDfT6PwL3nWnRFyBlX8X3dU697TSuSQbfJ1layIqyuQvW10TKfK2ds38VOQcI4KAhW8c
q7DXMPuSk+TsBDGpQ1Qz/50Ko9AzWId/tyXlJLx2ZbFl++QyXenk4sRxMgur2YEPSgGQu143o8u4
jb90z6ihlypOtuJTT37HPrRg4fAB9EYdrWx6MOlW6rFs4qlJTXkPSuegHNLf3Vg5jRbrPqn5nrGr
akBAilBFn2x4F305dgfAcBqQuZ4cQl43OkekcOGrO/53kMvP0xbd2Jnk38F1JVosWbHlhovnOrjv
qqFEJtb3c9OJx9tuHhdSHI/6fIjYeF5/CmUMQOjDgwHzq25sMZKInX840tDIRrGMTsWmqP5GcMmi
/cxzlg5aj9NhBbiVHVO5gY05p3tkz3bXjDQSrE0q82JTVgPSPHaQYsgWj1HHlXOJYVhPn4wUGmnA
1iBLYMWM6FllG+Ex9Ni9GvJ0ecDul5pMcPE4kVO1q5llRyBec3J2pt2SKy0ayy2PRHPU0bKy7uHv
+8CwxKREkyWTee639HCa4CCt2iZI8CD+lLbpS0zv0dtHrSyUUmzuGPHJZ9SHcWYyF8dlzQ5Fns/c
irWIpGywqBUHs7/tnE73yObDqWs8p5sLYewz5FF6iRQcrMUHSe1/1nUa/fKrtUb1PvW6sjvakDXo
4AZ4rNrF9np6pbGVVNPzePLo+hYjnnXQEd+9tKROEP7ZzpwRSPyHRjAHzV/AE0VV3wzhcKWj/fZB
ZR0OSVd/wvmulTefiy+i7HEDUHOWa4/JHaZdaqxVxIbDbNDjRP5bg8t9/DGQbnsBP+a4JwS60d36
eR3H8xhHJuidhMPYsGSlbhtX36PdZoXJflevxSs8fKPEy7V+APUlHdNg7OSNITgM/DmH/XLa+gVv
xQ3J8O0hY0hJV2EAD6WD/gQwhZPLSf7NfSaSCKUIyMK2SXXqYawc6i9uMoDzAtxc8dNjQ3LcJ0Fu
I3Es6UoSVGOY3DHOgEq/0TiwAFZ7RyIlWrTDzOPkDiS1EDQRgB/8Uumj2EB2sJamkrteHxsY/u0u
eZGRurtqF/SdYdrRxbGOCqVFLPei1kJA4RapERN/fQkalU/XCO2S09GrVxRYwNNSdraXaFf1u2xC
KQCOlsmUYlLqUcluzSgq80MO6xGo4t17lG7yxPnHeSpDknQ0w+qMWZTntgfh8/k+S8UsilfKE2ZM
Su96MOMWgBz7CimgS4VqaDzlPckl+XSedvQCcPNtFCcZmrsWX9uUSSsSVAc/bZKm1dObL682EO+O
w5VQsHGz5aA3dnYVg+sI70RH1XvqvlIz0oXP0sLzQ1vR0SCdOle6zAGi6EupojO/oPKpPoIpazfG
gQozpqaW9DA2lk9wnqCaB9JlLrz20/SQStPNlDUvJCWAVfIuNI8SQmNPAm0EgIrrEEfSXYU3iBXh
ipR+WgVdqE0Ewbdul0nMcOzjsTpCeGJGKZgqK1pcZ0rEl3kfXRkmv5Ep5GIaHf+wYPbEKZD/ZZcE
ZI8TYPs2w7V1kWfQIcMZQMGSPoj3H5/viMxXe1dQjME1nyvyJDe+LxvCXZgouAXJRtmGGWvzf35L
R3SRc7p5ysS5jx5tsAsrfEzCpsYg4AU6Lw2rTV/6UJXD65VuMPjT4jf+cLasCJWVNsOloS47etAV
3Y0KZRqcuHAr9twxwMrQx9nu70lEnDeZKVTKjpTotHUFabsohIFvhaWiDi7NfA4ifr64MEsoGpzd
DwPHebcFwTQk2k2YAApszR39skbpr1UxyN4r1Up0ODpWLjxrKLQfTA58Dpa8BadlVH6GgrdAaXfj
+gbdE8IiMoSfG/8lhIBTCg0OBz3a/WgbjMW77/0ZeU8yqqco++D8owxjg6P93rgnw3IcgluplZZl
4dFKE8hpyhpfxlpVZBxaay6liv1Avl6WZEr/1XCLlo5C+AxCdqhisloXZYPY4a7f2NfKjjRPH3mv
PXBzWsxA1wdfTLdznZ5oNBU+E/NmJTmUE7KkSKHujFcHL0Frh0FYJz9dZk9bZKMKPg4KOHhGI6XZ
h6R30htrq23nAuPLbiMgqdB5F0xmS7zqvFCDJe+ROI88sfa7ybpgaUsBvm/c9Uf+TxKn25bT1R32
gaPGyIraEaf1LFtv96YuUqYDcfO3DdsLECGOW1u+AP8Z+xwbDcWuiNrtR7TucKxtOi67cI9JWiCr
+5pMlBv+uOLdMxdXbZ8vMNXCf8nk5gL+z2ItOoBakkUbsYASq0yOSzcXto78vaQnAnjehVSvJYeK
KOlNh+ZMskVUXd4vpz/RN0vGvDoi7fWSJeijlZ3hDMNUFujTm80Rw8JU6Ifr9SQ4VneW8LKgBEnw
QA6MdLsh9ftdgHQ1QkJ/1BZh8kDv16if/p1jMDiwgyD7TBmgJ+LZ2ey0neMTRlun1/BeT9o93nXk
zTB/J/W5I9ZPQsS1MqlLGZo5t4xSHH4JDXFjglDESDHh9DwDLYTdlAd5SPax5lQC4pCjOrKijA0V
GR1d+uyMN4cjbFsV1EOrL79xISsYEvyfij1AI5Yai1LNO1KlBjuO5ru6SbWotcVNgdDA+fVeWc8p
Lxx24Pt7gMS9CMv5hM03jlcuWn3mGu4kDyyLEYVp7jlcCrKlM5oA1H6E43RuJpstgRD35jHz7EVS
f03URruPMYvDGR24AYxgV5l3RWXZxS1AYQmWUpVUqTmV/6dvOP2cR2oPjwNP1Vb2NBOrYCUrIQ3B
zyz4rlKbvWGaCpT8Lp3Fb7ZrjPibrVUfabmJFnaQgZJVeU0rsfDN+Cyr+kPyzY6m1OuTRvLh8y+H
nRG4SkezP2YMHeb0UvVOI80IYjNzldTvPR4cAw0gFEIxP7UWWOifwRWkxC5oWinzQksB1BxHH8BC
jsRaXiARMW7kn/XSYykJL2BqKB0YyEkeWMvh3u2zPlTe0gQ8OKHOqnIMqBz5WvVtSBiInj3BNzMB
ZSh4XVGybr3+gbE1B7d8Sk/d9Nh4qvVnAXOJcDFW22R7UEEnZY+oVDU+mcdZPyFsh56komkuy87u
5OK0AtkHC9eLbv7VjH1cwvc0m6EM1c80jnHKVHeSyt7GzKXHY5geXj6E0Mei+vrD/oQb9iuUkNQe
vaMXtubOiNpeJHHp6YnFDCw8BTdD5VOEupaEISCpix1qWkCm4USifSHcqJra79kVTWA/j77GOxGl
unnG3GwNT/AySJgf/H5IuZDdtIsFUGw7rI6+dYRlbr8sEYvLSN1YTc6ttTu28valoEP9PF7QFEEg
abdKNxY/BG76sJ0VquRt1r5k3hmc7MJ8LEEDSejQYuwaOh5OQ9t1qP3P+ijmSTm36++JsrIra5cX
6FVByo1FXy/dCDH2Orqkrb/A8aLDOuzeR2iaQt3LCeRCDrbb4sKY8TbI1OF3kd7ePntXTwgE51o6
2GLwJdYzuSdPKcmiJiJ+cOtxplXrcs8KbchRnCFC3wKH0gsMoSm4v4mZ4y4f+iiXSa7r+mvlSRfJ
UtPRS1PL/YRO3AHQYq0mh3uxRLB8CgeO1LENe1/6DElrN+QDAR6ddHMy9kquoZGfY3LczYrl2ebE
5GfxdGJ9Ye5nvvWJv+E2URPUqd4lGcq/MXBjeIacBIrcbGoJ+EmODGExcHh8IaLZhyzJshswyfR/
z77XkmwnuJ4IMOr6qI2ke2ZA3ZVhaeeJh7c1UUTCDxLrlCK5OzHl6u5we81WK/yhfKvKpgXp8c0R
GIpJNn/wIbMiPKkg6sJZM5DxpByzXj9vrnJQbqvH9odH2h44WEmTFoyCYtK/jhPNSeRtRmaxq+Nk
cNnRVqNCT9/S56vbts6RMtlmVy26obd3/RPIA4VKLXu+LTsMrmtQ2JoT8mJIw9SyuaeLL9de9zYL
/Nn5SppXeODsNgFD45s77FDqo4aJ4HfNSm+nbIx+GuVtIiaLS+OCpJ32u2P16vrK32ScaV+Zw9gh
EwSToqMKJ4UZ47Bdg+EmIZ0aK4nEV7/u+XymQ3Ml3dwStlWCkkwVQjFRKrm0MlhQADiu4iOdZgFw
Q+TGSXDC9dcsOZCvnEks2wnP2oclIBbhQD6wEgm8HhstI6QVo1PPmkreV8eyArr5DYtcfa+UDpoU
W0Nf781asLjYTcC7LFxFZrKs+3vUKNcn/VyDdW55CEVtTDNpuRJAW8YxgK1/mGpLblv7CRVCrmjO
IDrji/c43+W2vFdOFjbLAPgYhSb/2FRZV3PUCzEH91jOpswO8NK5n8uIRKq791HHuJW/XQcfadh0
GFwnFg2SJKG21GP5V2+k9wJTSphabhTSb1M7e+n1z22+YtKZL1Amd+dflC905xbFVySZjeaK9Pzx
uIMp9Hx/AOztP4r52nLpEvIe7Ytk6A6U0G0B+rZtgu3B/nxXIlSqk2dmnjEaegd6fDjv/MP54f+v
Bg/hxNX2ZfBU3Roro9sfLFYAKnJU98IxEpJJeHgTivDmtdGatFGIqRDBpiPei3611KIzEZwHQCTb
WIbrCMSXQvEcdB9x2oUVETdXmOrYRCpy9URwDL882VsiLF7K1jJRW7GTJjY7CUTaylXoRINDSSEU
zedYN+dmN8bUjayEdFy40XOstmDAy5sP/IThrf086N3gRFp141CbpA19jpuyMKmB5H0bY+eXkKbr
32PvUkJpwk/qf/xlf59aJsFhvUd+5WCSzLXVS7lqZB79b9ogbwCg5HSUOYRlVfbCtwCk41Sc1uW2
zjyPfI9B7IlwfYP+iRz6gc5Ei+HyqLSRMztONDvaaLm7hypV9tYRAudKJKSmixuey0aJlr85LkKn
szQ7ReMePbJbDsJB9koURSsRkHiqcKHwmUCAUho67dJwcUJFS921HbeG1cSPotY/Zh7EKcj9+1Op
2Fv2RgxssJV8hNgmKusyE5MSDwMC76TY+5U0z7Wf/pcZDw0SPzrxTxSThXyvmynbM0whcUIPb3uX
6luxzZX62p7cMgw9EOX1t/OAt3ewZ3YgzdRHLjebac0eACwEr0NtqewBq+wvS0Ujk4ORePxcUtyB
v0tlPAegF+8XWQtj7tM/8AvejW83HIbOW7GaUGHpB1PehZ0xVHXT6APWQwqNQ1pw15vpIHIKrKTv
DJgyslQpqEJndx48sMC7rPh5IvQR9WRQSS2316jaY8TMRxOdoP9rLbnbCP2RdOMS5UskOu5/lrT8
EkNBd0w81Ci0kUHAhIZqgcj1KC/hmpy6ooIRgd37wqTFJBFlALKo/vmfmreek8dQSjdm8V7A3+6+
Ye0+RPBNWaUq8qAIVOOu4o8KQKhyrbucLI/bS40M8aX4Q2j0Izt1i/jQ8e3ctA71egilNBk5tFid
ixwlqkukYCtLn6Rr+mjg3t1ir2ZmoKZEK0zLWZr5wSubR/A6bJqMEmHRGA6xiiYw0vfwXWn30QUf
5rGqIS724PMroN4HO4EACleh8lJOE5K2oz3ISvT5RNVcbyJii95f4WHmnhuypjRh+Fl5KmgOcMoH
74KS/lt3qkKmjv9kTvGLq2eA87Cm02iEm/MIhkfetmKOCoVa6y4+64S9cDNMpfiH1t0Eyol7pqh9
7d7XVEcuoiV7BKkS/GDSQ3PIiQxWRS8it9dHbWkHBq7StZWjp3ELIDO5/k4Z2pZrD5cj6Z7Cq0sq
sruaz1nUNDzPGIoFWmlJQluAKFO6G24uIS0g7BYXMN+O1ITIwVvGL+8Dsv/bEN3LOYE12xEPrrMQ
w/DVzDhF/BI3zr1rKFzjq/cuOoXtK1ZeDq0Tx9UTxcgXFggXXzjGBe81pqixXYeqL012MvOuyDcG
xTU3p5vE/ZQYWlXzChiES88Z6dc238pgzN8MG8VyjuG6cmIEh9tKttxuTpDN1MzyPGF8MzWT3sH6
g95vxVLbGDo8js8MLkKLiZP1xk4feUXK5/AqMk+1p+3ZDEEVM4Av3UAvdnuP0Q1msPH9EiGEjTtY
3LAkZ0fGonycFqaYIqgc3Gic3Re8yUkkXiADQvXh9wX7L9j8YgIDGdyQGM671/BuQCZD/NBDXp4Z
XV56/yyK5Ji6mpfx5bCA3PrZWDx4gmKU5OElUWsg++RNWkC1fZnzZ3FsBMKO/SkG8uxl3C/prJI2
pux10gGvHX0bgxlA+AfEfYjuqLvDgMeALWr6XcY1+UZtI/KfPmPGlyZ5QWD6ENOI582ITSOqnatg
FCdEZPxCTuigrwMdzNGNONTDEMNc63AiJAKM5dGiCfnyCmJxDtAtE7hnLnJHbzLiRf57kYMEVNEx
rS588zqHBu4vCECa5cVAnrYhS7pafzVXJA6XjQsyw/HzaQ6YuCOFF0TZW6SKtqd7izsmcZUfTq9q
sEiViUz1vpXYKTDGfeu80K03FKNbrWIXPsXR4PEc4FetWKGOxqxe69bJ6N2nHc+EIEFiqOfFpXYh
S6cZ8WcCZEG1YuRazDYnE5fi5qsL43z2aMSSf5vrxCAcamsR7JbBaqNgUuswBbXFMcUyV6VQS+u0
aP4zB1xxQNcNgEvf1zn0gIMiDyD2MWE3aPT4fYR2foZmV6a8vBgS/3y7h9ID4twH/Vkey0pVJf5F
IqsWndT+Bg7dZGpJkCV6kWdvlLXm6NqsK/OvPSbjLUa0HSP75+EUJi/sOywwYjvKadfKLvjKgD+x
RFetw+DpRYEs0+K5FsVARLJxN9R45R/P0fincjSwIihoThYq8kU/jktHK2ZDJxO5K4UdISk2R1AD
Rz6O/aqATd8qtSzQN+DI0a7WXNtrdlqcVK/fOy8b1dXeh649l/Up++FDxZBXTOQIC9BXIv4jWc+f
Wg+1xZ9uSlBNh50PYb+3TfHHmxeW+uY6v53KOhjMl9ynuGL+OJi4rPSE3wNbYh9PzQhgBedzleeb
AF+2nRQyTLx9REHfvZKIJxKUFmL92cZVnzQhDdnw8BjZLzcuw9uqW/R3FClxSS8T+A29FLWcaRtB
l/X+foGNs6uj48J/ERxT2C9cjnuAJbKaMqnglWbOOd5Yd7WcsRt4lRefKXSGcUUBDFR4sUJD69ar
lnoIi58/rehiXvr9WHrJuadtwMREwxT+WwKWpWLOS6lmuvCnmchz4Y4QC7vFNerbYYHSQvxEVHBq
qr1jy6l2mS93J8pZvVIPiiuTdZppg24upr2uCuZ4eW3IcLzslmq286Kut6u4TJRYJ7Vq8XOZCKH+
BzOJMAdCyOQXafs+FMp5yfU7g9x7TPSQMxC3ZHmTNvHx3p+EtvcEHgbkq5wn+9pbr1uteFip9qmg
hE/cZVp5SohQVmrWFNKCDK7wcX9oRewgu7Nt/b2dTsy/7h+hikrnIr5qi58uV+C8ifteXHSQWRIh
PUZtUwTLXVdU/iaJ0wFJnVU5gwEtLd4B9wMPYhQPHygfaQ3RA6Y2bF60Y8JxeyAoq1YuBrlqP7RN
PrIlH0WGadqp4KzuG2xJ5tGMbHYjVpJXnUtElsNfle3FGPeOjVSxXgWfG0JbNGd9Pf7+FA9HbVtm
2BYBUUxmMq7CaQ7IicWWkuTbKxQQgDRugoBzTW4NdCmGgUi5TESJaLXKEjA0QoLGfqgT4PuZlNBV
bUsAFapObRrnag00VNfnxVR7ZVCg2+ITpieD2bMzrRyle2ZdemyauVlKikX/Gd0nzJy8VUf8pk/y
9h+coTp3aj4iy95OLKY40GhQElGRVPL0960lCSoFkgxTRdjvRlt75oKll50wA1NaSNryNkEgnKHY
1Rvla8vJry4t1S3IEDpT3HpgMP7leVkWk+AFTJmaZoxUZNZLlQ1emjCY3oTzx2jjGQEL4yvEvxfu
jfnQc/GPebr2Z6i57gbUpbzYHmx9W2tDAd/srqOh+yoEsd4uLq8BUrxpI6qs4Y6BgP/YXgUN+YSs
iI+Mfu8anocZ1AyUAbsAfVdGC7uF2KsYWvYbaiSr5VDpjfRTWZ5ylHyqmHY2olKEtCPlm8d/9C6p
fZcp26zxIS44rmaFCgYof2l26ynsnjoCjsv6rc9TyVj5wnjSrN96/XnVP+ruUwy1DY2kXp3sbEN0
Npa8wC8pM/00o9GE5l2HtKG1YVpVfNeDnopMD7YDJZN6ntYxBT6rZTrPBVms1+sOxeD8SIMEr14m
Yl9N4z36obU2x9pPVCg4JM296nrb2bICinKcAV0tHWX0QwBd4Juj2yiwLrHr2J1zCju5SDQda6x6
pIWu99L4R0F4FEoLc/JbH+bY8jZdY05V6UN4n9ui/pzId4k/I28Pb1oHhICiyo0I2idY82FZ6Tb1
vRCaHWl039ZrFxDJHewzaNTT3Rdbn/D6GTxBK504o7WOx7/Ydfkt+64mygjjoddmhh8SAiPL0fiz
jdTf54vr3OaPGvg1JaU7AY5WOHYaB0LKrEl1jsz4JJ+FH/N2NVBoCNsJYoy2pO5WA1r1SkGE5d8J
cP5c+W9Q89nrjrzQ6ib61KBZ4+s+S6k+PP/fZ5tyy+L9zYLVSbf0EC4sbuTtNVkmyq6gVAzV3ju+
uudf4vQGWYgw8W72iB+FC9Xr8I5vZyL0HG5QBmujQCpZUz996sIgEuJxtRBtZ66NMKpxXvIeGZNL
7IaQkW4wN9G1geKzWLbwr8dCiAg/fHCrhCkMXVrO4E6RvDUC1MlQqKI73ivTFfKZ77nmQ+Znfj02
8xChvUmx3DVraQGKjCUU1t9SR3HGUULMTwjII0C4rNv7yTh1l61U13ki34bF9sJUmD2n8eMs4BM6
XFlJIWg18DSiiQ9zMiS9z2I0Lyp6SNLb1IoGIiszOsPpeT9mA+YcKvx72vPsl1VXk+WeNEfAiv9Z
IPKHc16Z0pEg6OLNhPqLUO/If0dVKKhv5Gos7vpakT2FDkEvrMOb4spBIjugILpuFPrAegZUOA7H
4veazWuqDKJYcFc8C2Di3wRVW5VF4iPEZFM3kUvFibBA8ZVjIr6pNfjQRk2K1wRxOoyiIjWj+e6h
uQXK79zut1o6yUn086TeECKFjlUSPVnKnSb2SKCzRMCaa0yJDEqZ+BlUsjxdGK/eu8iSlQWfn9hW
UlZZUb4gr/dfZj35+8XZIDYC6CCfuG8s1G0eCxOUYqA6OExwxnGsxduxR6tqDrsmr2uQdZr29doI
ZTvAmNwngEiU9jsXoGd8+tE7RmFyxHPEMntxqJ4KwrvlB9e3MJYSF8IEGhR0eeZrMR43gcf4aFpg
/GuqVsK+eZSWiXJlVB4jSioZWwH1Qycl8Z1LGAHZmXkoiD4TBigJYd1CcEXW5yUmurq73okLeO2T
2RwzxB0Oex2Zsn67Vf2nIA/YKwKYZydbG8hEOdgQS20ADjdDOeSnzZuqyC16sy82+YwrX7E7WBpx
g5fGO0lN2JYi1wnTvra6UHSIuxKJSrhyuy+UGbKL4rFk9Y3DcCzM8CHdQDOZO2RD0MS1hdWQWRRH
5+EFdiL0qS/o5zhOpoojHl7ijRVdhNPtaoc5PsrWTZvZACQ5t4WT/8AVoEtty+9AQiCURvoUdSV6
u6nqbn1qcAMbpKK/bzpMLGYUMn4+lqwQyjdzoWeOsiorbw87tW/pJg19b928wJd8vpvtgy3kFEfk
s9/XyTY/M1D55XK9NtaFTCUP8HR4Ba4Xkgka6IweoaDkT5xVfvE4b0t7hKbvebyjE06eHiOAqDqd
4G+KoUGqAsZs8+rKHK1olqFu7HbLzH2NOmYQtUnNO/LPWyNGlyq/eHKr1KqZJ8FZ+WdsZ+xJFI9J
ZJQ2Fo3chda5IN9kbMJBdEzoOwVcwYRM7VKdmS1VZkMwAEF5wtJgncymBREHhRJtMhhlDiEtsTH0
gVSVmyIGxlBIp4VBou8LtxdKF9ikAIccwqAVGRp2LgRnSOJThY5zAz1456uv40tT5i+KcmbnYgpq
XcctQjPJ9ki3gsDXXjld5slhuhrC+sShxE4t4k5Oijjc8ktGPMlatrFLHCSjoECbo++qK2h3uuP+
zF/sCPv0d30Pv8iJRhLXw0sDe9U0rsPUaQPoZgtyKgyuwQfvgmb4Ou6iKdCZ7CFBfHJtBjBRHYCo
X3YwaHnV1eceSjfK2WxhVfVYK75jkqOTjz7GcbKMbHNtG05Q/zpyB6k4sh+vJy9xcvWAcwJQK0uQ
6uFQV9mr8u9sDa3jcNSG4OOdQIoW5E/v/8JCRC5YGvx1/PzcXZoMIdwHpEv2ahfjSBG5OElYp0lM
Yys0DHQByfO9QJvJVQyXdBZuiyUWjvSXfvJarwQOx0CVaCEZTFFuGfDkUxH2/mQeo+SQFE+NOSnq
qowIMUKzqcO3GF4fl7QbsH9ARYdsLQAloj+dnb/LnU/WT5Jewz8lsiINP/EQr++KTB9TNlL+S1dm
Xl/lZ6ZXUp8lZcXFAIKooCYFLYOsm2+FIIBgmfnscDfpdnzCzpn3t5zobcmN+7LBacxCkyDEpjOS
I/C382SPCEq4uwuei1KKN8COsUnNFbWlpiJlLcdkWUDpAJ6UW1YwT1r+UM5sBeU7UaaeIMhR2HgR
RmQxVWpNyk5Sp3pejEPDB3NWel9cR1zgzDO/h/OtFoLScYHRLBvRx9DifcqOXSATcFzLOKlAd/Q/
eiQc9UT0dyoeh3vXY49ECkPi+XVkb22CBnjKutofxcIAcb0AGEr/WhocvBdRt10NbpeyWohA2uMV
K+ttzAIYQA18buuaQzaBS3znT5l27LVW3f3vqr6/sLA75DJQDghqU4GF07J1uxYrxnUe9U5U9m5v
4kZaWuAhT6gkzuljAadUSEpYyOv3LWOut6HcXX6qwHhuA/GgAppxhTYj1A20GePgCMRcKXHOOAXB
rDz5T9emH9JYtyV7nXB2oWOjA2oN2RcE7laYezEjjIpwfGGZKQ2MI8XZrnl/Bnb81hayX1aBriIj
2dzU4HIU1EQn8FKj3ikGYpqBdsAEAPfr0YFedNw24BqnK8DmtMuZQ9mIJsGEtr9HDXB1FjknPyL9
mOQUXQplbutPXMPsWo+FjE/nKClcdTrE/VUGR7MBO6wE7efFlQMLOCEX8WgD5Q52mEYe/2mMoFw6
ZUVZ6AnO0JyH2areayZCg/6Cn29A8Djto3n2eRuV2dKGhiMEkNQxU6htSfJvKFGD/XNN0ObUltZb
ldIg4Gvu3DtKx8GKq9G9Ark9jNQMd0eWyowqHdGtKW5gNv1H7syIZLlH8XvRKaCuvUk+8jqfLULt
yep1mlfoc1+DDCi0MM212jRmV/hyc/lQ0b9I6eF9CP2JlRbILVTFCwu8P1G6OygoWtI5nZBihy6d
aq7DsjCjouUEFSWZpK9NQuUW+xAycPh2yjiheubtZzhb+U5sPvaE0k8s1UlmOqiNMCPZe/QVoXS7
v4Hzh+PTTRPqH4GExjJ5qh5+oKO4YBrfYV8v4FGAzWJaXOk/Q50Qt6mYzVdQ09Ul/hVJihmqOs+b
BDNeFxnVamxfB67d81Lvk5i+99M92d5venNaiWxho5jW1YfZpDk8oO49VnA/Fbh8sY18VVx3RJhv
XrtM/u1azpwrb6Piy2AwyIFkVsH3uJG2R6KeRE0ICa4EHF8jGraMBA4FotqeVdNVRSSGg3evV04x
cJrVU5LgPYIf/xRL8A0gvljwiYSRNz3EkkisKv8c3tYJYztDoylZckUltYxy5q/MDpmsKOrk4EMW
GneIox1OYxi/PfGZ7C+tH15YFzdF12l9EFJR8LN1ESNL4aDGfzQvtG6USy2CNY+2nRktt9aTzbeZ
vTCVis4qHKrElA0XSzG1EsOoSulmFRcEWj1Ep0ZtU56YD+YgF/3kza8w27ffFWy7XJ8G0yC6NQLE
94Py5nfG+CBEInVygrmjhf86U9f+B+cMng/cHyZiboZ8lwCUojQdtp8GURQUf0hzXJUu+hFsPVTb
q2Qz3ayh7fZKXDHvOEi1cSIv30sf6igwrYM2C1ktnnoEVOyfPbABKIxFn5yAB6q7YnhV0lteoV/3
JdY6wiNiR3AiflMS6XgPRk/CxF6jZQgLUpcn6plK8z3ZKHFGz1ed0k007p+v5+Tdl+BeoCuO1VaC
ifb7RSW4zynsnDioRNENf9nWrzATy1bTJdEyg3S4/bCTSkoeKs9TgnlyqektcrDVrkqofUhl4Xg2
Ot31ZsMIkCUGT/KiCS4Bi4+jO+oiLB04RdSrYQqrxs1+NI3c5mjW43XjAg0Js5VXMWORbfSTluqz
Kf9Enf0hBagSXiLZLT3QFI26kk2vXH3kIo7vsm2Bj9iZj6McV/HulH0GN8nhmY/42lcv33lxLJ8W
8dM7f53dc1wKReI9dy9Fkx5xr5z2zOeb6UpLVNrRCibofOrqFlTq+XfCIMisHbnKVoInyiwc2cgi
aXioN7uHHQqMnmqrq4+AT9GDJZ95Ka2GfrkgO/PZYScAdm+T6UU7XAQK6NNcIKNbn2+bvQ6f85ke
FUNinjHv+blE04AVRCv3xO8uD4XSqw5QQj1wtSohHIa2dF3wOr+kJXdoQZv2iKsWgWRGVPDUZvUG
zZSJ/Gq/3twiDOp/nFqASTmXIIXoeKoQMirVQ9XINM7uIpqHV+8HWAISYWwIoJah7ADNULu+IWWN
zrjBAPX/ig/S6hAQRIErUlXR1/soqiGp7EkpjCFzmEVUFVpnkp/jmA6IPAqf08kJoLdjW/CpFNpO
86iB67cjXPdkgr+CvWlwoxc+rS//+sRldZ+4h91LfgjT5i0/ptDnzSlpiK7XzpRNso/gUfVzrCJj
mKBY8hELKs0iW71Me+BT3fMzprYah5w++y4Q+aXmjsFIi9ZMu3xPkXjg1zTRFpbfHadFNVrK22Er
CDNK855ZGjA7z4PUiu2rnPLtb8HCmvc8UoSUW9Bnq1iMQEUzmOYJb5TOwUx1apr3y7RBrWz/U9ot
dPLb7+7tk1CVZiYNFkT5P5/PxWUSJ3fRtEosakGo8nFC1WqpE95ff/YY2udxk8IoI6IWzjSGB/zj
IafpDdKrY5EMbrH8EEd1oaBUnjdtvWti/jlLGkTMD/KMk9vF3xTWdOcFUtqlbx3g5dIhfQUeem9j
MdDgBBaNKzkygBohzuv0IwDKVmhNsVIdoZgkGQcOe1kHv/xJiSaujyiQDjyTxtsPNsAOmMgUl1PM
Cd8ITK3Qsl7tBqit9k0G21Uqz68FsA4hYz+m84KX6g4vTIIPkdQCsrzphvUifOkHG7sIP+WlmoAi
Es9Fbb9lWHfr97XYBjd2+VsoTMI0sps56n528zsJ80wW0urhn/BnBDsFthksvAvaoNOdxvaiclXL
efGA7+Jneu7AmRdn9ne6+R40ZPMbH1s8aCSR7lemga7GRQj21On0Exb4yEkdaLJwCL3EvIgONjcD
d+0uzOVu7B0P7nTycthzQ6mJXNEqIfrV7AVOQ9lL/RdpY7BpDsLhlNG/OUtwPo7VVpJ2pNXbKL4s
rKk00e2g4dX4IMRI4WBOeAQMWCgFp9cMIkbHh2LNdKbmJPM8U4Nd+zcOct16ecdiiN4paJkyKgfa
rKpR6LCAAwexBSzvnNfjIVnDq7Egh0E40fdTpa2c8OCBfGoy4UTRojXxQpBvb2xzi2duiWmnkY9L
MkhUo52CjEdBpjzfwmMBc7jVErcAdXTSsnHYmaPKTTrBy91i1Brz/DsCaPhsENktlcqrk8zGN3Y5
w1NRviOeJxc0DEaesSHkCJyevHf4a4Z/3cWOn576w9Fu2AcoQpnV6+xcBT+MoeBRS4UciQjNX0g9
MeZyDevLARuJejKqfgeQjSCxE2R+2airI44R7lJtYJ8n70LJF09zI7F9N15GLwv/04/U0xHkcgUo
J9PVz9HpL1QEsT9UyBqG512uF0zK/MisojWf6kfcrCslX/RWfL5Y/bGC2JAoIGPRCd9TReQ9yN7O
JMDzRUT2x/8zAZiSb+7k5mOkWTO6D6SbX59n2F4SPLFK39QLpwmtnoHBoq4GX0o8dTcHMzyvYSSW
fden66gJ1DBYJarouqD7G6F8A9P4QIUbmKHJ7SnGIwmw8YeodFLsRT+o2OL0zXGb07bKdIkvrPWr
IZnMDwT7xAvShkH3FtrHgNLhgip03zgJkLvmoPVXdHxz6ciVWdPEBOeSo2wKOQm2jDrPVP0O0pzY
mxJxM+9nXtbymFNb4Gq0R+RPTtB4sPVTXk1QHMBwtS/XsZ9I4+fBOjlaC2ZUVn0C5sRt3GQZFGSp
Hka8DLtnbgwWZk8jBSvqKXxvJbU/Vb8cUhYuUX3jxOboctHEVRz+h/FhDwrv2oA645y46Wd5CiAn
gKSCMIiI2X1u3IxU1JENxDSb9gJAJyIcCUI4KUvmj2E3so4srQR4JAonFhigQk3fRpllhIYC8ywy
rhd/KQfhHbN5MhvdzTHnnymTx7j/3oempVwcx7bq8uYc5rXaTXdgWwideMh+95c3KeZhPgwSiV+R
cbr6LOUKCMYZLbIsVddJMURhO5IjdJ53LsuXGH5dyFoYlKwO/Z2q2kba0M02LhtFbbtbWumURN7e
cDCf6HGjMUIAS3ms2BUjgOE2LmRwV9eOnL6OQIle6kyEAqmDMo2aq8BZfs7c5Bh3pG9/stE9D2BV
NGCT1vdthZReE/MU5aX0EdqtLFmiqhNafJCBZLS28j2oAlWHTJlN5tPPy1+nbL/renxySaACrqzD
B6DrjbT5Xg5smxMKA0zKu9wVk2ZRIqFVeSxFuc8udR6vkS93J4Xv6La0LrvGjEAeHiq/Dg3HmMYD
6DUEgmMw1eCSeO0Ne416qIGnVxZGb9YZ0uIFUzUCyf3ZoIbiklNFJrpMaIQ/FOvnzZCRcd5BKaG2
bccralGTWPUFTbPPWxQnQzKKsnjCU/G6dlpLdthxyF50rTVPFoCjFoA7PCW8ac7650QYVjDIcgk4
21DF/Jml70gg0oMjlVok/L1QwLnkrJAni5zafZu15huAqnE0I2ZUFOR/e7M7/CA2QfXzAtWj8bKu
1aTnx8pLq7mP4MZkfi7pADWE0aRUioI2Mup4zTkvORZop/7CZN3rsujYLhQX+IlDAP1LTRmoLNrC
ZiU6bXQcX+FnCmWa31flxhikAERqMHYnKvQbCOZLK60ZS8hJxJL0+gmGSVZSo8azAD43jxomuvS0
sMD6u416GYefCstO/jYXdYrpas4MIWegnMWMmfHRXE/5F2TPd6uWaKOxDWHxZiwkgI41foL+VZDz
wxQxfUfwFwbq1/u5HtUaPbif4RLI/6nCWCKHAW32awn9NtJ4VlNxUcPRONQBuDFV214pmckOvbnm
MpN5Zmb1ItjqIfkfJENRcQfA9gwOm4sPDC10PCHws+aiNbovDzVlBt5hYm5rZO/5JGlkHFCcAa3s
edtnZzbj+Qo63I/CvRDlxWgYDTkZbZ+oOCXupicliIegJ46H9bEIrX+8GH1HJ7ABlrEuSZ3WOnuw
D6/TkBGkFQnAAxN6fZQC+KudJ8VWcvTp7abejA3uKTQeuS6zxQI5BBTvjiE7ZaKchyF8wHiJOy3R
20ahRlY+8BfUgDxXdmfXQCqNhe00XAFr1YtcET0FZr9GOO4NVjpEzk5CgKTlUYmbh/G0fPMUlSyF
yXoEsPnElvpfJohs/deYZstd5Zu0T6L+OPCoScksYUs+jVKlTTx4JMN7BHpnKU64wqo6bENdoe8Z
SRF+wSJe8U+di7PLeAv7u9n1Q2rlA4oXKRD+L/Oreg5yaoM5kHY8oG9ByWXP2v9LCzAFIfe9Rt14
ntAmf+RVyv840DojpaNRQpqNa1BDKL7RLf2nylvPwcw/EgFV8A+ztuP6QwEYJIDBuGo+tuxdPO4H
ibbvDCcEA26IsFjEMktZeNWJZF6nhTAvgriJ+XMuWIxQDlYJcxipf5Ne+/Hce25tuzo2WnwS/L+i
MeVMrleuY3l3tjOM4Evdp7qG7pF/6XH47hSPEMoadr+j6JX1hNQqCEyyqt+gfbzxqQCetcck/56p
BmNPqL5dRejPr0Ve8/IC03PkRbrVWYEAeHK/SZQwGmDY7WvF8rrOPsqtWzAbPYcpYs6ftXubrw8/
zc3ITOCf25+M0qH2G67zOV9iMIR6i/ceXGbKZ/B+Q6Mv4FvXLuLC9SRXM34lcZMjBeguu1VL9hDI
DnaqQqLqPoy34uAsoPtD6ZjHzvnhJoRuWwBSCZaumoP3dLhORt0uzErfnvFfeYOyvpAr4OdqF/BN
dNawfUwRRHBDQeguyvoak9TK69qyjcuLfI10j5KB2s/HZVjhpgMFgZ3NGJd8ly8hM2gvVZQEW/lQ
tG7vKEcmEv5lzjyhyJ8RfTZAH67sX7CfovfgoQMH5+VCZfSy0L+uuxNa+cuveL9539XWLP72FN2Z
hFhrk4EbYgyyxnDISFMdFpdz8gmWsUnUBAiG/brW8GoEMmzCKg+5i9CUUtCEzLvJVal4nTg1yF/n
NMxJyijZB1AsYiZWwXoaECkFZ1IN+920+gtCixx7OzpDEqNKUuLgsBHolNlZdCbmh73RR+/Uq+DE
WIbIcXNVXhis2dTUXAZojzlCfE15yGaCnUlANwQT51SvOpMn1b9ERShx3+rsgH2wy37hAsYJIkUq
4r1ThLYlVwIlZUFDlGyL1fKUkFLADBEH/LpvrtUPagijJ3k8xuB8qJYD4znVh6biNVQVx+whhcev
IEe0mWfCjd9Qd6kFx8H8Qk88BKuUN0/xxK4xYQuuAxRan19l5ftgVO2qp+IlVI2raradHTRew+yj
Z2W181m9GRBWW7TzNY0WG+wUmhzVDj/blapGX+7/pHpF0CCSYJtZPxqXjMgM7DrD5wVdVqVtWMEr
X3Bu7sMy4pXqtQKZYiVMRZhXEDomqf+LOFxEhm6u/0SXiMeuiA2YqUvTSaEuSRQDYcq8z+ZdfI/9
Oe4cmi208/LZYT/BA9eVILyX7E/Z470CGXtcVuxz6IgecO1u7uVHxr0u5W9k/rFuqWOgg0Nku6tO
ja9Pd49tqPfU9153/G0vDAYuU1+j438tzd8BeBBQ42WLfHjTJm0SPPh2O/VEXsDiuChDDTSWMEeA
OouzKcfFSNDsnqIgrbICag8EoAMvTrCUKpO7Al9eIM61kDOuUMlOOb+rGOtH8dDlosH7zzpwOHo9
u7nuWKprKtrvQlF/Wi9IRv42r7GaJpa+BfeO/gEHb+CRsTaRUk2aLRSJ/6ckbhWUdwFSvjkS5PVt
XICwcDRQzoHDNCCKKtTocIFkewTMTWfzbqvHy4sICRJb4kcTLv+A6hv2P65Pa7BvaSPWLq2stLKp
xSTVHJ9ATLWBGdq5II9hBOOdAYQQX1EQEW50yzKbTtgJWSTEHXwwoocR5bqVRqIpKtOZ14vCFshV
TjdW9lMMUku8JS4v2xGhj0FdyqFy/CZW3+ptBgw14L7ss8uQ6xN0TZwovZ2KzUuNEtf/RiCrkr3J
b6WjeXpNPOpiazro+CFJvFwxLxF8ZNP99hcw93yQ5fgRksGOWoq8H6sv3fzBYXFO4Ogt29CuNA2R
dM+37pwEm/kP996GJeDEo5MWfSgaSegb5ss50w6hZfW6G0Sy6LkUELJUXGa+alFkvsZwsuty3rW/
EfYTxQo+KIJ7ohTDiHAuzSx9gU5UylGlxf5oVK4eYkkDnVhRchxOiAwavna4+qM8FvARow/6aBSH
GevX2KjyZjRcewZlUmbQDj7yR4BmiJ3ajNTe+ahkMl+o9kJK6B2asL7zXE2ldPPDroJbEaWMGoCN
zhcizd0IzKpJmjvqtkKtPxnHH3sqQ/rFHUJUTbGQew2qc5FyPsM7JEL8xdGEA+tY/aJJ7v8GP99l
mv3gvUbFxqGPtwtPvUhv9dplF7MrqMMulIYmh+FzXcoTVMdoRHZ5DOFmEtRn928D1BCZ3U3ThL2A
rOgTadCM6Dz8Gz/k/IQbfuaImMuugu8/SdwwEYKzwk3Ncnh74DO8QpK/1VK7cIQbMbBlBdozU9XR
HyM6Lr1UgqRxG5xjun8TgqNwsh/f24NHsnJNTNKp3ORR8GzXpkmNoJp3OrjGpwkn0Z4LNKzwz42k
SLMamB1MUZHkkVdw+1IqcBUntrDiYYwGnChetw6DFiCrt7KP5hQv4/869pqENPcHJ7gMESUHklPB
zKdIbau/Jqj2aH4A0MVefuQoZMMw6elMTo2PMj7Ce8585/lLAwPHAvbPpVmb2CYxcq1qtkDy3VpK
Nl+U6Jd8cCjwu5Utlo9O0wPPMBwPSGiUKfHpHcDJil6YCXIBhYio9qfRA7yAONkyuNZyyMKtOoSf
G+3svLhWAR2fWqnOV/wW5zbe6ciVz5TcfcC1knsHhXqrG4MI8clHFS2/1cA4t3dO7SHC6b0GPqUC
3/PISEjyfQbDYwr3DkTu+MAmkk05CJBBccCqTNbVo490768x6xOylhKE1GbX2OFsSF364Ya6/ecm
lMeFb+/l6hkDmsSX6EzVxFxcEIzY8SG7pRdgR/xbXutMw6qMnr6xlJ8v6p0a/HBF44byn4TmWVV+
EYB2kFoxBh2UqxsgvBm+LMLoAAIDobVvmfTGtUGEsrop/yFIlHFBg5A5Ck6S+Z/2YkmFOxylW8Hu
RvKp0F4U5TxQvyRHfKGOBDgj+fQpjgsq5Ut2k1tLC6+OpAlssrfq9XTjjJrrGZtmtL7gQhXdUBok
8AzYyhAEPed6MTrcM8vAPH917aM2Kvvc7wpeuwYqKkfcMnoe9XA11SMe3loNvUuWrEG/35dkErza
kOJyzt5Z9ujhiYZDJvS4d9Du/EnldC00MJ6HxGlK6mcXS/e/HdfS+QRQKK/WypxgKXoHEWugz9Rv
e+ow1qmS7pFIJuTIpPydbRHv0MkOxPW78EdrG1Ta5JmSX1CLEDmOgkwq0pH8UL0j7HCTuabLzmee
2W/1tZYBcLz8fpfKYAyZ+6wtw1paUAkS9ErTKnC0bTKEW1Ve7v9+kckyVDf4KkOsrD0o7LexniwP
vOQllYGR5nHZr7c9ug2145D99WtA4Sqe+1Io5c34E0wgTR8DO4QTstPRT8bPPU7L10Lg4mv4wU5b
UQzH04m3jPM3XGMl49NSc298375KMTs58aOyqYUtYkq7vHGnnB3CLhi10hOvDVGz0lBCLq18kEbA
qXHyVFXbVtAMap+ipKLRu0WTYfnmGB57Kf0ToMX14AaepmDhKG81CMfoBBEjUvF6ChhWiWbJHJLg
rIXiZNKUWPKH2C78WHlaRdCqYtcMKe1gjmxlImyx7Tpx6wVWlKYJs2W6FTyPYVLqlucY0oxEvVTi
nu55giE1ruMa9C4GHZXeBChaxtBHjLGYTuYWOnqx+WoYcK/2q2wiGVXB0bw4qHdzKBX/rgPo8wld
DThWwEjq7onxxED5uDx86GW4IBN2rUec+DLxWcOPRI4+mVId62oyaMHb9acItDGhdWwS8mFRuOZ9
SVyoj5Kg6f40XE5GCYU532iB4XRtMzKG0MWGvPFeQoYxPCm/Qd+TJA+yz9nVWhAMhLYdZbzo52eU
Vd3ZlmiUFPJ36UJdF2Y9BUhOEXZulO6vOddBL6wsEb2x0Wg/4+8kJKlUtSbuA0tPqDVHvvKfIFfS
2jO99lNhu9RcvN4fzQ1gKGRrPxp59eOV6epoPNdTkc2oUSbfxvdHnCwFzhjeAWcils9V4lopY4oZ
hg5VJw/ZiKQVVrphqL28enNDHeGS+lXyS+yNlfR7lTDKz4KyCuq/aRVs3ag0flOulYfAeElKe/41
viPhr8hzUwXK2iyYK7sO7xHPNEihL8eGzYIXKSEFItdHe5MITc+PoXczJofo8VJr4b6KBsDznRnR
hHi85drUrhRZJLSCnfYjbX1zdbgL5J+zKEK9vpoD+etmDPYJixrF/5uQT6WHl3eYevRXVldZua4T
e+h8GWBUlsU9Y/pNi23pqk5Q3emg6FC8r6HAXofETTbpfE+WwwtCACPtHk+8Gcy3RCEKExnpJG9S
o7KfK2vTNgSyXviYd1f0zmWDrTH/DrPpx7CNJ3pBxLDKBrE+8AzDal99zBI///6BIT2xdidNsYJf
s9oxtyn2oDewv226vPKCVSgw240XvMLkQEuL3yhqQff88knBYv8NNABHzqX6pCJ/7i7rT2pnDJVP
PeTPsPP3fzKB0kbbM/a61gJCEFpUAeKDlQtmH+FuIjBzPAeHa45LcqLuBKUNVDiVR978vksrzQs+
EK+8hCKGsuxj28tx46efZRAJF2z8RFK/rCududn8llS2EpL17zLleOx8+63hKil7bk9Tc9D2WMp+
MAGS59aRelVvMdYz8nnqm9bTxs//TH252IHHAmi0SppkJMua5nbzQdOAjbLbWkTcpzrLJCgyh544
Twvt7+QCHUFcUTB16y1QgDXcaV4OBsGtrgwZ5YFD8qQItd+yN/oojROYHkCSTU3bVCMBSWuDdSa2
pzel5yB6PsqM9ad9y0lu8xRFpLyvLcRnrYnoJ2aPVlqYB0cbD/HL5QYxmbQOv0uU3eM4/fm96q+f
B8J0mUc12DnsNPe62updoS65i51mKJMsLECUALd6CtpjpSZNDkUuiwzi0B1asANtikf5viIyrk/B
0tgiY/umPV3ejWzQAqlnUUqk2ZbVkOgPUyyO9XnH5vfFm/i33Mgx9swhg+Blwrc0fsexh8sbP3Vc
1FiCNYVpL6yKuKwKtvypFuhoUaNHCA7WRpfnts3HQUecRX8cYkXNiEfmQgnawwoxdoU3SqQuysVt
6fHsnWJ9C6W2NR3sAxib6uJdbbSdSK7hjk7vX4h2/kRTNczQAzzhW5LgpZitYVwO9Womo0wGk/xe
0gdal3gfB4rXqwEvpphBs/PMCyBgUs1b7s1AEYv52Bb3WqxEGYduVUOh1ppUDrzpBPSAqyCYoEHF
rY/AC+oUSN1j86hFUof4YR4n+/hcIVrwYlzaIZ9trDcr/e1RAsRD099pDIwlvs8b4hZT9FViAY6x
phc/0w8qqRg7IPjmAgpERDIdWfe0JKK9t4GiZtjd3vET3JhqHSfc1PPiL1mPzWPSpBHDVtv3Db3s
Tl3beLQuJqaEXrcSiXS1PeMxHHEjVW+FdfRYdcvs9wT0IonXck8zRVVFly2FSC8aE1e2LIAE7CHS
QY/dCTMt72X0Q0vXbsqzkdCe3scsJkVqdhpetLoOKTVbLbDorcBNMps3YYITsKDkYDndEYnJLg4d
Hi4LGZwjoW8c8Ax0RB4DCq+onzaqbwAxOeTsjLJ1bUZkCQWbRmALCaSqnDLYu2zxe6ndDjyohVSr
v6YqxHS6cf+CagkmH9+7+HPk44vGgZqsWRFP8FAcyy4fk1hF4US6T/xtYU8JfpOnuEnu0CSAmQU9
Oxa6gaFOtv15SWYViCXlcnbcOrQOXO93B27KF5GQe5C/h0Z9G/Jivs56VkO4Dck45/ynntdl4PzO
hTpEOkC761oj4oAT17WbXDiLsxmjl5FqXzdXE0KtmgymwjV3yQe146gMdsevkWqgGCkvZXawH+eu
HnLEBUUL6k/+dgFqZom1ClHLgHia0KMXoUJgyfaP94Ia5bnIYAa/cJHtDKyXCvIjCxQ/Fy4A/GjI
uYveSiXWB8cJceYz8owhnt/EvRb01f9o2w5gDlXo/G2wLh73EzlEBYxAQgHnoODz3dsN029Gxkbw
JrZ4RaOcCl3vYElT+gii4ID9xHPNAEoDkWWmRqDZNtIJl1xCfXsZKK7SMbwqAISsZP1Z22VIPm9k
loKRC5tqddLVmKR51/e31eO0OG4V83qEfSyDN3V+ROEWReJNEQ74lbpRswbVc5MAsRRxzfKiMJAC
fwZmVGljALKLcpvQz0pHZOMA9gRs0fsy6tEcUygYUqIoEFs59NM8fWw+4Vd7DWw1p0ERP7cIotKe
UvGT8h62PuedKEFMWB8PnJDHJTJ0NzEBsEFu1aqhJZ99R3O5a0pUkrCj+hMt3UiJCwQlYTaD0Wc2
caxOOGqM/LoYBhLNmhPesl9FZZkNS/pwrFJF9SjFmemlcru5Ft9yh4i2Yoc3/VlqKkXA/GfUBXMy
TguleG2PLTFZeGTR6AAmtIAlHL14dzGGG56UFmFQSet7uI4KjT5CaH4M5K+2TKtFIO/iXnSm4gGU
lg4j9pRxEx98I+c8eXAqkfa9jh9ueGIfw4xmaRX+oPvqATTt3L6W93CqRsa6PO21mHB31AMO4QYR
3+nIwd6OWHT13x8UU9KU+WtZ+kT/W/gQ595B/Uuw1pTpSfwaghGKsox5KP1PAXYqtOCX5T12p5U1
4MJmXJdwsOVpBR+S5fIrYbz4C79EehDNbLrrXgV/A0YsJsg95/jSe11ZB1Q4kEcRMW4D8cIXIE2D
kpwN9x0RDC01wx7U6IUwdg7MhoOpJ/7HlgzkwTorgCFNUAVEh9Df4woEvzjYE33DlCrsOP7qVDX0
ZnRZy68EsJqrGfurJY/yMuzzjwVina8reaxKCnNw/xtcBCpqgI8vK6/s+mzGNSZpviyGJnU22ul5
Qp2ZBTjT1LJ3SvqdwdmXBkVW9Zhuk+7LdCWs17rIWyX+3JOGXoQcC2JqytJBKiww2IuLmFm5/Gdh
vqXpKSc6AW76ngIG44lYkXIlHxf2AO50CffI7dYarVBSIx3lGEi99GlCNpyqMJAG42F0HUiDefdk
bke7Yg/KoikyWDUr95HuHnchPacb6ZzY/TAOCwLUmesJTUJdBMu07HJF2VqOdmK/bdIfmRgngsvO
yxOFmw6hjsAqAX5flYPXPRtreywsBp0WWgNL/YcIi/fBBur78LxizZXXfRk7MHN/UbxJ3wQZKMa6
61MB7gjgM3dhOntM9mM8HAiJZ9MndsQ1lk2xnEe9ab/gHe0hnbJJCFUxeQ+C3eRU7kPnxJM0sSM1
hA2p0S1xIv5EdcSttQPIe8+GjMjlbsIWXwLNFp5IMkO72c9kEdQx0edC5jeP34IIgxN2sGW6G76w
ZGJcNoN6oWOJ/Cjym9ith0XKVxwwqK8Hp0JnybnMmo0QbnJIW/Wv6NDtvaPUVxlJxAjiwMu/S4A2
LKkb5tZJP66itCPsERMheR/9PPny0uKB0gM9xPq8Caq30gDFTzg4y9NpdSoXfDg8DjxOREztZ95r
VvcIGDLvyyCeQnpijWQXYAz8BbMlFtEgPA2471LRY1F+TQkiqgH02uYn50+DmQQS4aMkvCSUIX1E
S0tZnwsyKXrDW9C/tIlSQt20T+43QBTmMhmNiFwapLoSDAdMwNYq6bLdvcY4BadB5T8TKADxrli1
lLGi8u//IWwXMboDVfhpp/i9Ob2383gOd9P9iQhfNWFZwKYthCm1b5ocYjllW4tcq3mHnt4UGcT/
O2MY6v09tby/cDd/2srWLA3ITZXN2LCkWUbLL/vjQkCM/c1vMvP5u3iUu+UxxlO5sYjjPO43e6TT
gGrN27qB1Vmfb1lnTqG+5X6nlZTpkbwi+TId3U0Dy0iCiPhD3l+J7H3Gn5HB/CwAtCHdFdOMwh2z
07e3CsNxY5jseg8z2OG9lYfZ9XMcNcYtV1J6sp2iCeecod2rn8+UhMkkB/lgT7KxzLInL19I+yk6
YAte1o8gyh+f8LIZ6UBTcIIfQsf3c5dP4t4oiD5bVftHgx9q5+pSnX2yo7QVtOZP87VFAABi61uK
eLrh0Vohn+FyPUCFke35xsQiIC9R7I7xRy/OSw2Dl8PI6vevox6Fg4gLLy4uxr+R2z5fsa6Xd75w
3ytetFlCN4R2JqMsXu54luGfzezu+OAwbLptGrceP9JJUqQODz0qqepdEs1aArQNKE6uiZ1IBD2D
No9yjtYAqlNJXgLyBfAIiiE295JjtehsgJAwKhbwAqF5KryAAn4CiJKAOrQ51TZeukMehPSLrh4i
w66L46sxbX612J9S4eU424dX0uBuWsxwpc41CeH7Xpl6PukFywBCsjUM7j0he/1H8jK5iEjk8FOV
5A7U4rtUbbgzyS/ViuucNXLBbcQS57sSpVPxRaVgOaq1I1X6e/7d8CqzVpY6GL7Qg2Di+RSWTN+i
qd13Y4dSROenbObp6YElLwW+N2CDve1qO6ahIkDCxQ54It88Ds9CyGLUhx4OeVFQQPqssvxoCpyT
sj8EMHXKItntfyHft/oq4rF10tjk57Z7uJ5+q2kk4bFYm9vVVFRgTcyuYI+rZ+Sr96Oja9YKpJnL
0HdpI9iEASMl8f2hfBvD8C+4NONisM1JuTSL/3pElMRGRooGTxHhIpYK6lyNWIg9t4D3R8frgRRu
8lG3D6HsIBO7KXVjm44yKvp6c+Qa/KuVOGJZsfZ5nT9M3TV2YCBy8VLYWlantKdK4iXqWTTalcG4
0+a8o3mSDk4esYHZua6VVIOHlc8N9homqYS6uFmqM1dDY1ReqQidTz7iyg7sz6/BPWHNSQoBNV7R
s1FLHKM/iWhlRwEzB0AdWT0nDP0sPDv3YkBmQtP7Xxua45Yf6Do4MeKk7bz04K5voXSKTBz7vnue
gj8OjSYd+DOjGBSQv4kX0kxpkRmK5TRj3nVvcOMU3OYubPijbdsJXeWxJwUsuSNdZw1nVsHUMFz0
eDUCKECPNYNPBa1E1zr1/MFHjs+4ZW4nXFR3zP3tT1OFWy10T2SsCW0Z5fv2wmqdsQJYVuHDDdkH
byT7C4PgMdJ1KtwTqp4Dj6+AuAwpYVKiDctp4+Pnll3989Pzd4yq1MfeamD4a9GAvgY/j0cFR44q
5Nu42UXBPXw9z1X2nv1i3YSsspqzgjR1x3RG8bABv0V0+okjigwr+rLyqPcv382pglqIqfL3dVrx
UP1K6Dv6/ZbKjX8UeGeE5FXaNWIuj6aym5Pi9vgHrCnqX+2jb5f9SLfHYcPJ//5opvMlCp+siOuC
1/QYJ9dH1yoyyyqrVoCopmVyMPn/rT5aKbhnOqIGDRRYPsRB2sFlA0JL/+8wvj/2hoUqUK2yLL7p
HGy5KSbknCciuXLBtrsn7xDenrjpQ4/OEWxFNfJ3jJWV5mdrxK/itufnYJ0edIO2QJRXbUeFD04m
r5irG8fAXR5iyuMhMB3BVgH9NI5fImc3UWDtrWStwiMBuWk0I/Otwnjf2V1AzJKWPixK1DBN/p4W
h24q2srZbl6yWbfWk+Gzhxpw3NRhvjqYmQqHxVPtuw+sybn2M+GKcce6d8DY7Gq0/Nfw5OdjBWVX
MOc9JRf0lUwjM15p0es8H83kREFerbDzVcIBhH5tZI/J6YY86rpjH9u2FQ6xIh7tyUg3eePaLqj6
sgQLOwRtqI0OHpkIZY3G3fJ+BXH66TBy9K4EfznTs3t2fmNKMOcLmio2yu9H1Q8DgE6dCielkfR6
y2lqqN11x8Za41tBbIzEARuqV9e+LugeFopO7Le5A4DHZWGuuuK4cEg6nB+y1toOlVDWxo1k3LYH
Y4gAdxFdJuE4Sys7DcoyR/FU3XSvzm2PMHbOFNmeLvUlLfxo8CmpA5SKZFGsVRq5/IgwNXyfkJDU
3YO8migBaJo/HOQqWEaTmirXdqdNzFdWuiIFqc96C2Q/z16vg5MgMR6PwWfJJEJnI8yJ+S4hfj9W
9/FLXUmFP8J81yI+qoNYVkdIKEUvT0qkeGExcO3+/Id6X8igdwEO7YGk6a1QG1npqh8wLDfOrWvB
jLow7kyc2y5kHo1pUylpF+hp1K/QNV/Ai0uVQ4o7kBTCLK3jF+zxBK+XZVDq2qIm2ADYWT8LJQ2Z
nV7dFBLTWUxntra6o1xpakp2/DClCxb0LOhjFhBKwPAZ7OXdxbIO4WvJ3F2Rt6Zv+vV0/gn/J1B0
b208aiLN/nKYwfqzSELYimMfu4wZHPGZtn0dyJVt4NLFBw0SJtLBMXvPB9Qv8R0fRIDaQLwuvcQc
qZDgBVaRSXPSNLYEyzxEtd5XCRHZ6Yc3bKzsN2gplQzQR9swPlUz62grI2TOXwdqyZCB1e0aCoxT
kVKcNZkeV7VDsE6GNy0H+1noXhzN9UtnlzXZTwXKcOCKiDcv/i3kSpWgQfVr8Qf5RubnDLDWX4YU
Z8Kmoty0s2Hvv3bWfcuMtTokqDpxGjJft1GJwBwVUhNF+s1xD9tBj+A0cV5KP26TUKVuWg/S6Lfc
2qd/ZwAFBfOobxytopNuS/rC7d45m2z+yg5MClW5PDOFfhLqI1UWNPyABtetaboMwZk+OdFY1XGA
cHGOtOu3ONu+8Jp70I9c+Yrs5N7hc9jGGn5vrHF3P9rEQelM9pBg7HRGdpTw1YfbP11TfYYmm38S
uoJHH9ex4pYJWwAd+GEbWUH+VFugCHa9HG412mxbW2VGAZvr1uhiF+cbYbRMoJm4Zpio4eCRQVzd
BSn6KPxebqQskqEE5J4IK9ScySxcVOA4T9o8zLwKMhRjN1YoM3dWnj37mFvnhXfyjzAA1DtZXQmC
uPWjxQ2nurtJYmO1kJGjlgJpWQEa9ewCfGFtbpH74w614o+f1l6V6QICobIJE4rGyIWC5I/Tb28W
+93eV+Ru2zLB4sC1s99bbSgOWI6eyuEluKwoZknNQ8LYqoxdg6rUQIOS3TnvmhoSVnsDLHrFTiFJ
FG/yXM2P9Rq4VcNb2B+GkzmSf2bf+kQhcSP/Zg22LiHAX1bF+9X7JCcMCGHBpcPJwAGesfpuqtsf
7jgtCxDnRkluhL02U5O7dmsndWKhWB6CvjTskJ7Mn+rDVXeiVFgpqH6OeXAdg8M7PQyq9o5HtCPE
yiWnspjDx8WCxBmG4Q1ZhynrbU4GOSGo2LvWZX2hIk+SGa2The1VLaOzxBiAgGYIXRGtxH8HFj11
UH856FPvLbUxK4faxf2jJ89CvaaHDwt1/yCcMZzPFfKy9HY8lh7ms96HmY9aITE5POaLcya81CYY
JzgcjcX4t3SH9AFiph2fmAmYyatXnGaQaP0IumP9qDRAUrTG9VTa/7zQxl9nPqI+w94Qs43Qbxiv
fR26OhP4fbMErxIv2ntOFiDymIDpAAX9jojuOjPdLFRjnU2OrlHMZPDN0SccbP3V9037lD4iUAMp
liFb4eGLdexyoIPiBAd7NmgJ+DKO3fdOnGvOOCaolN8WAR+TQAixjplAA54nYe+p08mj2TjltVYy
tojqjiw7bvmzqlu6Q9WX4WIp8lrATnBUtygXSmKiqfJNl5Ca2wNA2nUhsifgKL6wX97dlsU91px5
M/yrq6SPfAbayjflyiXzH+eXK29JAPwAusTDYyeJVuWPEmScb2QuG62nDb/Pltjwphm4dmHbZZp4
D4eDmt25ZYAzynbyzXz6E0GAOsss4FxfkdOvqpl6FSF5nqqYKevmbDH1l/s8hr4tq3/GF8qQvevC
zGu+uG3AeeoXb0bYSuAFbj68NTvTgEL7h5Or/ICibehIhBtQCbfboVtr07/OhXTtaCMUjD00d+5u
tmQzOcdtq0NUkOuwcrzr9e7tUZWdpC4S3mJZL3yn4oM3TLOLrVV6IVqa6BjyQbKboKbRXdSVjWyl
mR+gC5vBOa5M1HNzN1usXfUVfqKcOof2vk/TO3+plqttgH0wZdxHR/U8OZ1xoGTUKvkhkQ20jnpZ
0zp8/XvLxEM+vDnF+FmoJJKTc9J6U9jVwc8BLNY5smUsqPIAxS278FhZql/7AGtvC/2ci3GOG95B
n0qAYzPcVTJhamv+bFHabITMnefB9QCrFauqnBRISh5s46r/NDfbkn1dEl1LNVIIiJaqBgQioWCd
vZVe4CXZ2lP4YFlJHlmuiy9cK97ljFNw1vh1CkyaSR5qbTzFOJqM26Y3a2xILV2uj6aYsw5WwgtU
6G1gTu3KttbM/5R6uGOGtluubTrRTKHhNthitmGJHzMZbKJjQlEWeh163TV4kRBlmA+JrTrGrPEQ
4o7DjbcTtoPcdnmEHoRUnOrwaRLyksDxro25mpJri4DC0bbVa32lilspwW9nsBEL4hcQxMUiskAm
lsAMmwxZNF9WZ5a8nI3IRmeqIfWmdYVPen+9Ou9XW9mmTuU8Hv/YBLE8DtKFVqi6bTg/UWgvWvdN
3Xg+QbrOsDejsFXGf6QplibI9eFtKX2lVodDGE0GBu+wdLUkSmN6IGHdQyU3xqziaz2LvyIuoCfw
BYrRIFyj3HKneZlehpk9BvvX+XP/vbs7q/4Yoc+xCDvyrm6DN1bpkH9sqHnyqOirCV0DtxghfTF3
7s8sNLxiDDIVdnkxNYj4Hwm4+Rc9PQWEmcHglWPjhByaILOeoeWEZz/Lz4933QdjvBUoGY9Wfj+I
v4dj727/TwmhOyGzbzqQKK600sz4vgC/T2eZ32NexmYP/YuoEpOvAhPf/xwZXoZxlXKDq/37uPOr
nH6dWPoNB+bpCQQ3amfVNSk3mTueFTJw9aEFCy4s30NOYqa64/xFZpi51se7msksMBoYTPrMuOIc
ZYGog2naIXIbY2acy0x10FNmK2jIDSzUFaYX9DsEC9QqtLrHOVn+sSTx6b06lCIhWHv5JBOEslZL
oKmE3KBI3bimckd1aQO3ZkFdQ6SqjTamRvQwKbmQbyB5l4lQ+G19D043Qvv+aiod/Umr1kyW8QRK
XiwuWOxU5djl6IpSr7HhuYu+HmLiDVPEVndsM0xd4BK39R30npcVEYQG1whv40P6MV6y7C/IgwRh
YWhcXlJsM/CW519eR0dF1d7BIroI1bLEU6g1In/uLlM2HUxTLhL9kk7sCXihfSscYlLXyu3i7PoK
Zt1J1rtTf0VoFfH3owI07aUBz68HekSjVsk2ORUzvr5aXZi7NIVnNLd+4hU1RVZgAPCF3wNBgJG0
YBJdrzgCANCQqD24Spz8oyNI40tfMQuyajI5SEtwujI6aQfP6Kvh1XdD9igmoVVJp6l7Pf9tu8vV
wZyyTQ3iAIt8I59JihvqFlEWyl2Fx9n1Gs2HVkwvjdulmwKvfba/Fz+06O1LFJxjChTwvyrPc1zw
31InQtNwWBU5HM3BMKH2fqESjVkQiwD+JEDWmO5U7jw5ZsHwJoa5NtIWQ/JukHKtJBQgGk3TZ5Sq
6Yg+zDwniGlpT8wkSIdx0HY2ZWuXYp8rZBmZhTdc0GssY8KZ5bjrOU2W33FdzjrbaZuWAw7lh8yV
XcXgYMv+lFYzGNosSGZxmUw2m0dZku4Zc6iNOFdgQABY+/2IcKdUTFjUA+fjrmYEo9kRdvWeaxeE
N/nWbpJx6Fh8IntiIV/Lc++9HAoVqNKvmJoP14PiiEZsLNjlVGPlsPwdJ3+r548w9RW/vDdi7E8L
nrVuE5188HoVKzcjRNC5ZkmgwIyD2AKErsexIwGboc7S2jZ4bnBKKbhmBDJCXZ8wRdtkUY83Ya9a
mPZUyp8Hf/+htTCyPoNBT3GSt+0hKXerPBDegj0yFZrrwSha9V93eO9yTsw4TERCDU5QolRnL2j2
rbZlUoLiRaOszTRuAeRGPgHTY43JSH2CvpiPdIN0/2iOXHbI8a/lXCHB9l5RFsjZqqI+KqvXhPJU
Ya49meAv4w3B7ojfzwCY7Ye+zKQeXvTnsOiJRb699BNZ5Dey49tCWotpz3i6f7/9+mB+Fmrq79Gu
GsBWxgcXvyrsHrD5PPE4sLm55nMzNG1Qa5VyRghnPeGGMpQUbOpPf93FqOeQEaBRz2G6aJ3Oyl8q
y16GmGtrGM81qSnM/E5XcnDpGwOBJcXItoyp9ibBkvUV3M+bo/tYPCl9uZnfLS+n7s2+3FUP7YDj
NMDC80Sx+Xnp+zeRMw+F8T4xwPCfyVzuGLR3cfkYzOlkcBZ9ee4cblNdO4ZX3Jo2MK/Dz5Ql95qR
OBGjrh4rLWEvd9SbzPYFczaqjZelJuqMY9wWZUhb43tXtCott7aSPfRF6ArLrcaKPi5nnVPJQoK3
L1ssnLAeDDeS7ef1Vw5jSEauPmdnNiYlcR5cg/NKMqdWOociAIA5odAmmBDVTzS3tmSsqlfFd7Oy
cRLe7mSv4Ag9YCGPPJ3eMEXoF8gTJnwlh4yF9NMgELA+/tDFicbpVs+xAUKjWfDR8IWqhguzzjqb
r0b4Zg7l3dtB7lHtP08hYXCHUQFIZQW8TOl5OC1H7sEtg28rgEtVNsLnvWRR2Oo5L4Tzb+6gaA2r
aNinXlhroHo1tO75n4h9lv2vR8GjkLjErm/KciA2+Zq2PMlV7t4ybr4lgPMXdbNO9Z8GrFh7NElH
AVBUKk7phUQ/QR+05f+dsDstCjFWQVDg85TkLzvwZnJK4qEUG/GDRxhAexwhlAnQk+y+FKcyIDBs
skDwvEBYC5mRsIhJBnreO7U5MTqHKz6vek9ZAgpK1g0NtWwjpxAYkSKLvUU4SUNlzGHA3i0PjlGP
PqH8jY/ZcuxoctI5D/Cp3iFDwB4ZS/lGpMLjUqdWnMWLfUM7pJS0eej/4OpMTrVQR4LN/jteRQzP
NsYUQnCaXgQQbWSPPyZ58xO1DTaVLjrryc7QlxHzH4Q3N8zKdefhXXZss09J7DsuWU5Z9waR8lWX
gtn/imqMAEimZaqu4lE6+UvUJ04OKbFa6u/73r01otmFQ4UVaqQ/67UKB4qKVMPzwl2DuAozAOFc
HDAzS+2QX5bSj58TXGzCpSU+8A/UoZnKIQOlVo9nNz3RmzMVx4+iL1ENAYGx1P0vATT9Y41I5l4s
Grv/2L6r5mqumCalmK4kn7td26wC7TwyaBxQaOhAJM/P+ASEmpcd/B4l5d0Lzm91/kCtLH9OVgA6
Nond/nI/0xidSTo55hAPqL1CCsUE/xcnxHo6sy3CewzEJSYOw+eqasZ1cnKgN9ZMq17qKcTfyFT4
H82lu+crZM+Whp4eDOFQyPnZ1j+hnHV8hXkg3uLmggW0Re/bx1NoM/WqXZPiHqBlvKqOXLSoFha4
GFPYf/HhdsZPyfWWW5nAuqEjc8/TwGg29YpOXvLTsuFDNLb/pB+6HylhceOOYjhLLZAX+FW4Ma55
7jkoa3HK+ANznFW+OnelQl+rPli9mwR3qyiIzgnJh1De9w23IMhvA8/7iti04IUYuE+WeTQzkUsP
IZwpmR7KZxcaGQU4TZUbe0RSJyaUh6oNQ3Onb4sFzHkAHOCNw1Zjk+9DxMS0BHMA4Sd6lb+1ZFCC
IZBN8+ZrtndAl3ZoAQdW2l5DvX6paR3OQjjTKyCH+WCbyZABKDOZAwio9CP0QtwlONV0gJXts8RM
0BupW5NNrD5oWwsqiEjXj73k2IX8t07R/tSnH3cM83YrzSKJdk2CSVNoFxAziGnHqy8VdUtluJCa
0RSB4bzp1WQP2cYR65Qt+mG0AwW0dOXLJpf8kOAfkhu9RUZsvn+4ZTkfObfgOHnx0If6ImRszVNW
76WUWjjfP8y/Dkb7/FLHZhKu2ggJrs2kX++ahXBZeyAgi4kl6ImDJtIEAsCc+EYKycAlkNkwWiE+
vGAt4raj2nqKNa/SH+hi6SDNk7VEKB4f73BIfrJR+FYIt5Xnyjmhv4LiFC/589p/RgJyTyl+d5rw
b/Jd9Conz8i+WF9aUJJ3IY8cC3drQ1Wwe9n7dqBaJ14DjGAyeEZEQ+VCtkuofPQInZt0NiBLvTA7
z0+dRK35o4Xjea9AQBhKK3EBftD6lNHOtP3TlsJB1cYGCOXqR2bTsNYxiXQfGTruNX6LjQrSepko
HOPAOdfZ5Fy4Arifbr5h0ynr0DQMwrCJFKsfR5p90V5BJRj0MhwG0hSVSElrhTeaAGLArmMIRIg7
7eAGH83S72P0f63MzvEBCHaFV3IYA7D1ONIF8Lz26A7bHWRqpWMa9zyOb7qWDQgJ2ZZRkhsnVg3Z
8YC+wIwuJzGUUYswIFe9AhpXWz+sw7nChwV1XXFu6gaqNhevKZB2+Sd1Jj5L4MKnegC5dWaoPpYQ
SDIJjlnjiE343u3cg3PztwPerDJhHLDQQ5lBGvS7vmnERhhaNW1dBqBtEB5Q2Yo3H3w/IloDwVKh
zKl77I4QmpCGSuUJ1z7+suew3hyir2L3Nboux25II8AJDwr+1zS7iwLseE7k/hDWB4CSCTdFvhIt
/thUQv8jJ7Bd8hgpst0afvjjiE9AX7srNIRnKSiJj1jIQw8+Gx18DdUD2ecfFmE0lwnhMjcsh81t
Sp6Gj9mr5eO4T1GrIcoFUylDCP2PBuTQn8KD+TAbWW8RMD1cwXvSd1l3pIYlltUkY/Blh1lRYYnS
r4waHGVYeiRbyc06j0fAlDqTkXF+++/o1AZFq3tAyoT7xHQNviK08hdetdggxFlEUvQoD+Sr60CL
ic8M0HAlilA1fVrQ2muNiR+u0RAG6125vzbZzsMicJ5vGjSzjQpglvIuq+WJu/qs8MZeuC1k5LtN
iKUyCO62c5eA6a8UYWeo7ghDS9coSIFXbJqBqv3NZVuq58hzk4XfomY+7bg9cZuV+x9jkxweoJUC
e56hIuJGRfAwdTkq5iJ0LJW1+GO1Drl3Fb9vk7xu37pNvH4i/rFPqvfx0ItbbG3uHVMOZ3HtoYex
vmXqrd+WASc99bU61aLcmA1vAQs4Zw3orttBQGK20y3t6API9L+STrlDpWhxQoCEjj5bNffeTFt1
AAo7oobwQTqwAFzZGNqffnYpP+ZwpZBPwuXmhHc1KDMv373UOJgxgMk/uMReV/ms0ffFAgRGJdCe
UF9cmec9bZJA4snTZjehdpN4iLnV8Se7N4sB8IPw46iPT++WQ/CBn2vkdWMVKJpcu4fSPumnxe4X
BG+HYBzTe7Ds7B/8h4SYnZLJ995hDjPnAPuuyRV8DeChJjSCL05RLA/poso2A7rTqxWvJEv4FAME
HCpUc4Ee+jqbaxDy83lw2MZ8y6ckdFKz6ZujE6L5jTaUcxltYUmHAvX4L3VdW7Z4M4Q88vsdsDnm
ug6h9cO6S7EGza2nCSyAhfW9oaHx7pHZiuGS2VQgPFm5nZynuh3AoMo8hk2iKKeVSFxZRe+xN3JJ
GAeCc7iT7+esWoennVsmQuV1g7KBS5IMJv5DwFj4IvWMw/LLnChGCIVm8vxoz29xuDKu39KIy58h
MkZ9KpITtsQoFxbj8RW//F1za9dr+v2AHM96BVmgzivyHxRjXhbXeX0S7UVgZFqG3mpBfHe+Pnc5
md/BIHcwR3FpkfYyWDphLlNc0OPDy0c2ilHUjPiASHlXC/PB+aeENCHT8NFyAu7dUQNVWshcrj7G
BLZR0UOLYefWbne66w+4XmGimS6H8U8hsoYRBykzQIvXulYKb645wrLuVv0NABjRN94WkJgmzUeJ
vkzgV/jUR8YlmwKgLpUdv+fcPeFL1gYhj8GUz2Ksc3D3DKAxW/xkfBspeCDJyTGAiQ1d7eVYDNha
RAewX9B8rW6v6UK8s6D8IvPP6rb6ZsGE9zr0J4+aDgtFlotXRgbYncFG/sAB5wTSmwDpbWju7JK3
+mk+4tv6YSN3cAvlRiooo/nKnyC9pafnyrDAmiDEo95nOZqKkB6OBcUzZTMVhLsenzVBy8oJ++pq
IGhiPX4ubGnSB0MPuQk0CY9yteuGfAl/fzA0uI9jGTWBzhzFWzWo9mhcNRTFG7IpaQOlBKtSsdvX
/FIUviIP1aMXVbv5jnwFi/5s8qAO2oQhvenqrfFi11VwMTjZ++PuqSogv4iuBfG4YoBNIT0bYSwz
mc4IF+ul1jpSQlU15+8BYS7pIaqrqpr5hC0PcVrI1dqTlW+z/r6SavSZyxW4R3byCeo3tq0px3lq
b9QOqdne8Anssm/exR6YEMiiOW5ej25yw9B+qJwCHcgGdjPwmsBEUX7HgHObc0fYWBy3gRNmeVyL
f00HdvVPZw/UkuJOwVy7jtQPEjqrRPsNbejxzeZI4I7z3huAAycIGcK4YX3CpS3f7RCefBB5zBHf
90m9H4r9QtyrcT6rOcSXcVSRE9/2AbI5/11ScPnPB8SxQEAchWotE+9OMCxaaTMRQWa6ZP9IAb8Z
hyhbfX0LKg6KaHjeUa4uE2FHvLtWna9GTSUBGztyoNzaZHJ9vfVqDrtPR2FZ9lkK11sogdYYkd7w
kaTZEJf54Ho72wQJBKMoNEGpdTLVjbC2iBs06/fByGQVg642W8H6bm53qmF3H9hcU8EaO937ObPU
G+xI00qgffPIGpI2fAhz3oyyBcVEUTqze+Kjx3jYzqMFcw9NxnvliwQZYXQ2W3ET007GKvIAw6rM
Om/UM0B3OxX4MQlUeVAqQvuYUzj8yhDgZmWffOH/2h4+pKFCdIULuOsG+uHIy6KyBzPNK54oTqmQ
3cOWoqP/M4aGNLXlBSeYGLDAZqs7AVfKuvQKEDoa4ogrwlGl1F9s4Me9VeUtYVbaW0DQpwkrcjWg
pwd2rBauDnZ3DEl+eGOFWwd+UbGwWmwouuFAiOr84gJMPxdlQwOU53v1jU4bxVcJvafnaNQpI0ZQ
5+mPJZFptE8ceWNEHHR7V450gMsB8XvlSxPQM2gRWEYaj/tj/m5PvQgs4NC2REJe/ITs0yBmPb2V
se6WfSkGiWbzq8KXpx5feF6lz4AlmHaJcnDoJ2NSo5Nz9LAlsaPA1ln1xnWt9VQxU38qd7z9jPzF
ziy1/ExV05AoQ1Rcfu3Bb/o5r4qWOX7QQfSea465QMOOL05b7a/cna3QYOfTav1icFnnypCsB7NY
V0U5BNThas1ame9hTt+mOW36Pu1JnQzHwuDjGOFie5zrM72cnDZniexDJx05e6FG1fiTrXtCq38y
/uI21z/rT2te5B7lOMjBEzgwt3rjxIErcrxoMuZitdJKut1eM3X1Vi+2fdO2yauBoLwwCp79+VAc
FQM/opKha/tb4cIl5yJYio90OsGJf0W2Tm0OD0lAHmYwA9MGY8J0gESnnOfCbLPoFF28+SV1WaxG
hJmtVmYz11S2kMtsjqgJWzBiLtkRVrijd9YgWP/I1e1f0VXYVGZmCLFlYJU1n28YVQ6FxcI4VYnW
XBaffk0OhwezF3sHDOyynodWSqN1RicHlOSR1NV+4CiH1uAnAiM8+onPkrRoxa0ueJWz4ET2nZxA
NKvIk1AhcbOti5Sn+v2PvS8dcyyJhYCZnAHMqOE7B0qb5LknG92K4/akpblK6D7pNHifTwGBIhta
JnosvZbFZGlbo7V0k1S+7HFT5gJMyrKG/DImyNr/m3afnQYUNgGWXI/vev5A+bvn+Md8wvlOHbOz
siAlyEeM4wRBFI7Y4H9cGEnKTI1ltNklGR0qqNg5PkzJkKegzSz0iNoXinENNcURLDEa0WsEd50U
ndHDnjGsAzBpGZxEXyyWwt2OLW5zi3bzpC8PQC7ZsRz2cHEgArXPeBiwI6IRje9DN2M2Ge4oF4oH
EwVac/Kq+j0x47eyc/Jh7ax7OyQyOlvP261apw2HCk6rsPWBsBxuK7hby3zi4hrfJg4CTV7Ywmv8
J5CQf99/rWCceteDwwipeUQ0DlQvJ5UGpeNP2sEX35lFRQ3u4cdTAc7esq/E5Fcvd3xTK/ahPXEs
Z816TTR1pO7kTmLu401a4guA1KRhumi/VRLzdMGRjG6Rl6YzDQ4rMP/DuAPdWNmwjzs4+dLoDKLY
3BGJ5rzvzEWkDJdHdRqC3PCyVr2PnqZlu+OSKLpoQWriW8WLIoQR+ZoKGnyfktgQYaCEP3qFwVPi
6k9wulzvM2yHbh2+wmyV1nB2spAoO64hi4KvIOPuHA+PpS56V9s6T1CUzhCNtsgwFMrb8VDjgWq8
pgf4moXEBhiYXzZmKx3cgAbuJwe8/SmmmW3Jh88uSwUUaWW1z/2gdBh2RvFr+5c7+iFOZGOXuVaQ
8/kWXF+P9x7QmTCwEjEvKXr6XIXUCXTJedWxzQnrRaGLq22tp6s+CCnLduDMc1EETV6TwmQ/zbbP
vHMTSCHJ5W+KQTRXlKUo1mcjKUTa5UbElBVZjxa0GS2uBgqDUktCZZcDntCVXiXVZ/gT6+hudwn7
bpNnyXy/4rtNcE6Vb9g9Gx2XCKzLEliy15navbqgfhjHWkLMH/ZVVHwvi57wxYTKv6WLJDawMuXg
CEHmvk5ffyvnrBwmU6cabiSSdV6qwAn6KnIB0dcf1bh9YDLPoUWPY3WKAHhJKNVIceEhfYlco6it
TpMioX03sGcQdOBhtX2ZREBpZoOgx8Y1iPhcdfXRlx5I6dmGmbqxMTeEwnHomCO1kLOr/2lZkhZH
BRV3cx0otGEIsFFQz9N4QoocyY/TYS8xrOJNaQQQZOVTuv7+a1t9GF5diC3eOoyEMaOT0qu/jPVk
jdJ3in8+RbT7crIDIN9ny+oziLuDHxzh9yWQFlLJSoDa6TXBAsc3DDuhvwQOGDhxg6RVNGjIU4S9
f3f9nRcj+EGkMywzB9Jd0rgK+6AdPCu6ZCQyPaNn8QXNfQ+XKq4zhffgNvHtlWwaUdEGed4yg/5x
zx8/VRefDdgq10Mfkl1wLrAmzHdBIJd3VPFkIcgBu3xYU57PafgLbgexEHvrxvQvJOKAReasnIjZ
tvNjhhPfXNNc/nyMJ49B5xNMT6Gy++u8w5YR8DRqc6bGLgrQZ2b59Bw3V+1aXIvgqmt09sZeSkZm
Kn91baCWKeY90XLbDmIP9gZ3EWyeiopQ4uTaGKxZorT7d5AleY80HE7+i8JjfvSUPxQse2cPlimA
lgWScsIQRU1anGdE6b57sXsvvrBEj6B7iz/s2caOHqUx1ByORloTkdnAviwox5f0h0T2syqluGJK
jHeX/9L0dDysKoCZatux+ujP9mOhACNozWIDC+g5O4OzZitFb9iZXcKiaprAZU8pLOoZ/iArDOfl
l6WAnVlKNs4nlpx+8QBY1HpuMnQVnWPcwEK3v3p6NHaZ+xy1mfzxjZwomZsk33fsHxPSMVZu6MQz
1mqRqvSw4HhCogTvNupR2btdp0aYYKbyxQbcG/0f1tUO+Z1NH64QeNTfbcEatyqaSJj7vS8FiLNz
rgrsrLvxPAmpgCoZi0ihKrPObV5goN915IgyhA73MtTvv6egrlJPJbTEabdIYoK9WSaeAWCB0BP8
QwcU0MeXYazfDssbyeutHKY+7MUfnLmL0HcYacUI1+qLjOtcXvRTZmbN8PE/+wMw39HntKnMG7kr
r69qSdNHo6B0Tt4Pttrrivz2/zHCX+3Mu2ClD1szd7SIQOCXcE2yn8niUdRYMKt032ZC/rCtPbhX
e7e8o6XYf39UBXqcZY4mN2lwyyIG9tty6npXQdxLDh2agUa8ZLkdYiv6F/D8yiQON/E6TthC7Iw3
8hD4QdwY1QIjNVN7w7h1N5FLmecYBEnbi9e4pceCdUHJcwyahkZtZYfxB6euvLXjv5qwMgjin+kZ
OQy+TLlrXxEsK2VUecFr5nuXuQQNQaPwB1vd+Bo3uYgx1789bHp/d18F9a5qpriAr7de+zA0DVS6
tuJ4U/1Rg9RjHROCtJd8LdZf/lpPt/pBcgED5KDd4zCB9Ec8DowRzDcD6B3cFCYILm8soYyDZbkk
q8WiZnfFcrvsP2fp26TjK7q5rxpTL9dKHNLkJRh7na4myw4wBu3KBxosNCVKuS4iV9yKiTFMHEbL
4qSpC3l3NftqQZwFvOr/IhdVSvCYuo7XXROI/yERopUjj2Sp6dJ+/7c20klMJDd0WAIRYALfX6WM
deHKQj7XkYKxKTpm/KryAtnx1+yVZdtmqTRJG/6FCvAG/EI8GoUXO4381oTpwaNQDkJzDF1twyii
G4f4oEBJHMC6eoBRHAboIBLEUfiPjIwHar0DdqnhZIu/d6b6+y4lzxTa6EIM2Tkreslq0TCDYfOQ
Ezt6rH+5IChoyKDRrjmzvkO8oRrR2bzr6OuHEAa6CPYOIKFXp2v3/a4sMB47XTyK03huq/JNzWwS
IKLrRWl48TUQRbWVmxsHHtUDBsMZzWHaYn0biEfbxJmWDiJGKYeEKqN7lfrowJ9wWgGPuzgFpnPs
zSc+/0B03Ps+3yATjF3DL3oZhriet7Wr5WzVbBE2Ynd3ygobYVuXGWtGMxkZYu8Bi7wH/QxDYL9f
iSPeoNymuaE/5ePcD2vvXfEXoHtlj+2+q2mYhZLnrW8zXZtGaP0Ne76yMiAGdDqzCdPj+zmghgNr
vz3aYc+lywrhR/UTX5aXqFeA6OUxCXVjZwMyALJGpUu59umFsQYh15db2XXNMXH46ORmbsLDdSCT
Sh+o1HRrD4Cvrn1RQIURGuQJ680rC87zusXlwbjyd39LVZMDlj+IVVWqamLEtB67UdMAfmIDeDb1
DNzn2aiDtSYU8NRPmO88F2zjqc0iU0fI+I+xOsOuEOzG+JZBZhke5yYEqesBs3VuBgUwCMeL6fND
HPuclcL++64133LldYqGNn34SoGjs1DPGdmgacu14Awx7xQoGf23WMySxixuqQMa37EEXk0Ks66E
N0Ib8fT/zbt4zxoxYFy9jpHJCiCRABd/43ZeNF+nZmdbpfnNwdoXaFk4umHy2cZAWTMWCFtbitvA
9+mWjIv2Ukrlj4Brws6DNs6oZbaTY0GxkHIB98UVuG94FXLKS882ep/13MBGUr57OvqKvW4htDRI
71on++kFkG3qzlEVwT4qKp4OOdqb+dp7dFWUAFJJ7+lnjU1mMGxWqPllqrpbo+XSTTH7QPO5c4W9
zbbulK2WOElvKcSySIJUS7Vi+KFxky4SFcd6FsErUJ0QkeRgcn/pcn5Y/GPx8FMrTVXM6kHCRA36
RXmi6HL3fOhoNfJzU3pjYpxRwj922VdmkKbq0VoruschYLD3tG5PQaYo21ocmNflkm2MUTHs0jOs
o1xkFk2H/w8H/KhKivzurRCTJzfTw4kK9j/hA7ZIDDhTEnSG7dGOdsW01Gx1XVr3OZZKcVl8jJSU
cm5ccona7UCApHZRHIXfjyKKTF+iILKNS8W9GoYgvhVIyWlBrO98L0wMqItVgd0+O97xPi8Vm/jU
5yPMOw2OX2BaMFx+GXUeEFcTbQILeugPxrExqNqoB4bivnqpwQj9ZiCacdGAENhs5XJdZ0ST4SZm
bSlMQeUoQDERFj0CJbkhhJXpS+ZUC86ZXW+p2/X41kOQx//UfRJaTKGPBht6anUT1IgPKTKQ35p9
R/T7ElbbITVXx/v+8dR+6ZJ9/nUIh8bGoIXEoY6EHyb3RctQfYUD2jKnk95pIIkXWpxnbSN/B6Jr
ej30vpicfPASC1guEp7M4Djme0ULhjdfa8tndsno9Z6b8hEt9L8ZxScqd9SLX6D67DAps/C0bjnb
ChFv4/q2ItyEAhfXm9UYz0NSWQsBBDw+2H+i4bTHNFPdinohIEE2rDe9cdB8qcK0jBb+9vCwPPNA
jWaUAJqSs9Qc74HKFd/FBPLHeAS9KOopcjYBrd9YjhPCwwtta3g65mKK+ZPQNY/ZhdqJdorbelmJ
dZluWUOM46myA1pQDvUFBkdDtLuJcyIE2KOjO7YGHog0amCaS31lfgBGs/tQ24bTrwOvojt5+hIz
ks9/8nvxck4dGp1PLljnBl/EwZTIcUCtfoNcoCBByDMcZY30rq2PJms++IE1QwVkfx+KZtbfoJbB
Cy54Mdqf0yI0P0I8gs/H72OehIwtWfVBFxxgzS2TpSWyN53plNp7Ffu29TMkaPOZ9V9t1I9Zx5Xp
iVClBCpRa1+OD6kCjycQE6SkYlPs3t2FHcfwHz65BeHz2sTgDJ48h1a/qHeantda9A33QgkvRco7
f7C5Eo5THzquanFJL7OHDhx8QcGnFfKnP5luiTUTOAYtxazYIYu8+RnnFtFGhs2WmYBuiJ7EcUZR
Nalg+HrJDCxNVi9G6HG8C5femJ3ZLPdRmZ2Be3sR7nGk/3wHAjTD4mK6dVZs7NjVt1CMttoECWvs
U2Bpr+vFsNqhxYnUQyUvAA7y/6AekjtnahwxPB7qB+M6G46mcGeUWayorXyxXP2bFPTrNy3GV6R1
N7mc4FpKt8yLWjs8aRSF4SacA/bUsJQNHHM+hLKuRkyQ9oG3mf0nYxw0Sxl1jmilziFuAiU5qmeK
xxpFTo7ZFSirj1LIYPtiDbFz/zFKI5QOW7l3sZT1jPiUbPGbj8wSCfwDN3XvEumaVXo7BiGHOLvR
xD8yiRgNYjNnFJvEKfG/l/D31shSZcZkz/MJYm2pCBwSB4aBjCGljIsYbgIvCi6HCXub2bawpLae
OlLVEym8ksO17bSZ+KfVoylrxbUlq8XLerEfqylVdUD34vXBLk4sNl6K/esfuMTJm3w8o00CIvHe
wd0kgmrE3MjPDvhSbusflw8ptB9LpRfysmYLAEx8lKBnoR8OtjYHKXxtAYS2m83/dgg0u3eFcCcO
1d+yth4+/EDrDugQ1kIN9ZG8jKdkbB+Cj1HjHPd8fTzsWaYtU0jPZOIJ0N7aIndJpUtX7YfANFJu
/oYiS836WaS4kEs6qMTNMJ0WnVo1Dxc+RqKe5Di43VIm2tfjm+v8QXIQ3q+npXC5b7OIqvP53YpJ
MWisD4vdU6w6QDmZJe0WHdtAQkf1fqIlJoCvuPzV1f5A1W91e8WhvklnaP+tYFdNyur93w8mbzz8
UXInV4VQyDNcqHS29OEoieBxGjUzPv+AUGCyIWR7OxXut5Ek85otHV29dELQsOnuaKGQTF8uyWe9
Gmfjp6MRWdB1MAaQuHYCskJnggG1Iv7k/cjnCRguAxF/Mc+q+/LkLQrYylji/9FJ3hqiV7vNzBWh
mtH2lFgqZT31lbF6ofXBAt6GL7G60dW1rptVAGxjqiaVAcDF9TUD8t0EPSQLl/FShZ+aS4SOrZYy
WzSDqUMxlCRN7Ec2Y2gPgnJ5+TGE1CgR2EO6zR4Uo6ov/eczU/RgSEhuKtuXfO+I6ffx9i3rDeLl
y0NpGwbYhN9SXidEdc7LsaIUwUBJqYyNXHj03LizE1M/Kj9ZXSNoe56UsEbow0RwtjuCQ0UoKfk8
sTbv4ibaWDZTss4CU9AehEvv5vqBD7f8P/SMPeyzE/MvJttPbtdxWBeuKPDLxzOqt+sYiN6CQiGi
/hrevmxlUwcbcobIg+5hvELm3tNaZtQuXC6qcU86VL8zptp/saQsfJp7LBoTVNYCqIc9CK5zZWnU
usYEB1bOT7zGlGZVbuat3sYvCR/5Eo2y4Cy+yTltJ48tDmoTJRDxBFIqzXT9Sv7b4Fya9P5/Ysig
dIxuMVSoUobsiJrC98NWetqOf3ruWlngUohEYXTyFL224gVTcpdGJR+J3L7Zuvj7nMwqhNrSVT4V
/lfTdFKSLHw2fLfWO5kmNIe5AdgQk1KpTJW/fkzAr+mzMn2cj7jwuYNAEgWSnj2B1YkPEHPKq+tA
wc97dl4FcwZmLT0lrV9iTCB7LNRxw0D9wxX2iXBE4/EYsvgAmv2dUnD+eLlzlvfrj3fM6/z+aK/W
xF9i3C9r3DmAyEsEnYqJeLauP2F250ZNyEheqvmLZ4DQClkz02C9/Xb4dGMwbzjWoVaK9OdIiXmh
bVXZeB/3gXEX/GUOhfVznIITpS1MTcRhVXpbKIMlDJSsEY3/yboOcD/21x8YWJVTjh1ZqBURkTq9
O48qz0wGXKbdzPF4FYtB43darm+prMCI3FfpqwtJERNhphey36+LZ/jfw+SLdJAdxhRfGkyiRjdg
LuBWsfU4gNWLxW9XjtJHwdROGjnsC1JVJP74HoOQ4EY9jquUSbmFR8xpOZELB1pv32HT4SgpTia+
ZagX/dmYBPzWfBx/pZsk5flRjb+O2MJRpYDjPb/Q8QQ8mhDrBahNbz9Qoupn+jtemEMXmzOsfniN
AWzNhi/ElaCOpyaecw/bGOrL9SF8DI/WhrEkuR+PQk+MJdTerNwpXr6+JIFaXGbq0AuNwNdjj8mn
Hw8ZhWmjV2VmQQJ4ibTs1+sgO2A5bKMPzr96Yqm5uC5nfJMfxdsvQedWd/zck9h815i5mlz9WP6V
o1NrUk2qf2zN+0e7+fo69j9ZsCvMET1zxZEpv8mWRrdqhAlum3RRVRLiQ1qJxOrP1dnJC2WZgO7h
ZTZTzgmnFBZjk4e2XURgL+iDI/yE2vBmGdAnSSEnh7uif4CuvtWHfsdxUlenBX34XrxelaoIYj52
AxKBn1bd3TFNi3LyCdzHskv40eF7ETzUQBnEJqBna686sEN5bZ3lckCV6tsKQaX1vKY8O4AJ1vS5
Wb9Lh8GbSYO96cjgTz9kFCMn+u98P1YSVN6RKZvJ/XymzZiJmb9MsMqBdIWXILZZWZE+wMYIHMCH
G+9LKKQdfxHHgvQY/gAj1ZleGv7hagHBXGZO4ker5VWJVA3kMWbFIQRO4e4xEI5IJ4JcjkctbX9P
DI8aP6EwksRV+HmtiSnL11zlL1F9VR08h4wAC6wi3Ig7g2zDSvkogLHbQXJtYAwwfoPRpGiuiN4D
1jz8bZfiE+Ol5APXEor3rl9zc9m4mZQpw2yeSLBYp59jgIdtDHJu/wXPOaf1CVsEY0AknVnjN12/
FXN1M7HPRSwKmQ39ZipV3Rw0XUxX2W88SClLFYQ55ec/iLKP7DFVrHTubmY0GldLNEKpS+sNdGdd
Ykrla9L2YHAo6uSaz9TAgqC302wHxS+GZlll6rcIWMckEd7yeVLLZdNYIJEfgM7gvZGROr2u8tLx
O1i9OVcn39jmOi3WI4t4iApwBYg3eERdwyxpfSjmPBNqiLecEaXxUAKZ1ND9Lpf9g/8cf8kJcTSD
j8Lrg+R8mgXxg44OXaZRbHxKtiggcb4Rh79bJatOUUAqxu6iM6LJlafyHHEn9MD/dde1XE6Twn+E
J+dXEvdl3LvZbJyiHNptWNhWVgz1zT1tYDYq1Wgws7/M4zneGIw9Y/39MZdNplMTcK0V03m5rBC8
zFbkgvVNUtF1zoCRg5lJQ0MfyD+CW/uJnJkqKzC7k0ifWcgQEhw7IGpSLxije0hVM4ovMSg1sRYN
TRt9Ygfw8ZKw6X1QO2KWtCAqbV9a7WoRQmE1m+GI4U+lT+ewGCkRIpoB+e5yP4IAHlloxTWf7/St
bitOX36R6ye/86BvTMFZ/xsFR1X0QL/Ts2XrdBonFxki4gGrIBETR1RchlcH2aObFUN06TDTTykx
rwtj+IiLmlnwEhXVZ1ndqj1ELkVpkqtl/LVFCO+EQzr+vwL0u9Jz+0zQEoLnyDgT/X42hZ4bK3sU
AUpflzD/3Z1053Rq7alFF18kgcB22z9x4TrrfogBgU4Py5zVMMguROKvpHFSOMgq0As2x+aQRNuV
QvSpEKTpdn1pY+3rTOQW0al/8xsnr5wcN9Q32Qt24QmoZA/crjBEzmvKLcP3o7jGHv1V1t2LHJuS
a4C+PNBjTK782X1PEp7M3wP2wrZTynZmcE7tyor8BCFLM2shT0wc5H4ib/HOm1v9cU22JkARpe5o
C2qWra7SGHbtZ6sCgHI+EFKtyK24aCgSp9c3eh4kPhnHc9TwkBr3ThZ4K6a2i2Ua0Q+CuW6nPTCX
v5MtQYZof4KNSe5a37qNklH6Rptz8qBSVrLayw3ThrQ+yoITQQQ3vX/K7ziOvfyf8qyaAjRiITjL
GYK05+Zl3ZKnnB4994DW3HrgV60xbFG4bwsMpCH8GAHlDpb7ibAwsxm3JtS26p25rSR6b6V48Tc2
93ff1QYt6J+hI3fRof0iZdL8cCH+ASLU5GOlxCiVh7ftFHN/4lBlbi2azWjYxIRe7/Xzn0vRtFQb
UU/pnQ33Lx2AhMhgIwvsIZlKcs81q9mJkZblRS+FgTlcF+JbOYKyOfEpNzJaLKBeoSX5wwzrrO2i
PSfHEzeEKTldbymxiUBTKVvy7LnGbhGtltLdA6Nb0SZVittqPq+bF0hwFVQGfeO47lJ345Hwnhb8
Js7FSU1YSKzc0d1bH3QaA8kY8QjdvLROwqV0Ihg1DvzJxYvvzd5rWAz8TLlTC8YyJxciJuAIYdMz
i/QYPaDQ6kj0BczcbLRyXzio4ccrOz6rDvjH1ruCLkPmZLwQvZ+yew74l6SF5zkpQj7xgN6ITFHc
o3V4v+VKHAH+dE4yTjO6dcE56D8RF+nCVzHZLNxLNcssCt9N58OKwopwIkJrCiDgIAG1eWwl1tem
yC6GisqIfw5KR4V+Nuk0SyMoOZou8WZHnv5/FWIrzMsNh50Ql3brALiiOGhawEMWZn3wPnwIu9Pj
MReU6/hANd2GGuyuVtrp3LDsLZ5WdvvzDatTfuqXtmEgskJsVT43BR9X/nVtB1eqwTCy5AhptZ35
e9oSBFwjXNR2QKa0VRMJZ2p543ps95iRQ40nXHytNqBRXH1DwR0r+pzQNvSs3+z8R+9ckEOB37Ho
8K/r3PyoXzRrn5Y47n7bACtzjXFeiA9zG9T/TYJC/8f6NyZB5yJbLiAJc5rCoOe6e/IbdyloT5sI
aHEvlBMXSX+fkmIP0LV3H1jSG7Dd6zfP03ZznJ/YeuF7Lq2NuofPCXV3bI6QVPDjaFhuoW5NIlpk
zWlKCnToTLzmXuK4W/BQyN0zs40OdFgS2whkBMoGat2u9BdURdemRGnlrX3CTLJKye7beCPzW9oA
hFnc5ogMwsD6Ln0S3l+shrVM0gvrRJeYY9nNzDoNfyfs+uX9DFYGh7XSqxcHatozJN06+XnJbBSi
8W6AjV3ABufqmCVI9KaMjjd5JFXcNFCkCkvH+PfBya76nDcYwfqwVUEEs/eUS941N7sQ2dloRtNG
aSoydkmAvDOhaqhVSH4awN0GEgjLLd21hUIQsr7FZ/XNK6cnVDFesaDgTtXYguoZjtmHVLLUKLfN
+0VGbxBpcMnMFC4tZDJ2Dsb3QSrEs10jhox0ACBlFTbOJanpT4e/8z4wZrq+PCklm/rlEe6blKKX
u2uw2L1s4RMFb6B98QDVnwnZY1Lk+6HYA3toYVD3mb8GbStMbJBKWoA8VKmbDgXfypp5anpoucen
EpMAXA98zSNVqqhcrmMk+lqIKsdF3GYprJ+PBVeeh24QieJePZf3ieKTlcKVd+X8cOYoZ1bYujrC
ly2S1VDLOtlnEIyMoFJCbRf87/GKHNP8eDjK+XiN6FRZYylKbuBbSQpvla3bpw3ivwA5cGYqUC+x
iSiDy/DhNrsyhYE3fsJXYYg6tweAPuaNt/giY/SLfOTvncdo8+ILCHcPak1ui+kadguKIBTENL1E
FgKN8FfrFX80xKvus83FWXiH0oHbEnvcfLGR/qA7bikctAz/b+zMSQnAoukOa29KriDYADimo7B7
YtEnAsWnFhB0e2TRpz74QBifNaqxejL3q9hOeRPVBTF5mQOnLqfwGuaWZ1dm7+M6TCoxeajNxzpe
MkLwEewC6Ucp7U48CvX36+4aoIRSqzfImfnxYOlV4LXAfnBdG7GHyPaOwM8AdcAzmjXeJWgpqbfG
mn2f+/Tlpp0QUIl2h26rUVh5YlPX7f28f4i7hV6gtTE15z/9ZYbBrasvd7onSOUhFiyU0BfpYHx8
UQslMjXJ4Vb7JpV0kgyALqkCmk3OIx/CiRAgRrhjo5uAU2KP+UyTmgwdwBZcabznMnM4C1J8+/1v
5sCHMyZACD8aiP8bunH2p+OHdYs3d8hhzvxBbuAWUmopvs6StBX69MnqOz06NkL8Vpl1fOqBNVsd
qxfco3s8THePPOfgsXIVGo/T3RlI4XY00yaMz0Sv/xW+oFSG8iNcULjSqa77odGfkAMzAxdGnKVT
h+ywuplRgb860xNH9x2J8LKjWXfcsiWJzR7cjkHwLDEsYnSHKDijFsm1lUOjeHZrQsyNsbyfAP6G
kV6hlSRZl1wH+YOPlMrLXE8DibJ82ZXSok1CtgtxZ4+x+mqr0aihB622sTDYWhbiLKBoeDsOfylT
hK3YsHlFRV95FPI7OUxicYsEfiosVT7fCAhRiUyCS6ypBrYFyM2hjEyIlTZXQXBDclwv5zevUijn
aD+e715XTi/5nOYwluA2OCHtXOL8/e1HDegGfDmiyR7/nXrBtuAlXiL2URhO7+5R0UG0UARjOAg/
4M48AwHdc1JMy+QSIBExoX6XDCvCYeYhuiXuVGTeF6ZIMDO2MSIJa2yD4UCwLJy/hNKL/ICmL8G3
Pm5yBejuexaGrl4v2zHaIKMMHL2ozNxyLO5qTWG4N9gmX8cKwro47KmvJDbymOK8IT6euazHBprk
6a0Z5MtrzdDr4EJP2KFTX9IDrdS2FGp3zhfHOgGa5zrFsb1HBCGaEGIbNEryA/gghpbcg2PH1oIv
ktC0dgnWc26gPafLwca2znV8i4V/kHURWigGlnN2vgh6/KHT6BI8Xspn9nq0nTIniKnP3CEp7mZF
mOsfQQhIp0piWC0sq40uzZR5N8ul1ipDBJBSWmRGslyO62l9q2z6eTgb/Doxy5mwYTidTCy7Qm6H
y5p1wMxQJUaG5218vpHfeoJajnbh65v9uaeYHstim7pu2zedS7TvPadI19RYqhn05aCd3HfTHTfr
QHq5h/IzqmzCec3uJHDL/dstK6LT64E++oMHrYBnXbMM3iwuMPv438eQ3R0XmDqHNb3h5Dc3GHJc
2pArc9XmYq4j+2iWmU+8ARYCl/xrxLonJo8mOKFmrQ0ln6cNEoDmg5rfYihoMtV+F778Z+ciBfUd
PJcu7JeFMhlhdembv9EgzB1kvr8z9Eh5l4ZwNcwyEL9EJqi3sujh/T7PSykRmO53Wegy+eVmQj0p
OB7dDIwcwJmAVnA507nG7NQk8E3MbvpoCL4Nxsj1LA+GmpVJdIRCK6QxcPU7JoNG499a3FQ2BVIq
lnCHv9PdFWRhdsX0Uo1VSKd6sr8TK/75/w7A9NWRqIxSSFkNglLnRJZ5JR/X8dlScmmosO/APyr+
yR53aIKYNsbhPIaryW+7AMtHIlCh3zqrjEWztZepNC7845T6P1Q63/uQJTFS4ro1S8UCLTzDvAWj
ufJOHBlGYFMb1eqMlViD8w6kncnTEhvRCL/BJTGexdlts1KrZh0ydeNqNFpB68UPVrsJYOceEQNx
LS4vImliH1B1D3H098mH3Ks4Oz2nwNYnXvvhyzqYUEoPWfqC4crdumAlTjMO8a8eHOR38RAG1DY6
knFzXP79KnMEhr8+XXDPdUPi9OEGbCgc7K9V8p2L3C6gCNiXbRNCWzF79UK1OltcFd6/ycQjQ7j7
nFMiHoFhGGhzX//oMJbqe7ZeQyBd2C8XWF3EHObo7WTBc7AvL7ARkWpREIB+Co1cBn//shupfb5H
RsJ9lAtBxaaRQiHpLs9AS8jxepmmQMuhoRPF8BmrJ5Pa+Kd2yQQXrpu2UXdtdUiVSkXrYVtd3MHY
bL6rvFWNA8WoM0tdGjltRUc7XZaagb0I426R+Gi8RrW0cX8TvRrh9WRPbOH0DV3NJayCUXqv9PDE
pZv9Ci1J5KAFI2bx20AJKAPgQDpqCpHUfBnOI4TJKpVgHuUFMlDJk7g4fyY0zbouQ0bmBCnM7d7j
uuJZlJ/0m6tDm7kCWh0RMm3ud5CqFAeetzu9ZD2ipQAW2VQC6w/fN7pc2Jm9dVMp2x7L4xBV2u/C
PuKpl/XGheVUsQCkQdD3h4ynpoieTi9hbJ7sod0sFVb5TVXoSgVWIj/YewxnQHpjY1iipYhWYf5F
/e8PERGaMOBQWvau5urJHazl+1JrKPMBYsBI+tzhLvPpTQ/3UKiLxOFLwcSoc+Qy1lfX9L5RI4J4
2Mw8WXfPEry97k0E0xMK61qf6T3nOo1htYsh9ySWU6Px17D7I7qsRVxhFtbdhhv81c5vvH0+wIrd
UQu2o6qqfoQC43dpZ2oi5tv+LIHcwhjiyXVXhpUGwEW36iz+VW6Bful+ve8Kd5o+UchrprfLw866
Rn3mugEtU5XKPNzdngdPRg0e5jndZD+mQRiAwSCq4DMV3d7WUQoFWkRYimTraaKyK7WlrU4ikM4/
CsqZ0hxX5ikj2yWmEQGKl0y3ABKJxA+LNwVEIfyxx0N9f7DU5E4+CAeIFWz+Rnljsm+T5UuyIWz3
ZQ7xvahbgAabsw6oxG9OOxq+Eqm14t+19NM9R2NTV+9lbTgbNyqzOoFOZCw9HiPYKpI6pGn8ODcs
XEcrLfIZMMUk3YmGkxgRT/IKk1wtoFqWtwJAbRKblqs45/3BTJpdkkhIStb/F4F+kp+qP+twi4/V
l0ZcwaT9Wr9KFwAtCOHc7DmFyYDdwDwgol3wGr61+ed/OYMilrZFTUi3fiBQc+FXGOQm5BhDZAYb
Yo4tu3h1/h0Qos8kRuvPqAJTct+tL6ye7VOdezkBKHe7iU50NSW6U8WnGmnwl8rvM08ylrsa4g4B
N6U4RRMIdxYcCQwWyqJDUjo7j3rfnBG0paI0/GIwc1IYZx3UWU6uNAaH+5FOMeJyvDOv8dPjSTLI
JuWbre57GYPCECtxDNk8W9wqlGWYvZHmXm9/reZwc9VpkIcXy47y0lc0nAGq9Jx3K38CeyVdo2Ei
35it0y1FOU/QZTlDZTS41+f9mJ4q7bGblNOT1YAY7kSstMMFBk3H2SEE84i3J3wnVUDjjtvl4WCv
sRmPUUCk7kCII1SXovFrhGROaxKXWgTf2+WPhQE3LAIMJjBnJ10DA4xhZywkViS/GoQ2sMBI7fV7
1xkR1cP2WWqQgpkoy4KQhMJ/4hmue+DAQNlxLpxXJBx1jsgcl3WHugDR1REuGT91K2FpSeeWrho0
bNnhh5YlVFDS7sP7QVMLHtGm6HT9jtxFDiE6gYQgHtaYKh3xL7g1Qq9duP6FUEaBW/BtC6gsHNQl
GV4sY5POAlkWobxNPzLuzeWujLDSKy+mOH3ozFsBXb6kDdFo5g4/O1zTSIYfbedropnZjuP71zK3
Pj+ltZVDfKwc/nFsaERYankmjvYKXnJJH967w/tbTiRx9dn5evNAawhYhsMlueWLNY1A8+XcSjEB
Ay1tIZM0AQJIi0wS/m+L3s2xWfs2TQau9JMDezH8SAUibYDlkGoWSW/Jash5Z8R2YwWsH5lPl8AG
N0JDmD5R81KVKq/YlsTOmeKvTImq8BPVNEjHhXdYqls/xjLy5Ixj+QHi3zLVJmaWX3Eb1iW0zQAU
mcrTuIn4+iWc/QZlHhET5ZknBDUktACTLjFHYAdHrTD9wVLoC/SDftr/Zvt7SAErfdjHW4uDgoKp
xHFtjNkaZT1canzqTzhN0+li92tjY+Bv+PyYy4eSBN/kbdCaLUPhk38/2oeDEVEGQMwd7sGURk2x
2O1QLIIldi8DT+jQlagQeRHfIQLmaQXh+J3iqCzpEa8GE0Gn95F3ypx50uHpNXRr3O0J6xPAkfC9
GeghgPyaZojYP4n22+3x0XPOlKn1tgndYEDkglN+1mFhGaZcsf9lySmu1YD8rU9GpTHXzScntu6F
OIh3/LSj2zcuEcyJ6OW6Gr6BeK8HGGwXoWBBk06upAyMybGKpIdTBFkf8Zj9gHMA2L4iowUeDUYQ
BoPBUnB4FTmgaFzXUGS7abkkGa4/ojLATCZrt4RpXHrlRVhVi7C6oRn6rGe7inlFrNYi44DaOyia
pj1zHAEeDvMYaPdk5ABItDm1VJV4rkJgsuMFWm1F3DxJK7CNRicK9oU3ABq5hoFiWR67q5sj67m1
rq7QJlj9V7W+wCCZFAX7lbJgPecZT7YMKyGixgW61ZXr9LuZ/Aqv4OjVvVhdGD7yTGZ9L+Qu98gK
XdeCU5TUCukLSPl89L9/PUSof6z5ZQB91mazBH27D0YwCaXJ5ttw4TTzQFxc0U2M3Uv5s+eAfnKS
g6E/b/kCgWf/jX0TA/JX5yyw1YRkdehsYyvMday/pUShPN9ana5MP7hzejk1Bb5yqNGQNCrnlIPI
VUoyuQT/N5BUh4Xa4G5wGOdIgGHvknkGjm6mJy5+ukUK67mb3yO+Ty7HFPRdLDQGpdxlKhhbnIdf
B2dJVyWZomyeZhGzihn1V/9DkIYtanfx5dm6kMedex77fyVkWC/ozGnaekc9HW1fzu77gdgtgLnp
+PPPYWLfiDs1YcOqixWlFkYD1hL/NRwB/P681NvqrjQaR7KE+IAfosErH4XKnx4tE+xLtGHt5qXP
r4LW2pyszQaE84UXLmrMr1UUi+LgOBc7KgtYL3yUhM2ZDX4C8eaOXmcoaDvr7POk3VmASuy4CB3c
QC+nEMbbUM+vVWF2qae8ch2GCKQ3rsdoxOIDuDU4FjPrZvbU6e/mRVeDVyoSgIZ/ob2eTIph/fFV
jMOYgIW0delMetPNQfFvmH57MpBH28MxXBVknZtHQkEXU8bSW9M3QVlnWkQKI/U/lUdx2wxpqedx
/kmZIhwNpqMVdyNJGFHepQvh3MjIoaTqdSgMQmCPce+kG6bXe8wAEkrjVOOeyy3JEcp/2EozmSxY
pBtNNjsfXGcqjQ8QM36xlkg982Smi1lsrlnRK7t7BdlisDzlLm3meNwPSPbWzNNLX07mucFfonXZ
Gmvwio1JdlZAOl9hrNaZmd0kwaxfLuccDmtW7bRldqtzqTkY0x/QmS6C/CoabpmKfI6DqkT7V1Ed
r0UsYHqEV5lbQrp1Q8uyuQJ7uTSjjkg0l6p61yM+TZk4assmRHd8+cUI+Uo8N34olC24d6rDSsZW
t42BNKzavcNNrcBlnAPwJMDnhRkD5qWRPMFeE02OEyuWOVuFQooDBLHuk3klgIQ0Iwd1aw16iOgj
R3lKgagtzYwp4Hp7w3GN1rneBTYKQJqH/tVSJAwo88PJHuCLKSOeT4Q3/LCzgQOf4JxRHmU+1UBZ
7gSzwYnDGAVs5QSwAL33uS4yhHVLAThMvTt5xTsYH5HdB6qOfrVRBZBJxrfYXvM87k2n36KiCThu
/mJFGOc+OrD3dffE5uR48jnRHIJFp/5csClGY6gMRfsVlHSAD5SEHj+2gLHfDnuwMznloQ+6pQ4A
XS+ilYVK8JKy43Vnxz4JMfW+Dqa9yLcLtEO/UH1ljD6Y2l9DsMKvAfgYJ4aV6KpUjy+HaxAtRSu/
tfHv6UpmgplhlC2Dtjj3Feh0eHzxpJUkk0/a1/p2K9PdVhuGebSYISLgD9BApj3Toy2abF9XHctw
iLJqVBmDDosuiKhXV1gXhU2pbZD5brijiaTJ2aNEBmZj/5oiKRrG+V4C0GJseu2Okw/Yap6HqMWZ
0wh8LEl+EnUxSyCB+QiTQVEshhb+EuJHFnISl5s0KDhSfIkAOyqyW5HdoWlmnOrZvr9/MHK4K9DE
waHN9t0BUA28PiSEtzcMP4DGcdsYoZBGqSGxNUpVEkAHMjLxjPY92KY5AS74eJgNfQ6zYjzBb1ho
2oTGyjr3nQ12EDThknzL49nVAgzk3aBDQeLmBfFmRJhI2dh3nA2FqBTY69H3KxZn3z/Hpyd2BJTE
HiHRAyOYjMucAaAdr6uwQwM41YV7hbyyUr5RZle+05kLVQ5ltUfn1Urw8PpKfJqCWkXNwpVnov4H
FlNCZaVfJNn15NDkci3Hzfzf7jR3aMzbYxI7k5dLWUva+CKHBKlMHmtYVHmTa55N0XvVxNitLJVy
5qDzRzjmUHUPFdXetd4zw8ps7J4hXXb4tFPrncdWRpw0tk05ElOxUOMmXoo9ga/MEdMTRdLtl3R+
aXJJsQegE1nWgVJ4Xs6towgDHw8YE3maI3cC1l60tjNQhDrrXfDRP/+o6mFtZpwc4mA9nBbrMvVm
GfHeqiJn3rvgKP325kkpy/++QHqqrdlbX+7vwER99b3CNhovjkHxRsINzmHus5/N2QX9+HDTB0g1
RXV63eJb5c6C4kHlVh+8EA8AQ6/WYOlVMs7cZjl60HiMZ6/dxrW28YmJnTYKHTHe8FSYApwSDsHK
ccXXGtrB/aQyg1SQqmS+OW0/Z0ktZpSVExYHCP2tWTGyTDEmiTYanMIr53HS3ZNyc45L3VtQEcQA
7tVxZola9G/FUfUIPUrJjN42t+JV5oBjCRogf+V7wNx6YAAbNcWjyLRcUAqx/m7dUTSqHxRN/f+u
OwNxKOoHXwP4jxKSkEGdHI1Wvmb7TAUiulHIl7zLj3Vvj9AmBUWjJqgc3TYMEGYgUneuWdpkEtjx
fjWHHvRdymQkURXaKam9/9xiXNYjKB22oiuQ15vjdJIQIDOn/ImmiYEL5K2kZplYNBANxjRJ156G
vBg0mtK3KWb6K9GM9uoFn7FFJYhm2TG95VcQlAg3WXbfPJRM4tlqFCh/IW4Gfhi7Iz6jcVVv9K4S
DgZJi0tQg4dYr4sInjlnKLj1ji71PHYaghpcrnlaYvxB746s+G6HJMLgJer7Xw7c5Aju0ydh4yNa
5iezyh0sfYZVZ62Moqo9QBZ8G6b/r5ovt6OJF8BRffExxgm80CLK43kBt8ldYZR1XhlE6lcwj8Hf
9v0kviWCNMtdunbcXQavqNvP5vq+Wp7nBXUaT6CEdn7Xn8v2XIcpnnuW7BH/fiPv/2EmKRrfd2to
8XLPghJKxojffasrADB36UcTm5QAOAyk8yW0HWnekwpxyXNyE7Vqu2CsYnOKcvpakkZpIG8XYmdU
FCBSTSur32WZQdm46bRhhAtJL5rcCplOAHdk83iwxyxagkeDmgX1J1++wxvtNUnOQo/lsLjTFpP+
GBOpGSbXiZmmLthtXKGt3LuIb1PaZJiHaAAKv7BHXf9iQz9nW1gYHHgLSBY0AsOdAbZLFsFtcPU3
tow1Hlj26w9HUzHUsZkLKT3jL6CH1D5LuPpieuhO2M5ni/rtsFRtcAw7891drSkPKPQSKq38A5yu
SFZCNLLZYv2rvOiA8ppykToVw3kDLm8mFCKA5r2pFggUJUKcsMFhS9X85VfBVZWv4xDP3NUb65Gr
91AlNMuQU86p+pLAIWWfASYyVM3brmmZNpFh8BLU7Y2CctY1cmhOpBx6GKvNu248rIA6IbrHnPHE
aiFOYmBFjMxPeiB382pOj1kX9JNoYyTRsRXd/uj0oMCIt0ZvnX/xopSA3I9eQAPCIjV/FfVaiG6z
0XfebQpw23WHLuexEgtDT9lxIw8Ftdn8UCc4iyAuiQ4u1sTSAbxiMH7FnnWWqGBGyf2xpp7PiRej
zLjo4Zbdz2HQgGy9p3nYGWD1iATf9AuTp88aRjsTJbn7svI9rCNa6hdn8h4BlE/AeYt2Gf2Lb08v
NLtjiYiywt/dogSbgCxPw8kEBcSXYMU0EvF2J+DA1Aj7ESgPF27XeX59XRbIdeFfI7tKCPeYWr0t
FuUkHH8XIJcVlieDZiKG1h+U6Dbw4qyeV3k3LygBP2C2IBHPSiklmSZlyQOUbfprdoIJG5lZlnwR
fGlvQsrzay/oeese/cMsBtJyAsci2/qwi4dBZIEy3csnvJQrK4Xp4pBT88H7lkbITSU2m8TUJmh8
VOPa0inDvCUW7zjd070BUbLrYp8BJPfFXzbfZnFussPp2f7vqon64NZGo2XHaGaCnx44wauUaiz0
aupSzJTG140DER1vhl+B4E85NdgMrA5lqhcf1Y7TjanqHrFaU7ZfySmk8muWGQeK2OiBb/67hVYF
HuB+83nrnoV2sTae6uRXCf6TC3brQmuUuPI9e/bKcJOM16GJczNZUnq+3aJTrY5Sq9mzfnoFqHoW
3bPJtJfjLONAwegiv0mpJUwlGSJ46/Dy6Avq81qFBf/+A26i582r/qMjyHBAO+tskPkBizf4osK7
370xWk+JppUyuc2Kui0GMsnjhWoYZoDh19rfyzE2xMfWOUu0Jb42qvlJLolsYifhQc2YuItBl2iy
SN9K+u5qeLFrJhRwYpLxtr4Ewcezvj/OSLYGw6bVsFA8ubsKA8neaZTgUEHWTuPL2dxX4tzDpT66
5AfCpTP8t3C43DTi5dfDk5n0BEdqVKbFcU+VAXNQwsetUqe1EcbfLLSSIrM/PQmylVQE0yBqrtHt
1p9I3TRbf9im30Vvzl1ku7ebpm6egGc+7DMixESqkGlyIKN633YpYfPsvnNQEMJQYxJiqs/3O0di
u+SF3fdSUJiYgXw/r2ocB/9uorHUkFCHmXNtxGQ6N7fxdPgPTkOExP7FK3BvRPyZ/mVrgqPblbfU
ZerBN+o/twrrWC4/5oDzIbSafFRlfk1Mp3VrXwMLZINdDdBeoJTPnA53ru0Sr7D2AM+E5OjXUkFV
hINLOm1p+uGiMpeoRGCTXJvHE8t3ciZ9sfsiwsbj93T/O4krKoJNOESK4AFiTG7xq+7nTkzM+MyC
VPpeAVxYA7nb0REBWw/DXgu3bjLgCGqiv2BsQWrZhW5t5SXRrLvSGdKWrWrqoRaSEkbRfSXybf2p
8UIJZoy4jam8AMJ5SVN03m6j6HEnmEtfcdWr5NBsf5qC62J3MrF/8m6gxCCJKvXnH9570Sr8rgkc
9EW7ZWMi/KE7uAltqUNf8/vN6FF8kGaWkRpvzJn8P9tVLhT1zwrWzGO1U8eKQXItU9ef/BzQPgM7
Vwy02KWBCsqfpNWI8mOPQBjFEB7voA9WQQqQAEvQ5NtBuTQhcRibsTEMF+wUMa4HUT1NWsbLw3YL
4/WbfMvanfcinw58WmyG0WRoIyyZ0xJvXVU4Q3owRi/I2TWcJ2pyHxjz1OdI+CnqGGQkuzKQWphK
aHcDX96rNPsnCzelvFU16kndYomhp2oKnVnjGK3Oz60ON7fZRURY+IC5sKdjcLH/Yv36qIgyFf4P
MlInHrZLiKqLbc/TR70XhYiPFXXtYVUDISpA6GQjVxhuc6pkXE3jXzw7+pqEnRWV0wLRMwmGXEpa
9FYUp8xu4cP+Zadboa31Tyxn1pc4d86qlLuxWnUpwN2N41kO9kZEbrmS/hxVLj1lNoIU8840JnDE
1lxMOpqw+9LNdhlgQEpyj+d71maU28f1/jW8VCcODFLbFXG/UbizEIEG2p1NYJqQ3Nx+HPGGSrX3
vG/Gez5Bh6n1hd7we2i/qLkc/XzBfecfGivQ7T+37FawGPNCmpBSZnzqrQfr9/A2PFHNNfk+Nbh9
ASd5Px4uflQv3++79Hq33kDDNlFPnZdUZADA/R2kEm+2cUxtzBBbfNF+KUOOkWxRMolbYnCLfeOQ
hi1bYBhGYnj/pjb8NVZHcww12wlU5oAdyGxOPzNUfO2cPTcZe99wfxYO86NZfsJN77vjCYRIf2P8
4Qiyv4OuipcpjmXKvmSeI7GS7miTi2uwUVO45cfYVW0eeQiW3TmBc38V7O87pjxCgk0nghHDBzl2
JU/s/WftY9UhG4q3skJpHmLoP/rAUUhW3PTjLLdbVWpL92WBM2hY/xX4eLV532yyq0hbfwsCQMKA
EQ3fwk4K7njD81inLv4R/jBrNBSBSLG/x6cllqvXk/1mP2oP0WPZpkCW7JlKaiQsARvjSzOglPV/
dk51JCLEYIInbaXZC/MasUVzIQKQI88SIvB70Vt2Yvq5ng53MiijJGbZ16bFoAlTPUSCvB2cDiXu
mlKzPhBMLYkrBhBTYNbuXoF2sue5iAk1skfLzNSWqn+Xo3mpGZqVp/Q7sfB7GDAh52viBmveIhSY
VPevaHicjAUrWqifgjEKe+8hkbxE8hzQHa9uLhoQtm1K5ibza6LV9AuAGA6wDzWzqFWFgFMWkQrZ
2phRqzxngT5zTIyYBpw9Dgw1ffWazzxqI0pLHdIxKxD5jxkozffLPlsy0TAirjy4FE8DUHg1A+RR
+CZXUo3v2W0OBuQ8+D3LS0uREC2D+hCYvxNli7Cs7d8FYmHQy4F7Oxm/rrkX7630cGgHe6d3rytD
E8ze0xwXoROHpa4tgqcx4EXnXBs5gFGN5bcwML/5a2k5AHP6aJZblulXzTiu8QGgCOTp9wUT+mIh
xb++5gnlXea9wZolGVGeRIW2FHpVG+ff5mRGZlKI1erA8ICJVDP84z730BrgW8meh9upJeepQmMh
04UiErLSc3auG4UpxGhcLPPiK8yxu9QCa/o8Nxjgx3qxicrmDve3Sgx8owRiKnL91WXyNcXgYpqP
dMhRqcOG6dig2WI6yZSrBPo0dKiM5wlPB7BS2WyzySsXfuKZKBn5GuMU8XuqgWd49tef8TwjdDrL
um9vTYW18ZQOXTe7G/hQppoapLFH/BgZbOsR+RSs2q8wrWSEVIk9iD/MyJ6fbM5P/oybFYcTIwEq
LuPiffDFsvIaiEQs0Ov1j6nEB3Zt8h3ot/nERGclEWYJAxVHhpL3YoPN4uPYa9H2yAEZiqNLDvox
ZRxpwbhCx+3QeJsdw+BUhtd5SdmXrld16kb8MyyaCSiIMNbRKtNViLcIEiiO39MkYN3NMhjWWDBt
7GvVa3RlPP/PcOzU4rUxjY+PX6HklmxHgGO3+0a4/cILHmioZPr6Jwlh9dr4fAxl0akm6pAL4HrZ
Ma1n/8cGODGuqwRglJ52Mg3g/TJxs//+2Y4ZGKx8dcheMhLmCAdPW+z8/lYW6vBPkSj7cF9oq4iM
FZ3Cs4zoJTBCuI1Vs3CBmxJ/SvMry2RO0FruBV38FXlHpdIsgXzXD7Eftck8fsKIo7P2AYbla1Vr
eZAbryCSG1r6zfZDGI+tFFjDjC9BcFR5Nfimwpr7QRMPy9X+bWGSZoqkEEk5dWjgJCASl38gn6IY
fl5sa85h7cFKxAQocn2nLqnShNFAAo16LwzKBxiTvKZr6+eL6H7fZeSMTERPLAWBocZCzg+qrZRC
+l1Ytswl7LA9UIs09ue6tJu++xIdjJ/+tIL4fBH7d6JYTJufYG3FrUZg8XEFd+VeWWURQAO4ZuWf
4COu9+kNmskHA3Npbz9nC23k5ayGzSVvczhoiZsGjkAPBgpmXQV7B+ZCsjsUtJk0b0UmijHHOxfw
GWUDgzPqruUCPHu7pPbL2aDhHwK5m+mOVy6vtN0arQnDfqjqAgBWlnogRYMuWpiw7yJw1g/kF0s6
VD2qRc/1kVvZ4YHU69ap+UwOskf0FsIoyfezuf3hRbKqL6wMWozBbekBQPqIteQVTEDwnE4NPVfW
OyGsa7dFEtv+VtvY7dI9me1jtLJpLg9mS91q/IxfSmCUFVhM4k4l0MfHVmxdLoDIoJjJwm1Zywlf
43/uj4Q/hz2acE8c+Wj/tycnLhrHES04dyB4Rlo03kY9letRriE3E1HcQXtuyy+p0A9+LPDMElvD
04V8/KJa5tdNzmR45zoVsIQAE3ShVUv+xJOXD9uREuIOd8cRWUeFj9FG74DUSPLl2hd273kdW1uI
3gWeaz6Is0/FRLUFptrHZM5LZXY36DNVXtqBgUSf1ydXb3Fi2wGbgagWfvDZWU8I4eL4qxD+cCLq
YSj8V9id8QPaUWaZuE8Mxl8SZx9joRsViT0iALlGQZWDuKUbdrX5y9FvasxJdQ3bD6+dmJb3D5EA
yxMD9LihdTGZzimus1ExbHjb2/J6/c8Rz7mOUe/AEDEzULWemsKhdH0tp+ipDKlIPLChGIpalfXM
uQQnrF89LbpALRVPKBKcV1PA1Fu2l5HbfriZZlpQbAeN6HQkYnTPPaK87NgOGxkFheJ8VKyklNCy
u0NaKvZ1mjQ2AJw6uraWQYDfUy8h6RDxosF3BL8tdFYWUXS8Ypx51H7dmW4TlWeKNVynX1aBJo8y
1bOcrzAh6bWLZFzirSUiG+Y6+hq96ur60nd1gRUupybfqtytxFNbCN4UB7iDUhNASbD7PYZUPOsn
YwVW8EkVlN/aPyhYTxSq6y+V5twa+oV35MFUpRidM6jQJYESUrgSsyMDyw69RpkfqZxTKS0CT/Gh
M+TsUIUb9B9gzI8Vj8otfP0Gwr954SVU8mjPWp3U1zvFJAo6gWkissU+S8pfR6tT8h3b0aJZfeuY
vRwAGWLzO6I29DW79XaPczSc1J/qFcmMvkOxS/T0nDhFMTzdHaXezZYLjCAju/i+fMhAzZ3bBp7r
YGtroAfDIIwK2V61lDDIA3Qb2VDR1bL0l58E3DTxnXL11Kc2yYR41SNmeIDP2aCvecpzbKQDmrZZ
3yC1QL0sPeqVMrwvQ5Ra0hr6P7c+/KWI1PhvX8RCdVKi0btJWmBB6WzI/uGPPcPgte4P0WJvUaCR
CzRuhgcqBYWtZzEBMy2CRUQzcYik62dkCjIJJNstTjrUkLVWoftB4n9PAAtBrvDYktVuBCHZZPzj
4bo6qZPFfh9HWr4xTe1vF/aGryrI4Vo+/FZ/Z0JbSq//SZ1Uy24H0L4CUg5LCMys/F9yVI+r2PHE
7dfWI5NM2R10uz9lVe22z7RXRbT7dVJGGP3oJoo8fsxayLntdYe+ovcxTYAjguT8C7TTWX8ht+xs
j7IOJJmEbyF7+vFpbJWR0qW9LxABW4WZBV9LXRaoS4C/GoHv4ZRePsE1xjskNB6YyRT5VaK0HpI1
H7C+gPQwFGMdxqP6+U/abj7v9O3wT9acxlyw6uIlnSZ4cEj0We5rrWup5xqDaaqZmojq3Fn2OaDN
D5+Dq3NudI9x2Sd1BsOZ6No8iDDg68/zESgBUg7FHc5V3qyXkYEGW2WxzDQeuV+WYSz/pYZu7cCZ
6vY9zehyuUN5mx4P7bFeBw7IKAJg2WmyEeIZ255OubxYPaiQTJGmVr2CEpzsH/cxPGPg8+EGdcJX
TjIst1nhZ9pnNOOJiYsieYzRzPeWfaChGfFbxP6ytmIfnHpuOQD1DV2O3eclRbMzAwOTTTQ8Yn/N
dTRR0zAn9GW6KmPpnv6CjjeXE+6556d/HNE+wrU0P4PX3W+tz9DM+09rJOAXTi8XH3ZfDrAFL34e
SXoLKQGvFlgE100PFgUe4pEhabhVyV/6RYfc6kagJ6BOzTmCds4Qa8WShardnOysl3oHViHK2eMk
MpSrNpBy/LP2uBYDQXb4d6yjJNd4+ff7S3KMj0FdwrVNR9vGEplySr5uVy6IJzEDbyHML3ETvew2
egNkj5ZH2Z5BQs6Bq8HdkOYL48lmX0vFosVO+PeHHZEwpP/XINkuSoCaU3U+L8L1JqCuEIWabU5C
hhEqmYcK93HQQxMkNM5HHSEMfQwIetgEOsv1bQclgR1C00JSosXo5NPDFVRp+ErzU2Efi5Y06I9O
2PjMy38deU6MchkCPrXDYC5sqk3c0EyJAPE5OKmr2Dt3LMNbe0K3XA4FM1GQxGzZVMAn2f9k1dX1
uj87CBUVmo+UJUBr0TBDcmv/KgGEj39br1N62uHmnHb5Q0NmjgCA0ruU2CX6NV1foo+zG1EHUJI0
AAZWeofEs4VssHx72kQOK1f73gD7RQFed7VFek7FZSMxRMw/MrHq0xenWUL2S5UvIxi25KzziR5R
1zeqBSggvwqxDciru1WyyFGI0K3VmoBqfCbtWq9eaIO+At6aN/gmQd2xp/hvZIysU6Yfuen7wJU7
NR+XiT999UWXZhoJjcj52ULkZ7tgW8MLMfxAYo46qIx3Bu2rWupuE1tv4R6xeDM+kafBDuYPqQi+
gjjhB1AtCHSOb4utr0uLMWNDcwrycWxbpABb5x36jzzsVtiCTF6HVteQF3rukdFFN3mFCVd67m4b
UCM3u/5c6Q3HmBDbCi94t19gqHinenO+c+qFlMYBOXkq8z1PZALTn3u4qbrSTCE2JuLx2KzxuE0G
HR18VSohcr16Ijh2DaW6Q0ylGas5kyJSKHQGtXzPs04SLJjAGWIl3S4RsDaW/FHFSLunBbfn5ZuS
dCs6YIBX13SUA+9CDmRAwWlKtlEnifLpDqxjyMDC29SobQku673NEPnpUgtMmBEkNEFe9l8BVRDf
fN8Bk6eHT3wn7wzfT4u2PNrZyzQzx56HlNSlDbiXc7Ha4Wj7SjOoXBZmC8M9eZNKrLW1DzMcs1Xa
5uSYrbDh3Kh/ffWcqcLW1TlPFPGtxaa7hu/bKpHiqqlS0FISPgkkFymaWeY5I9ieCSk10CpnmqkO
zWa6387zuNRgkpJyhwvMUokqsIBGkgMTiSCqo67Y77H4rISEfhrkbJAqN8Rg18AZ0ZXAj0DLKjRX
LpfdhzOHkG4AYSXHrdmGQlC8MovSqiKo1uwCbzdVgrb3ODBWBEcnZIT3m48AGuyPyVrOlIuOJ7mC
5wPfBJPe0y6UVMDWRnCX/SK0P76BoEjd8kZAalmF2S200TRl62mTBGwXKE5dM6Pa7Oi/otYgPYkt
6rhoBGcgZqRj242wINXv8Z+jv9+cCWFZ1qt+dLVdbv7awYZtpcOBPnGiERGlOPihWr7hrVCIiA1n
XJJYNTMeoTxbLd1g8v5NDJgEQp2d4nP/5xqTZlcGKLBqlhgcK8O82VH3gjYQvyU5svLIOnGMSE7I
8fZviU8DjfEdT1OZO5jBs4ifpWRaASYwkoAjeRArSZuA30pXCQdwI5Qv4a2ik5hOcnInPZu0CNbn
D2HMf56pdc0p694eq86s5W2B5/+pjogEeJnNgfeensSmEGR7bu2QppfoGSgMneUbWkvANWVQLECj
CD+b67oeDrI0HyGjY2bd9tVtdstqLLcu6Bd4YPcBp3ZL4agdctrNtIYXCrzlG5pZliJPCGhZbFOu
kFA+8WDXeDAD+NyNLAt7cr488FZLcClEUgTcr7ZlqBqCVsHHDHxBDAgeywfUBhB3D+KgmzZPKprf
/dtoSvwynhsBrPOC9dBRxClvNNF91QSx+Kx4E0ed2zgYw4YRv0mzO+INVOAeZj9hs4cdLGgi1cup
lYlu3XZ8C1sFH4KjdSt+Wq0iSFadTz+p5mDe4yg7Hr1JCHRdlk/mQd48Zv6bvFfJ0/JOPbDARTrt
25vXZMPOhaD8PO/lC8LIz+6hxNpWaB93ld1JsmCIHu1Q0GT/MGHy7UQ4wEJoGY+ob/1nECC2gbVT
nvNjAygexHfkuoKO+KXVIyxdmP6xKoNqwIP9sxTrf4VLE9B0VSqx2b1yjov48aWvJ6mMJFIvrLlY
DRmSJwCDXywkZDLku3QceYGNaNNTLJp5mtXfoVsTnQw7yqhIG+MJbOkNeDRN58btd4IpGM0n977f
ldVd5yoPxWucsV80+5IEERrqetxw0UM5r6eEuRPWpjp+pJH3oT6JJewUSihEP4omxDULKUoC3r6c
t7Iyy8C1e3Smfx02M+Jj5pi0qxH5VucNGBxtm+4yrIU9+lK6gMRiSDb3Im1Oqxl2cpKhWoqTzDfy
FlF8E47Pto2SI+eEAncQZpQqdYrlxbKcoxKD7EofB6HPMbT3z6IzGcCYahhOtFtHK+8x2JNS88LY
VEPtg1/Ny9gP0I/++p3Skmmk3L1Sl8P3SkQtSAx8LrIKoobIJ8JuqQMu/yecrzp7LIo2A8Pi3nNC
R6luYBEutbcxbTrCV6TRE9EmdZ1QzHAit7JT8UTzqbk71KxUOs8wf4487fm8t13cqZCHawmfyAnX
q36s0Eye0d/3NdJSynrzub86gyv5+g6wnn1B+bcXzR6nKER/HIgzDlGGi9LHgx17hs/6OkOtuP6m
cbVgoUS8/Yzte3fNzvxbA6ux5gqJLDfIV2SfjXtO+bws+YPXWPvVBPKVFIxXZ+P+Upz/ARO6XbiH
q8v0NZ5UhxboFA1RHbNB0xou6nmrVTJOka0WIt5NqWddcrI0Hk50xMqyFlzfk4vR1GjgSL0fwOOM
SQQOdd6ZMOg/f0gzQCEJXZT4BH4mPtpVRC7skPNYARwuStfzCHNoNdsxWGL5zjgaB32FoeWJyQJZ
LlY/plY95/aks2HcfiCO8F1qOFgHmHDZBAbI/RYa3PYwYo2qIY72xw6XIrDkTM4RbrsnuFPHzDk/
YhIfJZD+h9kwwp17CACe6f8Kz/YQFbOyel1n17gEjm0APAbk+Tt0yiMSGh5Upzq0+SWIE2VeLJ/M
p8PnkQ7UubznntjcTgbAnOK9yaRQ1hY6a533bSwFM/4Hg4Bl3+y70Py5hTB71nx1nyhm0y9Msnj2
eMAGtF6gtPLeKxaFL5uHilDUyQ+EOvUdLfdSJ+YQjIbCctB9x7godvJ26MCieArJnKwsUTy1kt22
9ph9f8f5ujojiDbpDSsV0VXqWzd6SatarM9Q0x7Wbd47JsbMxj9cqn4Ttid+3TQt9fk1MQHlTh53
dE8mM6evlcH7LFe08N6nBp1MgV8Pp0KMwSazOwXVQ6nFRuy/tb0atWLBTFXfztqDkNHRmk+hYxBd
5p6IE/ktsFUw81WBvpGHS12Fc7zikz6ZaWi4JMnEDnOSfPnSWiu7s8ODLNZv+IEVLTAfwOnjkFp9
ad1yLFCVDvyk18qsyD5M9huzwjNsTdhxp80pfNuImAk31mqtvAq+u4xwen+38awrfkMt20xfuRc2
xTEehQu/PV1RJNWYLZUMwzGfFbPoqGVNV20HqBvuSPofS8Ei+Ou9QO+HfxjkK/aTtm8EqAEPlyXu
00pXtVgfrOrpZHTz2dpDTYY9B78K33vfnFT3q+O314qdXeTggmpdC7ocUIjmqyahZaaP8jo4FH3y
7fMISQIUBsyVV9c7JWe8Q+0tc3Qlz8cDYMJY1LLpuIOm4RZKYStYTX7qWk2lBuxCwk0hEWbzZZyR
KpQZmrITfo8zY4iIcyG2XUbONjDSLcM/DCsDKvx/wsdoAJpRI8kcLTa+kzHIDn6E7n+ucHCYyQDA
KMF0kx8P769HQAPox1GzYFRpvchrB+AMoyrEb+5N5rU8OOn2iLQFATmNS+QsrG5Pr1QdIl+F2Nic
tMURAnY5z26E111ieWqCNxjhQ6OsRkanfgGhQdR+xTNlJUbR1Nz49sXoig6IwUHjk1+hE25Ajn2i
w6QPbSILtRIxlfJcIlAULwUeLmnvN/qF3Op5S0zFy8iNWVgtFwotYAabiqh8y6d9wFt2Q1+6fKv9
apFHivD0BkSwgEFcTm5wDjfRcs1StZVncMDUeesis8ezhLdcSzq3U4g4AggHYQS7h2uUzAnQdUfi
vQO3a9LVoY7SJfYQ8WgD2W6Mou4IVSCQEVSy5lH/wJ0ZDF0YjTfpjcUJGiQWQb/iuoyxiQEUJLSG
cUlmvTDs9drjdkT0gZiuONmS9c3UlwniYpw0xZ3lGN5yVAm95NQjpvcJ76PJZrSNTm20LT51xtkP
diV4zLT4Z7ZPKlkllfx66nQ+nSZYQk55H5Cv+AV7ZTdfktpAbp1CL/NaWg2JH1eQ01iAQINx6ojl
A/DggagjGyKQXF9A0lKHBX09wRAsNZn4ELNlnkcfDHcFC0tQasKF3y26HdYbujsjOG6ynMFVHhCl
uMv6IUd6xkZpqI6b5GNQuFFtiF0OCReTEScHs09Oc12A72UrTsVvnrHWdShQSTABiAzBouMUXoNB
aLY+FDrUICC9/fMWtWq64VMzm4Z4CUwnRtT/WfAHzAXo7HGdIuiD0dlrWHjbh6bUAr4oOE8DA/sF
ExGZRHJ3ZYTr/Z0uyE0BWGnk3wMwGeJnUDEpShTNKwSzA9fsWqTQktHAccQuJRI9MgxYJ0GeLmFs
8H1zQO9TvsuJfkIHkpUcdbz3X28s9g2McY3AO0QplHyVyKS24xZLUZkxsvRFYGaXeo0hadgdbx7B
MEGi6oQ+MDII5eNzydp9wtP5nBUCHGA6nAP9THrhZTsR3GNJ8wxSyplPMGyyPKQKyt7ubx96Fen7
WmBaXaJZPes7m0/du2XpfBVonP5BQSqA6bECW+iIy+iC7rFJ9zKMt+aEKmcxP7nvdBe8Q6IAin2x
A+OStka/QUguXj+hO4xZqwwEUZTUu3cs+qTtoTljCdK6XI8OEfg0WTlhtpS74q6TpF1HZ1vKD1l/
y5FCVCyAmq2SBZmOmVz6HNRoJ6/e7FrI5zOR6NRpZwlM/cD/7yfoev8lAhCo0pcIPp8T36HUrc9g
yZfvcVUfuNUWO/r1dL7y0fCzMz7qbH2pS2yIUlkCj6xQtzVfs/6ObOd35UwWa4C22EkQQtg7stT1
vfrjVKM25Fvm99EcOSvc9xChDclv0avXbfpYSDHzSafFC//UYHWSnMIFhE4bbfaovxUyZAZjxnBt
NQvthE4g/jvb5Z0w0HDhbJDf/LbV4+agMKGkXfcL3ct//mSDJVo9JLBLvxPbyWbnwRQpEpJ/lmje
+BauKYRf9D5tcWVo/UMkH/3Z69QgheiGSx7gX4CtrhZ9zYbEG7XGAA4Qf0I6c1bFXHK1+OHLLFPj
Uny+gzsRK8CXW7TQkTR4DNfeWRZoku4RS9zQzlJ5Gsb9OXgCP4UwW7IP5SUaH520vl2YeQ4jlEG8
fJ4MrPqQv9306RVqCsDor01KEPjq7QKbIt9xntlDvg6Cmie1kkciM5Y7Ga1p0ujKWE2mFxZPjAnV
OjbDSt6AzugS54FnQrLMJ0HGpQjDseguL75K8oAiWL0ho/bCPq80UupGY9oqvvydaNHPtaI65QiZ
94zE00vAb84BTbG0EdHgPl2J0mUqw1xC3eiGAQYk0WQheWbDEEKyFHx7lhA2+cls3bchfGQjJ/cV
lmY6m9tsim60Bqzo7KC2gAvRf0xTTcpP59BgeIsfMDs+YBDroidZUkut3jSx8SA/kd+wIbvi+XYS
jdlqFocqDQzCgX08MA+jGb2I8dJY9D7UyRgK+W5Wu83oK0ol1NlA8Dl1emJn6TSv8Bjhr8E2gRvC
kd2AXsa6CAloMFgIv+0rLomRJlzvALDRQa5ezNyAmm2y+YqTKyadmwNdiNIyemmImp64GWVTjRUa
3kHwLT61WUy5v6sRGyXMJgbQPLeBVYJSgonp5vektGGP+DvoTA+ZkoyNGsZBcei6vXzGwG7eNReL
ptcVQlIsFNASs0gf7g64TanmaHzdkOn/tvQjNU9LWcQzRdCiqQtBe6vMwL5690WYBdycdzKc97q3
sapNIG7zUV6JYjHgqAdS5UTzOoOiv0Y4X9iT5N6MMvLKKxQiTTynf3NJ8NsyZgJZ6tsPKjk0EndG
M23po580mEhL3mgJSitDd1qxYrvAkjUzRyvWcnrjhikE+LfSo/vT6YKsN76OTJY/RpwjTZ4EGyC8
+i083iMlAmIkau70InHoi13RD8GLb8u1JxxQJPdsWTJo53OAW507DTxUs+j8G7ofKWZpn+OLw604
kEerlmuAIBEBm5rhspMNXfm4ITZ1OqGFZbmMmFJxbhgZaOLb5u2qVYCjM0hAW3KSztoROMIHF/pY
2TOg31ectOYepvTzu8X2C5XHZyAy8so47NMPcUZV1hyC3qqfIc5OEBgt516K+nzOGrRUAOo9AFZ8
LIl/wgJmJUqjvHuaKw1tZFYSAxD3bRqTgXoT8Eg2opIziqTL9v5aBBddBLe4DRwLV8okNDDOxGKC
+HlOXp6N2ACnmmxgVdZm+rVqPQhjTDuSzwHdPzw8yutqGFZlOuYpAjEuRgejnnTZEWm9gxgm8rsV
eqgbV8YLlaH9wQawgNZRcQdeRl2AJZn/O8CGFfqoiomXxo/CTexWl4aorEKDAa8r4yXvQDP1yzCL
CDfTsWxINVBaoyeWbRDfcTdFywhznW5ICmSmML00flGbCHmjL4zK3k+y6zan1FTJLiams48VmUT2
lDn65K8w2jcK9YnLkDUzyAAaOS3LtVWwXzrdfqPA74pUYr8GUvg5lp5y5j1qPRDLdBZtGw1IgXVN
/eubLWIr6FWCvLglgve0JlJnh9HENOnfu3dLgsBh5/w3w25lJxpGpqD2C6mNqWuCjV8nEjBVhjC3
Es3IEqJ5ogYFz/YGqeoc0QuRm5hMP/uCovkOiUloUY33TqmEyFHjc5pOKX4pFQjJHQD+se6wkkml
7KJeAiI1bBnaXVM9il+KCWELHiROrQI2D7XpyI8m5LX+G6Hz/zEMBfTEd1C8oRkiK700a/KeYf5P
IPBGfIwdgR/+3OPsNptpxDE9AlVNF9iq/1UDTY8ILOZ1rQpAN7V81Licl6VhUPbXStgrYvysoA0h
fnJBNweu2Nfs1fngMb+5Vc3vANPfaEabElQB22RRvbcHNsBKKN+9xPq+l4w1JLbskwg1zbc0Brto
L25N4cJG4l9Fte1LOnxi+CNukyMAosYZAsRElyoLTtFfQ4X1afJODNH5C+IHj5G6luJ5dY7+OMv0
sW5tTC6fH2iQGyy7s6OOfCB9zLAXAKFNP1kMdX1Gn2Tb5EwgRTVy2DGrJS5OAGyeySoOcA4mMa85
kYdk5gGD2qN/xfCEPuw+2/aT0Zek0LHFLr/XV05xnx0leMYsSNrSgJ/+G/UyUgFosX2YbXdNMus3
bVcSmK0IKQS3fU5O1CXVupDqR63xuSptxykvkqLodAUUwp6kX8qg1TvWmnaP+iry0kCw8Ntpa8mh
hiYhPU9jQP6E0AaLCRPoheKd4OzYx7DBCF0xaPzTtY1tusKK0leG4hJVC3knHBMpcbz1qdBgDpOu
fMBz2vvJS/2C9lTzqV0iPyb/u307wZLSur8EbMq0xtxtB5AEX4AV+UkXExSeL44Mw+oApei07DC9
uQb4so+qCM/tkjg245EUjJhKViy65cMX2ZTIT6wA+soZPWV+nbT8mEunldpA27e5pnKoaSR1X8e3
Qz/pWoewzI21f3ZTedA+3sATWeue9njCMJiir3ilG8ShGX1POi5UqsVeLFn/uf1eofLHm+eJUAL8
aOyT9lSGCgrvFL83sVU2n0RamgvT6cswNG2J6t0zFcXFYCgKvQNO7jVmGu7VGFeOn0aQ7n0uLK3n
3fyxK1RAH+2cbe1aisTuTx0WBpAC66nIzSjT/FMPr9gcaycrdCkeX38M5S5dwNUec2FK7BoJizw+
xq+6OND3ky5AsN7Zr/mgNlcoYSJabrLgqLDPLv9SNycN32evEMJRFoIUm5EKtHeBsiPIB7glHXK9
CFi/G7xqnkn6mMg8p0ifUNGgaCQW5QMZxfmr2Tgl3dpVTtZTX2j34De9SK3Zo9ab5UYFXsMh+c1p
xDkyUPZRPsvKKTur+KfQdMaHZfeUgAWj/9ocMNZROwwDEqEMZh26tsZ/5epDO7lpHpuaAhaNIXy8
Nt8Ko2pJxXASlehwVoHjAJ7Dk2I9X05O6NmdLlSEqouI4+wX9V4jSYtXgGq1+TISQ7ImSgTOVwbT
xGR0nF5SSY1ijAong0KYSJPtFix/6mlLYFXLAQkKC0bBN3yqI3SLQ/iOVLGdvuQ/M+ji2jpmb/9X
Dup2JlRM3PuTrbAxJ25EMd9c3niNhkTH2MmDLUELT6gskpO5F/Ve7aV/sr9cSbZpENTSn/WjzmGc
BtO/ZG5IL7IXlMWA57rfiUyS4GhMAUjwd5KjmK2Gj+zcHTT9FGW5yGOBDnmr8fj8oiON1K3QcsS8
z9K1eV1hIwXW7D5RVugZIjWUhf965ToUaxo4n7ziqEQejFL+dRm3tdhX8Ptspv8ggAXAXxJvnnnT
hWMTQTR1zHcNQJ6HdLzm0g/hVsvWbVY3Fmp9dtI1/V3ilZO/ceaWYhkqDEemX9+ac2W2JYEwVvqm
x0tBPuKlv66tqedfPsMLcswfxYBbwlYhHxf1EO1foDSOFhcSsuRS2/kMSyQ+mYGYnrl5yXa79fGf
DM/rY15IXHXOHBrSl2l69DrnJrKG6hdK3AfkIR1goFqMAhIdzTOq9CFw8Y8quakR3+wRYdMOZOmV
CzrRQkAob0tuLx4fp1E56gD7ILFxhWWS3ghmHUDpmDn1jxs5E7dTSi8UcLaXyS6SrQbmMhYAihB9
rhq+ZJ/iuBaxK/TjX0KvhzbkjUL/sCZNvWYR2IDE0Pb2EbrhUDW69EJigQsC9XvPTsYxrAwZ7a1Y
G2ZMZvbvUupniT/pKxD65jmnkkVxtWmnvdk/ZS+5LqPpx5KfFeOQOoYbJWSH2QVM7T25Gi3Egt0B
4rryzwsN0alFlTlY5ZbF5xXE4uKXcPIWDAs/T/PL6Vdg4gi6AzNv5tfWiTFNkqBN6J7sjXK155U8
EJsHm0EPjuTzKW7zPmU4qLnOFPaXA+87znyjwz43mJZ/JSGi9qXJcvsjKLAain9yIJB3VsEKerWf
UqEsgLUF43VAc+uPL+PPMpvdifvD7eTPlA7KHZPm6xROYloOgq6irsQpsrrCRDIH/DwfIOdqb+Ma
m4e1XOnUSYL31Gj94eUQlqFpJ4aDabYOi3qcnVHYpK3pkI6yh8mr6m+ctsOdOb813Y9VaXhQvidD
VAHHmM3EjnN26vjBHGXQzl+JQfasYUdT2o221YfPZNWMCGbGs1vVnzOl958m+j0mAgjeolxgozEO
YOdtehCu1XiVnefWHwcP7akPxSA7wCXnU/cQbVUuJ8gavYmYaCTtvf4yeDsQMIZVe/19WQ4UCzEJ
weHEzemVGxPPor6HdR41s2C6HINfF0wVW060P/vOBO28Xsgbnb5pyqeoF/HFXMEELG8edOGBZTly
tHuK2UJaP/pOcw/xD8bZBAV2V+6o5CSI5mm9BbDo0lvYuv7o67nnGG+tB4Lv2L2WAKqyqH9VX7ta
z36efA/ASrdViuk6TdWnkDIk2Oyd5qr2MLvp7OyLKiD3CechXBCN8X4D8byMBohAzRFtTppu0ht/
LsTZuTvBei9/p0nm2ab1PYqfo8k7RNqPkZQJPtC5ZemKCt/pl62+AUF0dtJn2TaGkG99p514m4Mw
aHknSMHh5ET7b+dv0OdJhy8Px3gPtuegvtEL6hk1n/QACVJgFjaRarcm8nYJtGmr1xulDEzDiDQ8
0rvyvQkFSaeJMGom7kxXnkFV2PNi/PPwVf5PMzo3+Pr7gpJrZMlbBX95jntTtL36Q9e+BwOskN54
AgNpzMfDtgjlBpLHtdW79Z91jfjGJBgWxUbtXchwUIf2VC9FId5mpg3Ccact8Fr+/5qV+zU/LTN2
6ZfbZ5iz58zpUDvTpWaruzJLyaQYtGkKqUIKCsdZYW7OWPQ+hzfCIranwn58UKoR4h0i6OgHPhp5
veRIRRTyCCJClVGO64X89eQivezq/VztzObrCvSY5q5ccddE3ezkvaBehEXze9z0zKNs4RelZnsl
xsJJ6FkDD84wk7iUDQ69nkA0LL8CvEINipfRv3hphd1E7x4OUyktiGgy/NzIP62OQ8LBMmjy6x7D
W1mnsc4fDVCAb9bReGGsvD1OxTPE72+4nQX2Oa+al6SB2y0vHPKU5YZlUTjCHwRiIyK5Ck73/C6G
ZLlRZdEkb/K6SVIsqS7EOcgtmcqDr/gvRpEJ1wiZLjkFCLY5zodSlSbbXHPUf5mgTtFkR9EJ+Rwb
UarzVmwZwu4VNWSCdNQM/f6pA1hZ3sk/VwQvL1xZ28agcU8Kqc7KrI1wUHJuhBRRxFNLeDIowbcb
onQMjULtI3VgD3XWbRIyy285an0jNizB22ucunWUglU5A9MDCGoI6lbDLi404H958g53OjTKPDmQ
NpcJgmz4uSXxQ7g1LD8p5qzn/OeMdUP7yoJS1EvtUy14pYldMKsOSVQAqdLkC62w3dgX9kdUhF2W
kSyVnw9fp4vT/PqD4JgXNuMDVrTrTC7nIEeKT4NDLi9CrB5zDrU3FoTzeVDekcQrWU74jVbdFcHc
oJV1Gcrk/+GneHonW7cJgwmHnM1CrMEzaIYtKPAdJH3LnLjWhxgsUURSDi3UmLP1Fm3asNZo+0GS
+e9bj3B+aBKPgqNMCkVqyYSmQpBh031qLGXaNsYc6zUDhq9liQt1YUKXv3HoouqHUtVjS96F8fiy
S6VSUClKctOiCTlhqaeDj28McZtbI5eqP7JghHBf2xmIP70sL2LH/bJqlqhjqi1SGaG+TkAHkGqd
wmVAwYFZsxtC4FSnvUoEegOTsJIkkDq0nbXabdlIl0Vr+WxH9yVXx7EMVp7Mec10LtIJ1CpSy6/a
XhZ9K+O9vYnnj/BS12pVIVdo9nwW8RIqRHoPDC3lf4py7R9XYmKNMpNiUsCeIJU/q9Gma/gUtCcw
GAQd/UazUsoJByUo1P5KLbJgyXVTKFOiyLvHumvf0gpdVFC3gVk3FRq0HvnEp/u37TFWZk8bjWt/
RlQmZhdY/h0aDudovz+f/bYq+PEzet0HUksPEGmpxXp8o8Jqftj/NZn8QnDV/hd/tF0oXwMAmMoG
GJr1x9HxFMdVKPGA1G855TaqYSiVLGlUwgsxyQ9Fz7rel+pSyJxWO3FweU7JaYMAGJ1c9HC8keea
vnvlBvfaXazqMwsihO++HDHgdfDkuTbIPPG4wzLdi+SCTRn5t5uSw9SXCdwmNQkVwmKO8GtrARqF
0IVWT+L3xaf15NRe6s+FOZyJiBSVkw0ksBTGapubx/HJZJxg4uHKSI+7LhxfcMIlMPWN+TIkvAq8
YzItFYw7AX86gt/ygzJ8xF0LQ2V/CQ/Gownt9UMkzs9bNTP/KLGcY+usp6HV/7SHDM7E6NWUVwMo
qdh039xdlEGyg4yUz795xKNCTxdZ9FbpY45A7gyCnZlavqGWNKAupIrsBtToMXBPQ3sUk9gNPqvq
3W+wjMiQncw0DFviCG3W1Skr6NYxZ41h92/YzTx4UJLoScYIvxpZ/AppLEukxrcWPv3QaT2KFlmu
0NTp2taloyVBO6vdM0jSW28Juc3ZXOaNwtA5DUGqxA2imAiVS5aGXdJ9G8d0r7u/T455UDL3HBrr
q83nxqh8aqE0Svv4QFFPEAI1YqfO/Ymv+FgB9yORlU5cmKIPV+1nuwt/C9/drc2tl5qtLgQilZ2N
KV298rI77f1PfTS0h8POHOkloNSZB/OkK0LoCCFxrTqYvCZNm1LmHoCF/XrSYWB+IaniYT956PPa
CF/oTSWxEWNcA69GUzF+ZHAoDP1SMZk5gZmvn/HEAPWM9kM8h8EMgRCY1GPvn0a8HVG4hvIiRU8Q
0jR7dyVidE9b9idULBIGTI68q5FtlNjR+vH5ghwRnjx0KQhvHQCG/QLCuuJD3rUsRvvqpgmISs9W
Iz8325ioX85tjmKKAW56QyJiW0N6Y1BI6TcIsst9yYQnkkgI8SK3tX06SB1l3KiESbLeBpz3N7dy
a9EsTzQcOHJfapu0rPD1mMq0dZOxRzNm5LS9TDeGiehs6Lkix+DA4rMc0FOVxni2LHJ5dcGJxWnX
aP4kt4TolSMtkZF5nFjAevMLxbY5Gm+x7tFR0mDlHd6IycizIfGYtE1AjSkfHhVCUUGLiZ89viQp
2/1Q1GGkRajSuld27HL6eI60Ar/ZdIwulYKjxeAOQvh/uVTXI2w11KWi2W2qRgUVoKxTAwoFAgZY
SU1fok+h7HM2xUf1DZgzWNFn2PUWsqcSAFP+dvLIVJNPSRw68WZlDTzCcovoKgOysxLO6R48BXIJ
l58ZFgqLfuHAfu6NdL+rFu45Us0Os+oyxI6GquX9ZI45e1tnf8fiCG+QcwdWww2wWX0sb/dYYeuh
iaG8YGqciI9B442XfJVBoJ7VYks4aebeG3bkoXKwMBX4Jq1KQcfdUt5II2R9h0Kl9YM0XfCLQA31
FE1Q783qmFF8P/0lFFe9kyhQtDWpipFjjWnGsL91HhZyBHc1R3OpBwoS+gEvire8NSed3lO0NNI3
pmzbyGD/qVek4izYjAIR0nBCFWoRAwaiA8gEF+V4X3YD3YQRZ/JGDmRDw62mtXwzAHI5sE0Ileyy
zo3JzgLImgOPtQZq3xyxk12l4nNeTSE1YcLatNjqy+K88eM+CvnHIsrriMQDbdmlbetXz9rtr2Xt
qm0XK4ssq2nuPkxpl/YiYVQiFFy/CUNSsnOzIS6mZnRghG029DNZ8GZR7rnQIzlC9ZASZoBacvx4
EQzRXhEYUxVw9p/2HztSDLz9k6W+DYSt05FzyqAexzszglzj+UUG6nc1+nDBf4jqTSS9eDnwI+3E
4jUXuY67Bqt3dhtKc1qlvKFstlSjB2jsgIfARWlYCse5NNeK4IU9vANCgnB1r06CH4hDd78bfIAA
xS2dVXX2hhEYW/kxXI0WbjXKlSoR6ziRon9dlYxjlQkVnmHE1vwqAtqSkX3Px794zd/K7ar1xH8a
cXEIEnAautjIBRrZU9fDQQ030wggFiPBzVF60bdSuCJDA6hJ1lQSm+xkddpq86CiQrlBJ3A4kPh4
RSPG7wSv1gx0ZJmjQ3ozGXnEYXCDFO/PKS2Bmz0fvEmtyCKJFQTlwHMikOdv6PJV0rgS4OVkVzUm
JeD+leZVEfvOMObZAcmXhaHJOFZpIImCC682cI4F9hT/u/pGEyHgrjbLHUAPNAmTABsCoQga1vj3
/CGw7RESEwEofCDxQRR4BLdOCXowZBJDBtJG+cXL1Dx4b1nso5stEKr4v2hh53RimGgfSaXwnreG
tkdU6K4kintUiXjQ4HdJHQo6RGjepWHZc3qkNTcgWVtUZ861ezzk2TRCx2gXKQclIu8LkpinQETD
3FLyoDlV9FuEKosTXOMGTGhlaweqnNmiOiRxogWLq8Eq8PZuT8soGO7Fl1jMfknmeTBRYIrc+egg
Se2YwdLPIFOxDwtpJpTVbUYPleyJ5hYllhgrftPSYOXOvuiRlrPVpmU4BppD5odn2zNUEsZelFlB
yuTHJcOaX4Min1lYiIY5QBOvIWM0OiugbGH4WKKpdIMYL/GCCbMjMN3QbZCoL+hZKRmXMuwK9DpL
G8b0eR/y4T+lEVuL4OwCSSIawUW0lryhgJm1iHHVYZlgM5ARgy0YiPHplU0P6MAsOgFCr/fiGk7K
vjLZ6jZocO1gORRSnDev28c9g+7bOsLGPMPM7K5+U/lVYHpliVOMEkUPnXbPFjL8teHNtB8Q2bX7
gSJ4wYyImTTuL3e7KRHbV2VRQLYaHhbLpPUSpDNxXXPUSiNzhsVjwLjUeEI8N99RCELkCs1Cee/I
EIN7IbkLy3ZxkPF06DF9qe7C11VFtWi4P5ET2R6Y0pXphgy4AW+j9m6eekmkff1xCX2iJJ5f370l
NTaUbjBzhOitujn9i4oPFZIA+tYte/0le/Iop1WlPnP36LYPOTlxZ6qznVaDw3wxVjrP54UeuvYm
lAdvpAbIj/AqMhf6fQms8HN0a1OuKUrz9QGd/YK4XbxBvhsnEFwOVaesz/gNspYuXCUzM5JWogxR
xi8jtnZrhQveVxGZEliT82uiFmPb4pazebqFWUyIRZr7bPCfTi1OJcHqbDWmjKNFIT+eeNSSycYc
TNd2TvkLZNwApb7XVKHPfKu4rWrwzHENnHx6DFiPuvVg/AiRgEzIaDHcFw9grI6E63X0oWpmtLST
GY9xN/xv4vz5Hozs2UKU5XtJ93zyUCLosCE/C/nCWemI2/YYWl8Z5t4/admyRerkAYV8zr6l0ipQ
219l3+fwSpof41UF/68+yyJ7Q4/wFUdS+n6GDa5snjaS8oV+xrYE9wOQNu4F2IwO4dfoMg7FfIOS
QbF8wdHYmFlobyhdRtyQr3AFU+JTpz6FaiS/ZHJnbQIqPSe3j9hfnClfS5frref56tvI5GXbiKyY
Jqh5zRcs/7mESxMzQkMvf85tvEtOmi0Y8bt0sl+sTpk+6NxlBAsS7dX1BSBpqnGhuRPfwXpmlQx5
VQKwFmiIOHRGWeF6oUW/F6uG+NgcINQ1Gb2HtlvxBUsXHH45YWLGzYZiwg00lzbN31E3qvpQgB2+
8RWm9r+pblUpzgdSvf8LmkqcF2taBvU0GnFdkkgspgLBMQrI3x8EWtHFsnW0LXabECrA6knE3hkL
bw/x/aXP0TggOt2p19BrUSklxBKLAfaeMa8CbFUF6ELHLWpmK4g/4qgDznA4XwvWYhxEHGL93lZ4
OJ95pBgVUxtJsXrm1/Oj5ryOMmA3xrxQl++hgK+Ks7x71xmqg1cmapD6cxcfXbbSNWEF9PEHCIj0
4LIv1YXvkA/N4UT/KIHudUQkqd0RqjAzCGa9h9EOWelrJPqR3RWQ7KkElslp0hSgBcDKadSKnHGy
ifVmKzTHVCSJOBAAAtCn2UeZqb+CuUqSRNKwU2AY60j9X6AWEnfacp1XYbjfAalski8OERXOR7uB
oaVFryhmHOheL9WOG45lB7ozUduQD4tqZv9yzp3Lw92M9Tze04faVxlL7qwNpVDXcTybuMCI2wq4
GOlXbYllY8ki/Z/etx96tnRjx6+EG1tpdDL3+aR0v6u78nrju62PdiaisSaFVdW9xTPKLNd9RH9y
Z1LKIq0jhw4P5vJZIh2lBjRX64lRIJy6ISKAQlcfiQ7w9AVUSmwcFSPht2UPtphL6wYsO04lcZSp
iHXCQuzAXpzmAbSp25BXp6ng5CIbAb0Tlvcj4l6JwoMvSzUeT09BH4uo9U0Z0PuFEN+lHwAnFZmj
NAugPadgDjj7jNGIQP0jFaH7TEj90O8CHLp+gGbT7ANGmkUuBdj2PWpnPLRE9KYCvFO1SnT1FUs5
s+3UMn2IuXR7ciKI2tw+ah4/35jPebHI31VqwKP9WuHGq/Iq5GKGqITVIgTmJgR64jYCjDKmCXFp
UEi5wMyAQeeFLpve+w784N9NNZJVSVUCesjV0FOOZxTjn3Tm/RLWsMJo+VH4x6K72xJ+I43y66ve
0cONhLVcd57e+Ld4uewdaYOWDD1Q/UJ0vFYi0ARU/SbLpqR1dKQumlRNhCAzG1S2karhu5v0L3VW
n3rbD9gTDTvQcpHxOOB4zNKNugQH7TSiqmOBGgFh/RTcIlV0KFapuq+rCU1n4kUsElwgquAOX2ru
GXfouLd7+radYGJyADQ8ZfOUzL9TfwGS1QFMllo1KWDVYwKPApKE/In482JIitSzuLrm2JU5j4V7
J0305OQeq3wGi26Dbo8JmJWlQZFQa28AFSyC89h/Jo0GfPrSeJiZIMRE8/gTOhF+dbpWNq87T6VE
/v8InOl8ovnuf59YMGsLKhQlFATa90CdDpejmzKovTZ/4foDn230R4/CIwRKiH9O6qJREswMo6Hn
3L1nvRW/tWX/+E6QcS7QcRdoBEi5dyzEry4GpOvoJG4s2lwEmBxExGT4l2eI7z/WxfYHWpLqEAAf
RTpL7MJWb5d2nkjYm5muFQ8smcGuMDnOtMdkaNJ2fgvzEZNbZZG5nHGgvLeitvroH7f4A9hejxEM
aiheTD+dsmzMmILPjPloD1ZCAsUK4hLqfffGZPMjslTehfWDxOU7Iz4KlclLrjczEX2kUGbCLx7L
JB5RZXN8ME7BfWggs3E79KzrX8AO9QD4DLKkx3UKyp1DcKn69+ZDa8cFlRieog+CsrVEpaStCoWf
uMZbX/wP87AgF/4kRjxXarbAG2acFT5xIPxIQoFrDlp4LXNLoPwbe+1xlnN4ljFARCmGi2EvVv8C
cOYHoSECgYE9J3yrqrVw6Cxr/7m6hRkBA3fLHemhM5Vf51p8hT5GFZ5j2cSvLD0w1M9GPJmHeFTY
PU5Kc9tAGqsznEpBK5qYjbBBTLl/0NHlk3lKbGbjfcqKgqR7FC423G+JHF6Tu0tAWRbngiYuy6dg
niXywPgX4aNgoTJm/DMqk/QwFZmakTENrB7QhAqxq/KNgHdUdrrSMj6JZt4cMib95Fs+U+vlBxzn
BKYXlhebyYn+Fh+4leUTXC7IaaMw6s2VeokaW8BUCQZpQyKiXInVO9wxRkfg+rxpZxfFqJTWn30i
XiYKwjGcmJau9sYY6Y4EgbDMPjrt36FQM0QCT0QdFbTOyUst27KTzTubiPClI0Yv5Eg3iRR+Onjc
oFcjLQJ4XCpGmsAulLVJl/JYqfPQ56Uczj7CBWI35Xc4GX8QLqFwCBhu7R913Kewe+kI/N9hslMS
3M5Sn6OC6Axz33uHoZACTkQ/uGIUg8CvZIhDWKxuYPNm6UYB2j7+Hrxq3M1ogIq7Q+ol3hNXfLif
7Bmn+ZYqZebn9a5QoUSbiUDGklrVlOUDGPz3Z3/HV5Y1482xN6hnN8G93fQ1eUnKMkK2Z/n4dloU
l3yI/yBRbkUE7V7qBQhCrdBWRr64BjQleRNr0tmdeL316YUiVDESalbqeEEEMdM4esGZBNl9sr/p
7xEsGzMWHivqZjQeVixqGxVF1VIHn5X9no+yNqkZRw0Wlckp3NUUxV8+No++rmt3tFTcqadHWpTQ
VuJj0vyX7vrfWyPoSjapyB0TkcvC0hzPcOae05CRt4QEcwpDqhjhikO8vCdyfWwHE/FaszKqY9iu
BcSHNOqKn6NGK20l0feyQnADNxN7B7r5Zb61IRTXuYMnUy2v+UsoWgo1u3s5KkMXwwOvieTLSbi6
hvyku/BSXlMUhndewEKgLANzE3Fjd37qaiY05GtyuWK7UaiSB76qK1uyRBSw49b6udNBDjSZQPUg
3MIeO+WoCw+umV0UNUYlNlI5dcmG3UG/8MNpYzFEzbXRspYA3QrPFuOB90fA7o8659/pfmNEQKox
ZsibSx6lzCyvsZTaAIzCEz13tf7qBxumGV2rGI0SgT94h4U1EraWqojgs3hSoqONm89Rli2RpkWo
Jk+U8CBcvum8Sz8ya6xKRbdwjqj1v1pzux0OVCQ1yUas64pNGTqaI+R4yKjljR4y2DRNTaF54sKk
jhl7VWwTtcRe3DqNu5JOCCLzAv7isNa4adZub0sQ3AkfciV4T4e4yfIYqfs21QXNLieOSw3C/sHc
joCr1YRpW6nHJF4teeHCQQoJSa/B85po68wKB9mizVCjCTBEbaRLX0fNEVEbD1AcgA5kVktxLOs8
Sp5hpGL8of5pwq4BKs3mcvjNrT29P/aM0uwQlANAPS+XgdR8IwAQ79s6ZaV0bsdSzIkpgMFjrcly
n8MtyP1TbYC2QhVCwzRxVyBGKKtnume4zrd5miNqOzrL8Q89hNiwHY4tK+XtBBKSsVARz6X2ufLW
Cs4L1+DjF61JVdrXIhZvqu2L/yiyZLa3zMv9bGogNC9sogC5BCxUHSSdFM2exGhXk7tBYvK81T8m
mRQkPPbzjGudG/2pnXwNtuv3Ep7EHQHvHeEvAls+l6os6bJwgLtoaU6H3OGMyjW2Mxu8HFFxgiF7
koI4+4cE4oqUVxonyXM2mSfc0i/Y/nxZgx9p1UTi0xDUVeVSH7CsjBzR0xsM9+0DElfcGPgZBJDZ
ZFVCaDoPqc9pDMT/ZMaZ6PqM8WE3YrDHOJxb1+iKKqiCpmG7TqLXnpOTzLEdrTPxbEtiJSeiWhR1
wSzuaJWCyDJU9ghlz/LtgflbI+GrqJKOoBojhwPktPZM0+bIa6PfIm49DtrePL4HjN30niF++9hA
K++UKjv7JgccY1ISacp23BSCJSs91hJjQOb/rc6GO4C7KIfsCKQTYsS8TufUo5AWrXHqaR5oIkac
5gYsAFixPhXDS/MAXZXLhvmZsGonbei6M3EwxThyyt7TG1SXOBWVNuWQdK+XSgOxFMs4gI6Tm1aV
EmQTtm1AlTraE9NVxecXK8eCkoLl3C/WF66NtLm9OVvwHV0q9zLuZN/krfsClrCoAiPZg3v7MtUC
xdT1uM+i6daejLTRp9+nhPODFRMh9ecrmYT986W4YA8TrC1aPobyqa/080iKlnrQ5rm9Fu49BanZ
fengyhq/DOv8s+t6XVsgtmKdkff9ea/60P+lmGEEZ/h72dGaUQBArlIpzFxDDe3O6WABy6tEM1ae
szB7mOo9a/p6lPINrEpxDjaYcBfaMo1lUi88VUZcYifqp5K3kjRrHjmeDhqroQkHEqxrEX1gytK/
dy5VjE+CGxRi1yACo+aKvM2XJlX1r5pAFq3tF+GmxAFuSmOL2SMme6K6D3/46t9l+Ud2pehS0Ojp
JvszRwFEX1UpYiGB08eNbIDOiHRYPgeRNoCukvt8klP2FY5c/X3KKbT/kLfW2E1Sw4jit3dbSooe
KfYtdCYu9mtl9KQzfC87fbKfG4nECCzimjOcFSbUyPH9DjuxwZN65IPcZRk3RtGCFehKx0b4Njl5
EJW3dQ4sZsIeR6oF48zboGf1bgksq2Rg/d6O9LIuVZDP8fWAIzrOI4t0QAwEYiDrn2gnFrLVIcr8
feMI53nUGujzc6A/2lyE4ysqP214fvP1iQB5itqluRv0KzizlJseTwsUm59LGtlI/8xbSucrtD2R
Vo8mvqdTTHE65ir54vrRiDq+LsfX0lRg6LAmB/C1DkD5359225BiLzN18/6gMsbJmLSYiApDbI96
QJrxgBX4vmgHWprk/8o3eflY8SJqoFows8KhRDSLr50VaWzBJEADRSvwkygMwA6vLSMhFtLttBy7
h9ScxPNNw5XNOygVLAgNMPywkUYj/SsCZvorfRjCWab1zRvR1ltFcUGQP2PTPdDzgrkyE9MVJ5b0
Pb3hRQsmwbqfoUe3s/flMwwH080g1/KjK7aO6rgdNJyUCsUKA03M5dIN0TWqolQ5U9/xbfsV2D4+
+BhI6whz5hpsCJI7+ZJsZpYdPrmfH+WRVgObjlVGJ3Epk5sFnvr9Ip9k3opBrMU6rHKaTExhAIPR
ikpXzz5OvNQctXqpgWL7eyqjTGsypeXKYEMoVY3b1oAs85OZZzzaK4KYYvHMdBlo+zVbWrB6sH2k
6Y4quS0dl7s5V1eteIcYxvV7IvKlSRrejxGe09xvjQ2i6BxmsaF1730hWTb4lL5LNXHeMZ5eLkcs
XM84Ro4jaKRBZqha0xXN7OPMvR5Js/BZBT6l1URpUulw52uc4nNUeEcDc3/VT08oPPXxuERH2s1E
Oha394siCnxTTXQJVMNxuZs3zAp/eluhP1iZCHtDww4EvmgR0MUOnSwFVePtnQztjSdnzlgoAbTQ
3y91D9Bxlb9X93GOoa4Yb9n+13C2OCEhnTrvAiekGaVF4NNfu6I0+EnELldeRyuYV0AdcZhDFQpY
cM3O0wWNJ+5gWWMs58U8tOGVod9xKbr/oCR2Fz1qzVZm+lYl08zzbUziXIE9jkThLgimsztonzrl
yojYWDJexyyTswid1b9ENLEI26jLpu2yxRnVBXJc7HRsEQK+mCHggwnhvFnjSpe5zFXnWvL57Pa9
/HvHuRUhth7s0D9OhCMc381cLoIY3kep2SeB5edCKcnpABHxRQzoeA9xGZgVXdZqog69vlBv3OMK
eydsYbJnICoOvyxtHQp9i+w/K46Ju3GPm5s/YDjwlSH0GjMgGhWyA681VgmTYV/ZQTsTKR6RXr+2
As5zlAGuY1JhdzAxWKV/UtQivYZ2dLsViiAJCw5uWgW3g0ZeZ7B1rc4PJHGpESPq8Y3pr5B+3mJH
bVtiyRJHil6gSYRdH5GWGFLmnE904fecvsxRTxfYVvI9EQzrqE3PHDruA4cu8sfrZjVJzx9uixjj
kiC7ZhFzf5yTQ0KUoLEhIvmKXwJ9TRmCzqGbBmBvzmkZ7i9Jf37uSnUuL+fPWIcNbyj01fmIPNbJ
YCdonuceX0FE0x6fF/8TAVwO53k1UpvSuv2+eeKZc1ppzcp0z6fFP64RtN0//XiLW86/pG4XN5lD
pJU6fBBIT8mr7iIBVQ5FmxaZD6qi83WJ23FfrtqunrvNYrQ9UdJL5sGL+ACMpFyIz5ZCnzEvZM01
ncB7VuZvpv49LE4L7rqWxd8v7KdoKFsiMnOpiWz7+eAiXSUNj3adX7ifTMN1FfGy03vTMv+dyASr
FxvMXo65EeWX0Zp4/9e77ITjcIZQkZ88TiBsHv+JWZgQzr8FupW9wvvNzG5Hes9lS4EPNOrFbgh8
rHD1wrUbfeGTHNwKcRmW9ylwN00PnkzqlJ639HbWDSouo1In7gf7q4f97oQeeSrQlwLsH42fCtfN
Pf5qHH7eX66sDRA2XDKLvealohXUvJTuxmeWLlAo23e4DmRYTck86n7bi5+IdzaZwh/NXx29ddaC
/gxyKGMKP7gU+xXwtiXoP4jAGJcvEWgLM05aOVz4vHOLqYbfFak7/YaE5dtLN1BNoagQGOhklh1o
yoSrwrLo2up9bsgFYmACqel5z2xkgIs4jmIAzkEmC33sLHw3j+N1jk3WiZD0pDq2VdA1GYJH6BVk
Mn0Gk6pnL/nO9Tu7bwSZM+iGvI0JGflghGwxF7BTwLciabaUg/4m8G7edCfUuwKdDGUsO9kokm1u
sotzB8iazyzZjwz0ZdpQsehPRbBj44FB8ieKvi2VC9rLn683BnI+Ej1cWEkuJ5RuyrphqbzXSZZv
VFRejha/P0lwVp0zOhLGKE3mZHUuyIpZ+ObLstRg6nGhSVydycYPsIx3yMd8vwr2H24Vek8673zi
Gvt0Te7Ah+AkqiHfkezz2c7gFjbhg+KLSLcwAP2mQUrBOje8mop/HA11WSPIusqsDlfdOM8+jEdZ
S78GWYInKGg0UaZ3ySSzeCyav81A4k9vl13ThSYVAXcLx0xXYYHGuCUFgxiYxvP0PF5IEWDqCwoh
uvievJkyLcVKMbMzfeBDOVAOiAVs/CRYmzAMNnwoQODEGo6JZ9WNURTfq25WxirWl1OqONoGqL0u
eHoGdSNZSNpCE7aan6xErdTDf4blvb5gcOCQ+YZjSoVOkTrY9Cecsr3T2cztXD5fGqCnfEm1JtJE
aaiBer4kyA+DwuNLGYqZFCOVzQ2rCyJXKhlxP8BulDxgjdWl/GNNx0sIax10EA/5rDOL5RlKzAow
iDkyBWODjlUMYYqTD48rsp571c5thRlz2Kc8Qkfnc69PDBnwjaC5ADdD8rol7bMpiaSWu+mtiYJN
SkriYu1a5Lt1BkFHh3/o27ozfDXhvb+tWYGQKm1p5zxouMpb829zru1FuTqkUJFtQvc+0VnKVelY
IoUeKJpGYRYo72TySGSwcNc3gGcy8GP8YTPiTZzZT2x6dL7IIO/3ZHH6NvpOJ+KfcdmvpdNrh3Pz
9nqueWnuWBuEwA/LhLLc1TEoqwggaHUQpq9agntyTH9wDJ8x3wHZvVq3EkcQCp7n8FHxfOZwrmsN
7jQNN6+V9YB0WQuTnCrPSvF+woS72LLbpL5XgeCFzXtxK1fGrWi2LsLhc/PciOerW2156tC/Pubt
nE9OD2RVjMnjrBhDjnaST0LC359PykeedacZgJ4ZRIjVfd/VWu2RbOwHF3YbZzDpUBeFjJGbpa0r
PYmR/Js0Sw1yM2ciaLSeX7Q127rxAFzmK0gnWTUU/Nz6HT2fqrnuUuxDQpFBSSl8+kyrBjjJMhOT
K9DGv9UgX0+zSpkalNPqAADeCeG9mces8TgH9jRtmN2AVXoDjo7D5cE6ewXruFmFToTnSE8rmG6c
OacpZ90z5nBwFCbvJcshf45qOxRZI/CGxa2HRzETgj3wkg2FtuJPF7l3wJ91SW5o1Hh+C8Zct0tI
KtoXUm6yEHDUwnY+If+X9LwpCaFKpZM7TAJSsWexu7elWLZ93wtubxvRN8OAeoncywf2Y53NdMeq
R9nKsuChWeH0HBRcETBAa88FKv78gfhEFDk/rqIQ62iBFVTpWsOmwCvtldRhQNZjNsFXx1Dmgl5s
aMkJ7sa3TzfkZHMJWdwaL6bcff0UeU8sfNImuHqRUbLl421YG0DwZGzx3ZEjQo2vmuUivKJP7vXT
v0SJ+3JEFiJ5EwTszA2LNnaLOmusAmy27lCS5qwP7t3bWp8O4/8LmwbhIq9nYKRXiKpMJQKbDOKM
ZkCdNqCjEqCCwsfjauUpHDlDxqg5Psm+/IsAvup7hLMJsUHyrt+U/70pWBZZ32mRoUXc93gGPWTz
azCBqlrqTCrYes4XNfK/gkaW8t698KlwizAGIJN7gzK8/hl3sHLPtHz/xlo5jCSqOZys2wkqJ0HV
f7vrzyV4JqFrsZjIKHTgWJQ19W+mEdvsnTLkfs4G4IFmv57xTKIPOeb+Q1dKyrbd8YgLpdNkO/v7
8DittQa98i2m58tphyMofCcLLMnuujQ/FqilbJtPdQxyvOOJemQHjYVv7Y0acsWmypkAKi4Br0QJ
pQelUCqF41ej1nooLJAvAiCp3WtVe1fJJoMLZSXKLWuPn/gMh320CQgc+DB4Dy32uAa3tlkQlJaL
jOFlVFNlu0M4FZO43oUQzpz8k+6nNltda6QGhmRHocF1WI6zYPm5Yb7ESDo5IORLiP4sAtZ62N9y
7aqPymWpuBofHMyMss9Z/dXMM/w+w4HcH9N1rK9WfNk/tdekKBXrBWOZ6bVQipAhB7SfdMFIJWFG
EU7Vj5n5uXUWyljHMVE6WmqQ206PIrE5z41zOCtl9uTeoVMo1X9tZWjA/ocK1OnGgMHI58tMido7
qRWJ+j6ASUqcfnYG0BSu71xgUx8ux9QMdZoQzmTsGHKIbrUCvoBGFfXVzj5eSXsJ7w/aQjBeX77l
G3y57iuE39UxY2reX//HhRj42EIvWddkTaR+pd5MTt52HVkJA07GaAbc3YfFGyX4NvK8mN3TQnFP
xEIBQgJQBP8dHcEEGI1FYurb60h1WeZsj4OxrCFR0trf7BlSy89vwbKpFuufEVrweiHM4ZaZSvuh
24wblgHzgH6gKAhmkEXhLFJOFCBSw9UadPolkPnl6IborhfVzjPoW/xitDTJ2JZ8B+UrqnEGqcOy
3eIQ4WW9YVxnKgkQQ1fsCq9SR0FK2PRufaf8rQRiNoBiovK/H4u0+I7oNChGajWT4H3kB+ZTf57H
5H6NSOa7EmI7GiUggodMGVgYBM41H1S9KnAfislFP3VvNj7HbWJLkWAod5Xh7CChaVzmejjVkTio
z8OKqHSpBSBS14vRDC8nuFE4j5yxqbyYRJvLEppJ5XoVVLa6+BxqRNzPJfO1FIpcyREiHw/PS+/s
itgk+wYcLZnouDSJOifMA3o9ec3Ay8kRUs3uuyAXeP+YIEeN71zN6I8sEwUS8ibYS+8JvBmz2M2i
fHjRc8myJnhuGKuf8iSlSMFEZC7K1FHQpA6SSakjMvbqUr2LqhumTjHEuTsWC6x/N9DoGg7erLiS
S2wtHawGAcMb5obI8iCyuFBMJV84mV3bJYV1GmeLDcYRgRoTds8ScJVOXY4d5p40OH5MYbMJw788
hC0+3Kc1pU8xUfmqawGEmvQBnrAH6tatO97RXqlAQx0B12QuB79WfUu98He56c6IlmdDiFA8nYEd
w13/93aBa1kQRDZot53l0jkQEhfYKBjoT9iBGYBB2dSCTcVPEj8I9kIo4DDXvtnNeMLgESWQVBYA
ad550K7WB4zMGLmxeBuh0M0Zo3KdSEhEoKb90BgUVQtUm4axHnT8ZxrrQx451eoIjbPUVeS3R+a9
rvyXQLbVrAdNY/IKdUBZQUkxzsnFVMotjAlNSLan62HYd8fOq40HosyAyAyvlkRgPJ1MVTduHqi0
FOQ/+StcwYDkzoSQlcqfsYEIIe5k6XSbisy//Tds9kVRm+0Or5uaAHsmffEg+SCYnIdeOI0yh7s4
7s61nkvo5Top79iO8DTGa797OPwboMcQKcaeEMqrONPqcpxr6sKNbwUlp8v0S1brSNrqWdt2ZJpE
Y+MGAaye4DFPI6VRfKMJu6hWjn9mqC5mYVm416Syx//hEJ/egE6HCTtMBZd2DhURSJJD2kdBh5N6
PT61/UecLAYptjN4wLZsr6dIQa3BuMVCYQf/1FVo9J1FpKlQLfZg7jTqA0x05bEVsyfWIs66Zkch
aSIn48++lekQcy1XtA2zVjUvsfO+NVVuB8pmlMnWzU2pKyP4oWd7pFqyQL2VOIUtJqaPXJe8IHPd
tbEr/e293Bt9v1MZ/IR7GY1ARlbLGY/udmM8CvufcFKp9zant4hPRG/UzS1EtwIyIgPIgtNW7PU7
nfZxaaOlZbQ2XouP5mqx5f8Vvuj8PXpOuWqFcqP/LXKKD+FM0x4QRXcOGRaHLtzdmf8lSZ0Y/5Db
7TRDrPThBSVnPRXiYOzv+r+vKWA69beXYe4eQaNyV2OT2rSndA1DX7D5cM/o7Ca9lpmb66O6ohEW
NxGVg07sK9QMtaAEFaZ/cy9gpPopR201wezMCO4c0WBnr64VOQMAyIxLv2Sc8HndAQ579XXfd5ru
ETfqp2wN642SyRXIya4z8/TSF+HyozrEdmRn2pmaydvWNh3k4Dt5zHTJBRf0w9aRl8PWVPfEBp6d
s4ePSWElC+Ynj298Sw07SKS+NwR+ApG3vmwNdSrXDw0L0+X/+1OWpNFxjX40Kf9sqz+0ar8jo73x
mXlzryLZQkO5OXd516xrOGHhh0AIkhO6bezGGjeS7dd99Y3CK76ByzXcPz+OZk9a9XzWTF8eldEW
madRPcOJBK819K/lC1JT2visjqKnR3iX/33Z2l7XhJl+9TL8nUFAz4dP1JzTgGJ/4h/hcXME4VZ8
9+CBqKrEDY0KUMKXWFh6qe07mx3SsgCHjyIobRemsskhJxoFb0EsSsD68+BoXfdA7m2C+gl163FJ
tzXenBLSfc0+vnGQQn268B42vfKk3t+DRcZG/lPA3Jm8oNCXxAluujj3bK7dgtDeGREW1uBYKkqj
XLHy2k1f6AtFpkCtmmTMjoOukvnzV9CJi3FSyErO7KylPv79ueiQZyo6aRGci0syv5+17GPqh8NX
2FU0M/fXZHDnZYJyl6VbETn5YxaKUVcMrqkvwNa1rxKF8Q3VEeC+WTbLIB/BAsFmIBHfy7jW75Df
bV+q3rp2ZPkCp84sWrZZQUMZ2k4HopNKPyySWX5ik0dnv2GLRwhgSAKvAq0j558zOVcYM4gEVG9V
NXb1jbfZcyTaO4i1CZnl+/8LjgdZ4o1Iov2Fm2j9ZHrE29wOrE9HhKFQK3UWnNWQ8qU5mJNAkVkk
7elpzosKMxdabJ5WXKnqYbtDIWQfhnyC1dasUu9PuiiU0ayDz3H6ZvbL8PfCFWAqwnp+Qkl6Mxae
TRdFkqTg0PXQ0eEGTPOHlzNK+3vfDdtxipWJ7wOsEcj5VcooiRF9XXc+EDrW6KBQoiy6LcW+6ONZ
MNRh5kWCiMEtTZ/aE471+l7xE1+ETdyMHMKew+GOxsO2tvyoMkBofW1yIZyIpHHYXaYXX9D634v1
GzQ2xBD9CT0z0/UDk3X0Q2EV3DCgj5EMpkIAbYY8gJT9fl3lJornEXi7BuIrHZpfTZRQw2z7AfCt
l5rC/8LyvgqKX+jC/cAYIc8+AAxCuVZYmHwd5rhEqoQbaI7FLunVox5ggQolLunMz9pIB6rEEPxN
JH8fpwq17klo1/cPn7bnB8vEMIeqWJavcjtvfGPJ5Nr2RyGyG9gsD7zoyIBiKJMJwyWC4nfFA0vs
P1XiPlmAqjFwtvQjbTqcNjn69SWmCHCzUURu6tXJ/K5ti1X8Ggx5BLqhoCFgXaMW2twWpZBCRaix
jkzz540F8Qn4Llg4vl/oHHEtRPoBmA1gJFk/oHFYzeoqeGREMJKvscrT2SnMkOQOvzoMHUYwb/BM
CyUL+UP3bz8fwQbhC1QWJ6s3NW1IprQoTSlleXY1lm+3LPkMuw6WmY2fqhM8+R2px93ZPOA6Kwf2
rYpyLQLg5UREbl20AsM7fhal6fhJQlohscE0YoHB029Uf5ERIBmZXcPemHt2PclfH9C0IBLj2CkY
MMuOOF4k/Xpdt6Ts8SZcimp0RGZCiLcrbRgQ5TTD7Kx/S4ycLOSo0krgUFLDDu4WTp5YMKxG5U3/
HuPW28dLV0rIIro97fBBFmxIhg4M8eRPYEKE/iDLMao9Ma/RxfxWxcipzpJ8DPoOeDQjA8bb0HsW
0/1/nu0QKctrbmCl6d2cqN6XXt/iXLEDbVgJB7QuycBsKTsP1dATltP8oPDryY+IzmF3soRrzwPO
ulGtSbJcwSp2glM9NxA7hMtquKG+89bmfKCde2eYkL2FS5PwZs3Ai0SxCxpSNG4Tnu7iqixP3keR
oJnWvrgqj+3HdviurA/gnsfHb/lxzl0hrMoJruB/pca1cHFk7L6cG1FtztS95i6uixOGnYWRKk7m
U5TTC8qfuaWw48g6HffuhjoQ5yqPHMvBUeIE8t2Tx2E3fauD6aJlVwbOVn35dk9xD/PaAOJKxVG+
k5Jy3XdsdVnb8N15Jxz74/jBjdC+PtWv/lQ35LSv0sYsd68BqsN4XXkyHfdd6Xn5AJ4Zn4ejRRXB
pqXuSRU+G216ywP3brRAViUuVXqWP2W51ayHZXxtzCgOfli+CNkGu4c4bQ2nD7Qu6qYioh3OZuSY
dTjl4RwiaeBN7xDPOlf8VVmrmTyOGgiVfPUHW6k1u50/Ut96gBQwloB7PcXSdKLX3+zip03yEWg/
Vz2g6oZjNl2wlaslzltelUOgNoDA2cksYN5GxBZlPydAAwetD9D6G9FOwmnfo2NspYcNMVWP/rIN
1yLee5t1LRJcoPNPkxenpXvf/RUo0OA4ojrKYdqcrXn5PF8wMv+0w0b6ls2UIljzPSCANL5iB0GD
tKlImlz42A5CtY1KqAfDCWRLyC+xJ+OMN4QF08X2SO9UkNfMgFU12Epw5G51Vop0Ot6FrtklW4Q/
L70yhj5icKHvLZWHokPYUOR6iJ0OTPNMzgZxL6Sw3H2OSllQnCzCnuIyPVVeuhNtebZltjzgaSnF
yNqRf05UCpLnVXMW5p1UNhA7crfxcKB2kQVYVv9PI4Xq6K2RXPDqFHg1yOf2Lbwzm2IR6cFDs6vF
jS/BYCgpJAg/gmwWmRMh+OBzG9p4ux70CIhKA7oXr3qY68mqzMi6/KNgmNYPLVD+Ruwgt9eYQBlJ
br7FvHEvpbsR0XxhrssIC9jyPzbd+Qo0fVOiErvzKud/IL6eMOVKLNdEmoeNZORcd7rhOOI8Dlm6
7bPI25duKsSrK8pQQ85yyD5LUVB2pdzMjj8QQOKaPjo5V2pd71L0icyNpzaf8+44rn1B07m+TCe3
2RkY1zCRoFYLWKyCO35loqv3PVnMvrqsLj1I/1G4+gvnvfspcOGKlX2+iGZuFS1a3Zwsd4HEFWyf
gxmvjJRigA/Itfe+p8TeHWrgpPPvl8qka0BmlbEC234SHmWKcs74v4Pl4du4OuZjtnzjyo6zOIwo
9JT9jLtLR77CCemHIJEry0zD1q7OOJQpxLufrIu67T/seHjAuUyZ/XjG2EqaRJX1mDHAMT0JXawu
31c64PPsXE5/NPL1HfwEKEZiuRKqsg0G4eOW2aHTQKoRv3uq8kxBqQK/Z3G4sO0RKkndVvdD/8+H
9fniVxpurhCXGc/Q7Ebf1o1W4ZPEEbSNGCtav1htfE9IcHVYQq1IvKilmA6GdLA4qkjuMdcPGPir
A7emrVNsrjXugJMGuqoVP5PvvCxD0TJ6wJA/PVMr2ytzm8tzrUTnqAgn26C9X5+93jQjVbbKa6KE
edK7OqH/U9k9E2gmMo9BkHUgHWOMjYhdJyfuZ+pGLEYvh5Hh2VHa9Em8myf9+hJEMeoMjVQbTb4G
W3BKqRLPt4xqXl29LSP1xBdENubwc0MCYy0YKBpSKYwKNdqzS6wSfZuj5SXvw0MHBnYzxyIYqPqZ
oen3LWaCJ64lkpQhO/AhU1/Sm/3FHoghVP2hzfnyo8ZAMzVvR/bIDH6hF8SguIjKyf89XTGVihV+
hFSpoa2ZVZ+MkfV3o8Mssd1zgXrkvSVS+NCaAxyqAD48bwxGkXef7+BqG0XpvOPta9pHI3x0DI/q
DIp0UQEDOiuKmQvAFYmyMJHksnIVsxhcoLs7S3W4UNPIEkkwS0YRgveYTyIAa+TqAc0xTkA1KsWl
CnJwFm42eWr5ixO+9YYLUfoHQ/vifJnxsQ+P2ri7neBm2GLNSiBnGboxiKh310TNad0iJlcfHyhH
tYCmhCahLujP3LFm0sBO8COrxKXppVGobJsqelorOifFGoHvRcWdfgNHUgaVM323/zrvR8VQvZc3
gXl9ByJ92Yl3sFY+csQ+/jCi2629MFez13P3AuGFD+xlr6yaTK8dmBIjTJMwDjo62u4eThS8VVHJ
K7egyRmK4R2+1GyEcjoVWgkZ5YnnZyowNfLPOlOdHw0haldsY1+R5YIcEAWwqGMGVVgtbZPYY0Zr
5aOjSzGk1auzeG0a0x8DF5o34Pmj49a+53K7bDqUE4ot+Z8tzz4WifrS88bvzY2kfri5e7zIVmdF
VSRDaV2hgtCI55SzovpH2H76r+4eZ3MpKylp6C8q2Oe7jv5qp7mNXW+0Hgc+6powH5Y1P8h9Vu84
Ngr+GWW+TNMi9PkZjRMUfZ8yHdBBPbhB9AI3AgP3fVrpV7mEWPxfeEsIZLt4kj5QG0fKzEenO2be
bS7Ib0papHnGQCgP5gLgoFyQCRRMU/b0gfhCfrES6q4OUwns6QDSB8XxQS6EklP3kHwZZ4+RhXE0
YVATMKSMP5NwsVfDv3ulrXYrKWwSuCsGcrRQ58b597wqWJXcxVuv6BjA8ZINErEI9zWHiNa9/jOO
L3ivvSIWEdW8P3d58AD65v214rbETkYcfouVu5MwoICcX5mFCRV1BqNBvnyn8Sfr9z/9qpuHO2SY
BDm3kU56qRWRyVuTSAvrusdODIEKI1urf+3PjxSr8YiRtLqBmanbkyJE4BUsksTwbpkpD9bZQOyZ
VJbjJ1qmQ0uzHPWuIy2nFwso6/oi5ZQIpyn3kYEE2D7+GxmBoG5IMRo6hGK95PvabevRl3LFqQ2o
d1VtoJLn6tEe9zSfaYIA3xDqUVAUcQ1rHw7k31/SoLH74pVb3f98bZrCwhfdNGmfxoxs/gOnr0wy
DqM3Jsin75oOwmJOYQ1a1J9HA+ZOtqDjAs4aU4kXswOEvzI7saeN5WIOUmDLkvsYF1Hm8fSqOVuf
90SeKZczhar9aNb6/psiTrZNEJMkSRduzLh4qYDIclYfSj4ZqQ7UqT3MbgSWHLJNuTv98MGoKMay
ogSGS+ZqcrVhnX/mNq3bT6V+1huPUqMB+DqeUNIED3+HwD6wdMFHu6M9DswSkByQE5ynKxvi0tKx
n4InXN3l0/CwJoEEg5jwW9emHVZa7JwmkLJyTWh96gQ4w7d1ss9sGAXqCP6RbsHByMLmfGqjyLBC
1KY+fHVvwwxGDqdVCeeIOzHBbpbgJgPrQib8vOoA94H29FiF8k99Gvca32uVut9oDhXhR0Vil06Y
gL9Z7wZPUEP3kWSgkq/mWkPLUp+4VDi8FFcH/9JWHKnMGJLYWvxEPeh/oVIdlB49gMrrdrWZzNM4
PiTMyy3Hg6cWCfN387TAa/D/N/40HveRu9HEBrHpjrt2s96ljnyz2DK3x/bfTWMEvglGYDwpBF1x
XLViLs/vE2v39FIuq9gQR4cYQX3Z7iMNUOeWzKgWFsUgDnGbxGK0WiVb2uesSXe95tpMDAkmiHJC
sw5lN5qzqQPDB7CigrJn5Q+x1QE8KhcY7so2HVaIo9y8ijfp/NJbWw/PKiq+zuby0xjcW+Jf8p86
lqIv3GzTLXI9XDB7IrxIZe9cppmfDTnD8waDZfK+mMFQmbhP9BOpyK19SxU2KaoS/qoyOtroIISq
3gKsJAh6dFdIYPaO+Ec8EieBvyRFEF7zNEIGj3ltiQlB7UiQKuIKuoNpDQVS2LEXpK6Fv5rhBitQ
oLT4H9ckfEWSpNvuXHE3wBquDjvwpE0OC+5xFHplSEXYTiw/EwwmF1HRURnpO/4rZl9eFl1gszMr
WUHgzJsr+RCqCK5M5L6i9N7Tbl1SV2HaxSmoh0ZrO4ocLSrIUOFhNx4JOLZV3NThFugPXNcZxYx0
vhIifbwiNNT7Ik+u+DLIzNffRR3Hpj4k8LvRYIOudlpihCqsjzR6uix7oEPV7s58HFADbdX72BTO
OPybhevJWEgOWTdpHpWQyls2wdaG7pc96iQemMZylLs5n4pL7yJ3MeTXowpxYLCBMfkZ3+BZwqU8
BAOOPU1KMROQ9XkEwAc+aGCb2pkF9TnAe1RcLnwOKZXM6mZge/ABZCqihFaQJFJEjSxQvS0L9o06
UmZero3Din9M57OZGTbUQ+iN02llb2SJnzZ/nMLOWA3c0YOcGept8zmkgROWgmBTtL9VSyxJxtTa
nRV+YY971gEOY32uj4TML5mVm3EXqbq3k1cXigyQoi00/r5TIrA9GeUfL+6ofIVkmR41pPcrNJ1g
RFDXKmfHlkQJ/EwX5r5kzOvppNYrMXrtw0qcUyYWEOcJdLtNXomIpE87a8N4RfjtbEbCXy4AAimb
W+RaMa+5y9R61wd7DgNxRd7kyTP2186CCkm1Hzy4FmBiJdUSgB25vL9RV2NnDqQyzx3RrNGxQ3oi
76qXG9jRcCUYv4exIwwGGXdbuaiDitUxILN4DvFMLr+4b5hHjL8zdB6H5viweGQqKeRetRPQe6++
nGkyUMBoVCMcFxOqRYzj9ahszm8l/I3RInYPBjirtHPsSZQO25GhoU20Xblm/4uq4i7IT/rFRTT2
0QMJynSlOrz1OdmuRyQPgdC9gXC5jgHOdykJKm3Aj2NAJ3/hFG4hjqYYykA81PZKve64QCKZBdr1
9YijVw/EAa4Ta1uY+sjxa0AD9/eaZqmGgj8h4ZC1jN5PgYkwoyL60x66UPIpSsZe1v7ZqYVyONqJ
1JwAvXmLpg0r+qjHyywFLcQXSFnLD4mkAs7Lf+nN62UV6wYKtHjI6GTNX8/s0LIqULB5qyOdgvWi
K77mDkJWLEvZQnIpQEWR2FYXPJMPaOhdtF31ND8S0fV78d+GN7N2FgHr4q1XqW4NlKCzKpSTHtw5
Ercdhe0l5e1E2+iY6Pvjs+7cPXyo6m6RYiBtkY3qDev6f3dQkDk2qsynEihdiCWYylMA1Dwa6j9L
OJr/5S3EbyhexSJh2jM7SCxSF7yiukKFgRqm4r5F08MwLG2lD0mPOys+F9TC0CAxLXOAVwbO54Wl
25W6I8GiET8DmT6oUedSVRMDGotibNjzur9mKz25RZBo0vEwlejg82UG5cOKZaYvA2WsanyN7uqP
gjJ8w71+S4lTrQdJLmNgAAezJ+EvbzsF6n9SstPlJ2d6xBXM/fQy9JgwUKvppsb27JxWqGas30Gv
3S7k/ZE3FKPEy5luk36vkoL3XiHgN7KQkPWD84faAhFAXDTUHo8RyjU7/9dz81dbGG0XVeJ0WFhB
Tt3+0MOJDC+p6oCynRm5fxLZ6C9FYew57vzSb/jMP7aJg+/igbVfMDEJKIlpqcXo0gEsONyCfGaH
cbCZ/JM7dFPm0Awi0gzpWgpa7W1t2o+FciM9PS1YBBGiU+ODCBbTrvOuqWuVQuJ1YQs5EEhvmcG0
jRFtkM0+GFO/7ONR6DARR5ebK6kt3FtgD3z06Lu3mWN/Vrx/+uwGeevIABajYn3B6ARL88TMch1h
n0djpjtbkXQb4YvG8WMcG3fGjgMAlUnYDuGmyPz03f1HUrksvTfguGazidFWSVUpyAuS8GfPSl8G
GU4lrUvUPoXwDbgBywSxhPVcNqZ05mkSt3yE6avHC2BAu0CYA2T9lLvC3dR3SDb6nEQiRsRlxg2E
BRKnavfRqeDAV3IinUq7+ZdN+tVHf4Oe1+TF3KN80Ezf5uOlwqxbUmsflBXZUD0RtKyJklH2TdWC
U5v+jq9A+TgfC5a9w58fk0xQs0teSlSdjiVbOv6gDkk50/mY4J1k1lktQxB7Q4ScxdDDqcP0LM1m
tk0HJ8sx5brt/DsJSlekrhFLi48afLkxIsZVbURvXuJX/T5j1YPpmq//PsKKZMAeYRf0mpApAUaJ
BB7lZ3kDRAUahkj0Sscw5W3r6wHw3CHhkIqumSpMvkkvfKvMKV9zEErFwsAJxZBigQWGYrEr928s
x8VuP9NpuogLPSybvukju/75l4At6JvI08/lgnNqUomxc4yw9MGF0PnJUKE0X/ZHKWpYZQ6FB2JL
9Sx905Gex+DfOmDWb/AvEGAxZ9hN8MLr31j4/WV4M4YUsSNw5NhrurxzG0sELJ+P6/iQjUHPPkYi
fISdFWETs8pG053I3GAyoUzrAaf2XQi8ImYxV+LoqQ/yp+97kCm7Jzr/jWFLXJVC/ookNkTxkzzY
n1J2eiFBlFDF4nl0MFXUX690PnnUN39kEa8+rxi8dOaAu2RRFg0NAMpwZIa7ynzp3jt8l/o2h1oY
wV4lQe+1/JdXOIIeq967QtnOvymgVJxpOPqVXpsTJXHrUAorLnZFST8LjuElKOlmRPPf0LP/FJTB
ifXnENFFpQkDAhBibsb4rhrPlnqZu7rWi2ad/gbVY3wL1p4C3NA9H68Ua2os9EdBQkyxm0n+imMB
Utj0hVahPyGcuDXrTnTxFH4VYcNezmZHElhHR8SIpN/DEvkMUCG0rUNoa5m22YpzSB2V26g6n+GD
N8B5ucTmluhh+3zi0E//Lf06dK4ENACQu1s3LfBFj+cmOlkESjMmgz/rOZGiQ7woySAGYuwX7s54
PDT4WghBB7RbyMcXe8BuzIJa+3dty3Jf3cYDbEOwv89Ad9fq2HrrO4LpGuWzLzfu5M2XRFgUPKLv
7h0PLjd6+2DYJpqEhK0gg4l5c02/KqfYZ1XdtVqFIVPe/OhKvaU5ttJ0mAhzybneVkSmUFCYkZ/u
dAcNFBAeiIRB8UOMfVCpNMPeCN9tPFv6e8ZtIc202NXliKyGG0+U8QmUxbcV8w+iYVQVOC0PovAj
IHfiIgeASdZHzWigJ9OGhgD3AeMoX5jFsxe/09vxrYTpnNe8Yv/8EMX97iANJVwD9vsRZ5WId2P2
/OcN0eoTMqnoBn3kKOaWTr/3jGVfLkVU2Y02d7hcJDYsi+8TqF0lxR9mX1wqGHAbplB2AllG+Rw4
D1qVjVsq59iSECTK5Eg4BlVG3gn//H2qwGBA+7juQhdljG0hrXnF04EzZal1qOQ3B2CYkQaJvS+g
b8Jb58Gxs8ZE/OOE0jDVgzhFbxZbEkcypfWQdQTLRGdwQCMddsy0JLdANjiF6b52gLmBi7WqZFW9
0IU4cEGl3QA5+0maf5GGgyvKkHGRLZA8IvA7DCmdBDSLMyprOpJr6UqG3yPM7o0vTZFulhzWYK7r
72O2KlGkf/4peUXii4j28DFwWfyWKXc4ajBTeMqga6WKOgcXDG57x2uHof20JrbY/U+MVsDDRED7
aTVCM0ZD6RG75SX/DgCzbQNB775oGt05DDwUiAuciy/L3gDRbpSBXqWIvpq/k9DPeQut4vqok02v
4FcoKSgFVG624klGjkSVy+GhIvCeyV4eZJ82M0/L91NrA/ur1WmlagSim+P3iG8P4hLBtzP17fB7
qz7G/NYxM51wM66GqbqI9cVczalEPQY/9FBl4ITjCQgPTkoscA8hXtbqGWoZzTQkahwafrFpfjPz
RQ/rUGXR5fKwkR4A+XBpRC2/0FB1uzBxVB66zKmmb+pIlAjEAd+2x3bFTt36jtjdHWErApkF2rJ5
ua8Sol9KmM7UP3eegajGmtQsoSztcxtgV3aytg1N6COwSx4BvVaMHzY19O2iTwZpUgTRK1byUlIE
C9T2E023DQ39CXCNNJ+objD8VR0ov3Fvy1u1qQGa/LiWr4cAxM2Q59ThL8yBRVE1snkHd8e+vkya
Jt3fFy3yzmPl7li09HHLzmj7CPn+PetvLrEB8F3jOc+Y8oNxFYiM1sWcZcbBuawaMTaH028G8rHl
UoAELkqMiW2HboTfKC9V12B///p7iy9XYn8OnyCqHhvRhPJKX9Q3xOy/tZlhhAwjf2waJm6ZSz+T
dWsLhGJkZ5WO1N6mLGQ/h8vmJWLtdaLvWxf9dGgbahtB1kumDfwz/MEb37kP9FfR/MTYj+x19IoZ
MbCmXI/YhOhfLHTXHG0Nfe6PD3l8AE5WyDC8oWUBIZ5+uq1KUKwrNxs04Vhj4RifjOtyeUneAu3P
gBJfyb4URrf1FbqT4hoXBcvFsfvdFlLMLT5I7syU9No7V8tXkVeUw9uoYIB6BoUZB17EMzsXjyWe
8jkRXHXJvZcfpGrXmRD168/W5Q/HFOs4r2yTmwGX2bTQsNWMolTXR+KAzQGavKnKruzry6T+ldIU
7oSS2b/1AVFxAeQBmQsmuJIMWoU7NNLhmmcq2coJsQ3H3ejZZjbCsRdgZQKYRmLYxrqyOxuaF4WZ
LCImPqQkoVoV86n/vEMsmv4LgCMoelNbJoslhFqRg4x3aohNxyTEmSR/7USmpSA9UjFHmnBGw1dv
C0TBNhNs9nPO8Jomqs6vEN2WTcB+37u4InDaZY7Hz+5tl6MDaPF8lCpRD5f3YQpeZ3XXqa1Jdm7+
aRkYxbwoQZcXEBG11A8wMRyurqnUjlkdSe3lMfjTvZK8CJzK6SfLbSzwbd8BuZN/zCKTM1JEHy2d
zkKsCv1Sau4UwQp3jShHUQ6K549I3uJ162G7RZmpsjL3+h9H2AU0/7d6dxC4aXb6HWQ1TPKceT6k
WKN0qpkW88SQ2Lyv33bB7Q0ooG9HLhkqbFIyXei1Q3Kml76lWPWv8DS0ymZHTD0SEAkQftsZ2M61
UF5b8bqEEtOy7oc/Gko0ZtuNMHBVzMBK/f4VomYRRYksRRxMbvCmlPzjmVXwt+lSTRPd21oXGKzw
klWWgTg+8oiUeVLRBoBhyg9fCZsjmhYGgY7GkEdiiqY+a51iieBlFbwSujbj2CM/k9dVKT5VceyN
ZVBeng0UXy2rM+3rvTMzD+NFuPkTcvjo//gA243Jhkyegre/iRotBOJRYSkhOmU7PgizRxERifvV
TdNYJ4O5LMBXsg8WPTFzY1X/DzkM9sGoDGVaQ7kUJuL2YqbWBVrqyYkaIVrUQpws0CnSq7GINJFU
q0zYa+Xk35xClq0YTxka37PckIFyhGKtdpe2Xddo/zeKwShzPJuRZ+AADzBfH3TZNo6iXJZNJFlF
SjUlmve6CcJYxEPGv2S/t/rzFF4DyK9bUBK/p3+lxQqP3/4OWFho887+CbaRD27X6hySC7M3t2LJ
9Q50xG37VrT/bkGbl6TQ9NbO5sIFeymV1Ke5Stbd/sVQrXpoSBOHBu2ruAX8AaE/TWOEKmGtPklk
aCApEhnwRqtMLWE5QDxT1poCRpswbu4P8VQUPWM1dTpu56AnMwBWJamTKNM6lU6jch74Kz6LHzQD
2OGVRIPpvyaEA2M3z2QVFPffeJJapk9FXVymRZkM/d1py07rPWpNXO4jJCpZj7hIzVHh5S0mg4mL
h0JAoiCRr1ArshExGFCUpPUrKDRLtGfxANIkmkf7bar5tcqGuE6C9Xo3Qr8MMKHiLZK9QCo3GmUE
EqlrPEfrhYWIOXWqZwJysLkGs9cXcS5GLjekggHBWKP8gqQxJiVFYOghwIPrVAUnlSC+vzXJAtaE
NTrcmRCa24y0W+olA0FG4O4QutJeEyoVCCSIam8jDFhJxvD+nDFYdf8G+O5PJU2dk+MOKlUxTzGO
IZPE+wzqYecq3I+A0r+C9NzabkOn/5JF1ekWlQUqu+/wN/DQZT5IxWnUj+kCfmOwDMNUdgGDbHu4
n0Tq3AlZI+8L/GTCl+80vj/yuHEM6KyIS7BMevL3Qvltfc6qKhzbq/lZ09mik6wvjHaDvtniDZ7i
lJkISX0i7BuKwUlglsbTqEaA4znLs+FsMcd323MS816dxD//dOnkrwneKQsDjKqX8nW4cFdDu+PK
vAQfwuej4YEH2wWLdefpOaD/xD7mVCwMs+JRWJPQOJwDZw8BsY4teyWADf2CY5kWdRP85m2xLKLN
EBQaqTy0TLbJYY+kUUGzYW29oEGt5FYd5IUDrVBKUn7eOO02ptFQ6EATDOXOkGPrjgC1q2mbjoWq
6u7EaB4dCS/Dw1It5Rwpwk13ux3566Zgh2rQiwRzk5IuhQEvhI+SqVeK3z+SqRDMZn3JvybF9YC8
QIUkNYcYbtRfYaLLKLvnOH2+tVVJHX9sK2EdOjGsc+lPwwxWfaJc2ZY+D8XMll3iVyT4CP70hhp7
Sfl9hNeOhcZpKQkZL+JlKspxNDsd8U1Qgkr+N1F/gNSO5kno3d/at11YEv6wTV85GAHpwTnTvRHq
89SpH9TJuSfOlDccSGsD7Ta7fllWKMusv7nOmG1BEzIMCLhjzIcIuJH1OAkuDADfTCbdlRwaZEhR
TzUKOA/5zIf2rvrvRFDz3mRKOuuSPvHNsOMPcArF7RuhPNSPAWjCnGg+BxZbZM03PX5NXP6HQCiB
Y1a6KszSn1ilocL2eO+JIh0/BZAi6NLpFyuS6OW7Tm+uLwAJzHCHuVjWkCKkOSD1pw9qZT6f9M4B
RTMcLPQB59U6FlMs3rExX6rXVcogFUiIFb1e3GzemTpAqeTl5YbY4ngrij70BMk+3ghPZI1l6IwL
vmFp3x/XcdbZh6oUX+73X8L7EQ4BmQiv+NrLaVCdHDRb0FhHImjgspwQ1J0q9y7L1NoUgtBOCf4c
RAX6C852mN+fmM48mmjgzLndw0rswHf6hSoWywcHJmdYW4oF53sAfz9QZQxrurqv79nqS4o6KE7T
cyloAD2qmneqHayxcKhZiF3rX2diEd0Lo+kP2MH6QX0vUpOTQjKuaUhroh0g3r3kO1bA7vLJ5PTp
xDAtckCdDQuouULDwIB3kYdwXceGCzMuYXJZPDc20yfIJB0sLxMoDhm5ov26jJuTkw1MbHnn3+4v
YJ8sIEylFGDhoOjxd0f6MiXJAi0vf+Q6+v6CyzzXocbIAwAVydzRB3A6Bzn0najpbd+V4QDL6ao5
eN99vu4wdIipRzWOhEvxSJxpWRMjB0kvOaGVMRJmdD+SgUzI5bWnuT6IbpgrmsZRNNt3WgKPsT4O
28i5uX1JlYhjkjGO1K+CCBeEjr8J1+/a2j7Aj4DmaEZeikobbh/92w3prfhzUiG/hQEB2AQdplsi
g2J9sEIG6/xC7/oGS8xxKWBuUv5ffI9CqvHC2mKjddUdavpeE2+m13Sg6LyPk9OnlQLEMJj85iDT
otNgqxlwUR+xkK/bkgIGQpUE5ePEhHp/Vj1UAyx+SGrvV9D3VfTBOTvPvLl1fBv/bNDdwB/TCMbM
tiFsQJ9bRU/N8bXZ/i/wTzEkRcnIIKvMgEBMhEY2X/gsLwk3fd9XUrB8MAZii4wJMFS7o6d2AxIa
fVg6jBS6jjHb2Q8eu6XnwnGa6clGJmGCwlFS/P1X97yNGtEu1OtuCRVQNzNxcKg7ut13xvzlyKH2
b0O6gtP94zKqPAgdRR4bSSADyEoVLJU9i2L9+L0o7sm5ef8oaGXgHc1aypyxqnkWn/uQ2YXgosJp
E/7wujukSgtebObMvnSjzsTO5AhOkEDthr32rS5QyF8QamzIcUv3oxr4RijDmuBdGE2Ot7B5p6Rj
KUGpOgcoUz0So071D7zwVuqpNvtkcfgYyskMAkY1UhLDdmb4YnIoAVosrDDumnOKelCWsQXEHvL3
gJ0eAFB/QA9hHmML1Kvb8ApR45JBR4ohDHbR+JaHzyemWO5upANYsZ4s1uPvK9Y91zSKobO/+E28
CRlOIjSmYwMFbILUj7ltXv9ql/XuLdiFVw9ehGkInUTub8IT5UNaiu97FE9jjMtt1WONRg3z8s2y
ZeyULJx8bcpItDnBI3mhNfzaAsEHMvD3itkYnHVujFhT58dmVrJ5Y15+IcEfAx/RgfAdqap6UeCm
L7qtDDUfbeEm/N2B7fAyOTu2ObqKCxO2VpqphW5s5hb+NFvYoghxH2lJDdg7XuV7KXF+XF+zSL5r
7y2v0fBhLYKS2Kqox5zk2W9F8KkbUUeinJ//pmjPF8l9vj/fHKd9ZOsJIaN1vN1IxxFAY2kkDcFF
zf5urmBW/ly3zyN3+3gLwqaXxF0ktSn8hizYwJtt4RoTi4j9U8skQW3XQHAIfDs/KUPcge6h2te3
6J7JNDg7GVOOJlsJufQtztr7iy7UGl6WkMrrSNs5WUDgFav5pIW+fRloowPYk2tIWHHNTrHvXWLC
3s24gx4+A1EZBj6WmIFD7TEe7ifSuvK2w8q1QzfX4FIaBOaN7w/aSwCnJPNb7c+CKDcBMedDDx5b
NnA44rLwg2Njvc57ssACaIJpHJ6weuzIVcCsXU31Sm9pBYAflAdJp4J8AZyrV7G5X/H7RVpK8okk
7c0Kr+hLj7ezfHcmnjWRGWjWb0mslUbaOrg0El6gOubCp1jNVS2Hp9NstGnxIg0qHIxT5gpmYlyf
NXV2Brs5Dt4MRhP+NdQBRAztXWTSIlA5Bxyq1YjCSxYK1f48BvrgBSsfJxBt7yeAmTpS8kL+Ta/M
l+WHhaQ6P02Z17QaqeG3neXXDg1bcWkg08+AocTBZHUP+b60OzMHdHp6/Et3xIEbx0xSPhV06ITq
8tj7hCD+ZA5vOaXfG/v79z6XhTniktFMtFqkdi7jVF/XSaT7nTGdopWYp3VkWhqjsHOH6os9zn4b
GjRTkI+QFpubgoYRkExZJHjXEAQNXZRCqOna7nYptWxbVy+2NiUX9ZBz0RJB8WdpbgD7E/OMDWl/
gbxg9gH7mAduVUDtgld/3FOGMMg7iXPrAhIXqkDr9Z9zL/cQm/3OIS/QaIDS4mU+3cja9JCohZl+
hV0vDUuYIDove25CM5pG3XXouO9OKZHzi903h7kRfDFznsQCW02VMQGruXOh1xnkxFso7w9PXgLu
VqpvzlVrz2kkxX07bdd57gAhqRv2bd1ybmhaHipiO657LAUEafQ2NR/sCht9rTlk82lLgtkpyNwE
v3/unCnm1qvRBycHsLasBVh6rNMSdqEBHqwAENnaCrD+LMRdJlUccRGTCS2hkF2DfGIBcg6Mf70q
kb0ERKFX+9MPfGkfpxCM3oOLIJa5FiBRSSfpLUXLr1c3lWGzbETz4WURQlDcglLb0TauIZwrlwep
1zjD3zlnHOHbn8J8ElPvCvul3uouO2rzxQAjK46QM0SDK8t5NqgdMFJM7+m2FUGBpwccq1yy1wNy
ihF8ABYBxyGP1VD6Q82YE7G7veP7TBjKaMtTNjGNuMirq77j/S8af64HH+IGlKOWBZfmAOeusriH
UIe6NspP/vxn5sWj5wmCIYD7eUkA9ZsO0NOsVzWqcCl/MKlMHZftiBjZBI76uxm5FKMKCNGFCnDE
v1LKVOx2yv2x42Zwr1Lzn+OV11ojqToYl59rT8tuq4rMHP9X1aP6ZpLw0hqmtvyKhTwVxn/Nxx8p
8CLqF0Pa6bkyL/OL8aPOQheQ++bX6L7ueAI3XzAfO+o6y4U1/DVFreP6ZSsPWkVBUdbyvz14zHgh
A3sBKKSEtqDO1nTx+AAIZz/UiE5mYr7QW0Z8ilTc4IbhWa5ySV2ahlCk5XIgTfcGHKsv54XixBzJ
YDSCdhCaNahmkvPs1Z/igndrri3tYZwuevg3YjmYbri92T37vpiDNPO7++dRIa+K4XF4yPyk3PuG
hRmFNSAR9JdqqT6Uebc9w9ps0dfLXaMEZiQwlv3UGDU8nt/bXOUoXC+QZWi65r4xXUTpcEhm8CQ1
nRiRwr07MrmHYH1fjaKDMpl6qwOWnMeItgrkw2ZaJrrWTD9UcerWexBb4wJxZ2nLSe5vIAZkrVYI
n7SGEtJ0PSR9MF5Y99DbNtpQnZHE/Z2Ltr3NQF/47E1pl4YVkK82Q/pBuRAAM/BZkFDoNCR2rMTU
p1dDsD5PWDkljDW4yENK1zfTWMAeSRNLvn8m/3nkA8UtARStzLsQ8+lVXw2bXO/yZYQwGH7ARo0H
EMFa5QQhe2LHt7Z5O7bKiURLc5zL5v220OHcE0h2z2EHWFu9vZOGrVn6GZ4+4iToG0hp4W/r3y26
/ioqhIubRqt9DqcYPuWxm8W83Sk/brcVR+V5HPsNqK0ATwv7OLPHyB9mgrBt1NxnJydTMkhRoiJQ
gohMuItKM9J/MAtz9P6iQYlLWjnlgyV7f4LwDBf2mWTZo6KMknYQtRMjGxMfU4Y8aIuQ+loVarDi
eK7dGzfURKOZ0QGVkqzErSy2m0KVSroYZLbSMaICB2OjMmAieYqV9O592dO3poCNC0BQLF+o2WUI
VESntZ6qUYp/N8mtmQA4I9ImOq3JPfFB1AtsvrJQDhOM6wdf3bOyvMcBgDAlTdXSq3JGEBy9YIuI
h7gRQ43t82GRTXTqWufDaL8G8Adyfw6vn9Wi+02KS2V8RCtfZrtieqDyLU3u6FQahktHoBBImXRj
J2PIWEwZFE/Q3MPDpXCgJJzydbT1fkN1/Q7BWHggxzy2rCa8a560Qf2V0TlXRalpF14UkOJXQGQJ
8aYElK3ttYyWxHlvFLGuAmvkK6IkG6BDzVIVsj2YS49BTcJ6TM+QXu4vMTP1TbH3TF7BrqTcmv5M
7TO8DMMbMtZ3C10RLlq1TU0HbTyYydIUjUeFgl0l6TPI8zQtUlayt3e6J4/2QyC3ypJTu7zOxapC
WJzxut9CCUrasnBWeAewpzjy2FboOp3FKnoJJhsKzFTRLP/giVyrGn3Jxb7jJMlFuq2xViM21GcQ
i9oqjYKaF+fCN6E65SsY46RMr4xCZ1T4h36/Jg9s+0Nu9qhK0JJOndeFkQZVt05QTDjXGkmQ6zUw
AuWBG3YxWYhyx+F8gqpJDm5lRpRIRBZAuyd+dRbB5jzHkS/5vm6f0xdP4kTy9sA4rjh/hwJWRr/k
CP/xGPVi8hWQ3BReo3WdLi5BMh5zHLCr+WML3NMJN/6oTSXvYlUSLZmqOEwtvE5nK7bUhRIkYoTS
WkXCodWP3keEjOEF9w1Ue7C9H5W7l8aUzBm5NB27SCPth2cQzAF1gi+aEpxKUC4Vr2c139ujN9Ai
y6q4Efn/XKv6R32RDcpyZJR597iglDH1Rg+DveFsVhrSqCGRBfEgCgSIcp9dlbXirRji3rPcWvgF
CXbMFQm6SRw3Ak2i5ukvlQ8WuueKZqFPnkcsJYfM1MLyXPdTteSPzF4CF1ah2tpe6bZjKkMjThWc
3eZcDLc+iKslaDxHVzWrtcRMn5WYtbxGd2PaaxMkZdsogcS62r4iwwxC2phtfh7m348BH2pO/GFC
6fxVf9R/Eh6Ia1IZ2puJcZmSWH6aXqT3QBmSK2SrB7Up7bZkqxTGRjr9KiFDKzFpo5TdtTgVeT/7
evr8KFhi+UqeHhdfZkl1L/POaf8VH9qhRvEilL4NgG0ESJdQxKyF/zaIz6lNzOpUWOj1Ek2cVTmF
H9m8b8Qi5a0jvbjeEjaMcmJHNetGOYZFJHetql/ZBNmSEdrumS2+d82W5RwtWniMvl+NIY70gSc1
O2ZBV/H3GVMPz9mnQ0ZR38ILh1iW3M/GVvJ9B0k8TCRmWkeZTXgQRr6JIMD0PMx0rbaiUxgCMDXg
YCnhiiyjaN6fqYU3k/PZhbdhFeYAcHGJR/Muuo7Idi99+laS4HP4hAGB3wr/TC2lxBg4qxf7yyvq
PaPXUWqdNSiYf+ZR
`protect end_protected
