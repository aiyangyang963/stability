
module Qsys_system (
	clk_clk,
	reset_reset_n,
	pio_led_export,
	pio_key_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		pio_led_export;
	input		pio_key_export;
endmodule
