-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TbAowgNOau0yzC/fEbW2D7QOZpdi6TR3/gZScKDAkUSXkD+ct10d3itZ+0tDOg+ZlsVAM9YBEmIC
4BwIfJW7tGpl3jz1LrXhxyXcM/JXhPZKqllHJm3Hnfw3CIVJjxt+3yUhYEVAB2jyY3eBZ55K8RuO
o5p40SAiCDnrzhZW20qiGtnuBEU0ZEEXzCSNS0nq6vTWJR1F1bVsuJuEciPOh2S0mL4u0/Y0qAF/
idMlkElbAuG++h61rq+J1phq2j//BoOYCMWP0LhT64FYbc2W7nQS9QB0c9APJZ2QA7Dy1qDf9sr2
z19qdl7J2gqVtC7Hplih/7ZcitKfLPRsJqyhQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9488)
`protect data_block
LQsxuUU1LFSvUJs5t0siCbSTH5TnFrO0mnUn8OrfUtqF2qkf834nM0tufcCgdUrVtzK7posYA7wx
nYjPOJX6/GK10N/tWO7GXThs/u2Z1nsxGHnsINqnWg7stDBJWPU/7b5rG+6j6T3D9pPIEg8AK3Sw
SP1bhRQbdPvBJGJHvHI5yTUTUGlekXCDoNMezqky0Reorh2GDpapQ/RKw2qn+i0ApxjGYZZb0MlY
e09L9cnF9vvpz/ZxhqFgJbP6Y7lAgmQk8L4q0EAp9X6Av0ZoicsVM7eSw1TCHl6oMPWMRg8oZhZq
Yy1D2hdB/o2gl5wcThc7kpl5EzXi62DECP3CbAe9jqXLClkC08IqTRogF1WO+IJJgXOhjs/FRHfd
S6aQkVGgXRx6xFix0nQgR/4HacrW1yuMY8cFFTDsVIwCoKzCBw50z458zvkWoJTx06l0EdcZA1U1
OU+t+QudL8fnbslhAc0Hga+csFQ3FakRT2taa+8zGL9Bu0IcNoxijPsi/hwGz9+s4SwV/W6gokoZ
fwBR8H9kaWQS77RPjhjoZhCwjSVUCJRPDbxVafAfU+zyJ6Da2w0xNfXQWCXE8vKJGvcSeDCpQwp9
iPf3nDpjsLYaaK/ZCR+bNzeBZ7hj6mNbch48zjsCJksIzRfFYdFGrV65/v79TW2BorFFWF+vZ1B2
NlwZutzAqFv67OOTPrpTU249oFwOm7GpuPrgyEzN5rAOLaSumMhw/kctJMOLUwaYZOSdIXFiZBLk
GvmnmRs+s+jxo5Vr5itecKaDi3mb32a7L+Zf+5o4cRRCdr/cEkPnEcNG8fyWvXjj/xxG+pTrbrVM
aQ3rFbBy+JOV9y2NP9Dxm6UExMZe1SjH3qdU4ZOpZSNxOHlI7b3UWc5GN1gPOcXZunV7FYA1P8ph
NNvu1s6dLK2yEchkDoUv+PiHWokgeKJ0U6kV/70Pnw8d8UNgjcEzGZHztiePprrRYP90W2AragHz
cVJCyFfryeW3Y9IXnew9jfnFcQG3z5B512/9OEMdMs/PEuAnjIsVbhlnQVuNYNWV1ir8dtwsFTgt
uhFpmIc+q2eNQbut4w9dDC4jevNQp4x0YIj/difkEMQ9LGBlr+pHrLm64/H8GM2dPcXztvTfLzVS
g3h9944sOd5YFzGFj+6M7g3uUMEc/nYNgeIDYU/Fepp7Aaow1oZpjU482H5qh9Ji8wzwxJaYf8Lg
QTocgJiaHXL7UHSR1kisnQrH1UliybBpO0exMskPG6PBXtFDak6AFd2Eju0FDH9DMSsXMIU3ydXc
RZ+3Te95M7P7+24v7NnfemB2EOUStZSQ2k+pmaUh0kkJZMr11jL9wMzL/04cG4KC588teTfquNqX
kY/rljhrj39sBSKvpVrw2UYfR1jQyyN9ujbO542apHktk25voZzGLt+QseKPj9aKr1Y6vHmaNQvF
Jn/n39yFpVgmQ6JhQwMamcu2DhBw8ootXeA/bfhYjeCQpvgaQg912ed9NBhlEGIMTxV8MIDkl2J1
zbSbfI3D+aOfc1rkeVjEAMs0obi9OGngOj4rblUg5wSCz1b+dRYAsDLA4ZwUhxLGO6uGQ2q3tB3I
737ehzIkO32hLm8EtcqkRSmxvaHcFFLAeBuzpVPp6+D+ROdikrLP8ca1i41ks2Hkz+46stSQuKCv
0z4iSYLUK3zoT5fodMq2UEDf7UpcNRrkPjdYmBkunr1I6+rpYcB2/wyDb6rPycf2w+COVA33+6Te
Fvw/Opm8Ayf+tYSEJ46hppSOy++fekWsnFd2A3kuIBT9xaCNmkar7aOvWIJxnGk9FftKbBw32302
sqWRXkBaV3JzTAjFhIqV2V075IhiXU6BRnGcOzpEsmmTtIRCNpgpLvIaWNIxlrYWJvqH8NzwoQw9
eetZRpXR09300q/mdiBId7wiwdLDsNKQuePT5fdlxmPh+jdO8eyQmelHBIvb8j9DofAKGSOEqAp5
xHOlFuu2w2QXZ4oDK3E8Es6mYUYAef/PvtMh431DSiJYLWaB/mOWbsVdWCiAZI3lwzxYHpKYrfow
B8CXuxcSKLfTooZ/qFvVZrWZQqw66/uPCekH88YnYO0M0m99tN4QHWNih9XIOT99GJbV+eNR+HkS
ufsb3atOufylemGezj7uLU+ZrNfptsIYwh/K8i+wSWoZDtcAKvUgGWhrRxoyAdElCLwYLXEfse9B
FP+4IJK3WpGE5u79leyxD0EW+vqGGdG+B0XbDD6+p2Mqe3AYN5T3qQLHZkxmodxIi0U1IrPD33gP
6E7G7BeSaclq311alVyHSlSkeoON1SAnT/3PRD86cpsY1nNaZDKf2vixdKRJOwrg51ATDWDLMath
RYwjF19VB+ba7gAtaZUh/n6mNIOKBZ6SpXUSLG2E02rZRiDiRKKTDOsL5NV4pK3Kjg9ttQyYFG+Q
NQDmbMCzglXcpbh2kLcC//AMxD5V5STT/MYT5tGTbCLQQjH/RsVVH8vjnEriTTDNSK9/R/gEZSo1
7pk7EXTVMfre2/j690sxUBbdvCh+kMmQJ9FkAm2beF6neTmxXfSWLMmshvMpvm1GSjsqo/RBiEHn
7Oj+grT4CdZM7d0wDjqkn5cCgpMCqlKTulZ+EEJ5eID+i9P3o6bNJBQ4pstwRXTO2QXiy0iN8WDp
XVTNtffVCaJEaLNgSVrSk9curmBCBcUhlr6MMr2PKpEB8AQioTGUVT2fQCb+JoEqm4yBv+iXNekE
yR5y/D0tcZ8dU1rd1Mb1Hb10jtuuZLoMuncFlDWhmRmDrRJscHjax6G/vHQnpPtiiqxwXwaYJZD2
NJRmF3LBZeGfffkleYBSo/HotnuH5pHueHG85T2LRBxH7qHADsaQZ//MFq56PdylfNw3ungcSYC1
aljK4jWrvN1PgpqWTbiFAKsI4005WTrSh96lF3lJhCcJnb1kZes8G9iafc1tb0XDYQ5nvuSfmElu
hZ+d7MWC5tmIrggJhmXXkpkgpEuNckP97h6JxJec8b30uDGRNNtvrxGeiruZ84ghyrhJOPbWOHy6
WxXTD4DmL7FJvptLa4B0u1FGALDIauN6TZgEbZmWzTnCsrVHBA1kpk9hvY/rQ5/8mZaC7SWVpoNM
FW3rDWT8y93e7LzPYseZtojzg8jSP4HLgVojLrn+1CN6cCjLJcjRPVoovGXEnMqd4hp1XnS/yRY8
Im9bUX3wwKvf32Vy+wgtHghlKTNYUhrbDnT00IL/HWPBWlAms2OORLaPZCQiAwLRutGik4F0HrKW
evLqLZrjx4tRuot5DJbFVy7Ov0QfBZkqpT8BlzerwzL3k21h8s1rgaEz3AzCw6Nj/xrWxidAL4mF
sS32GV7v7BIAttQ/Z+T16g7zpf1w7r7N5d1RETPCGQjHSSY+m1Nmtv8226lrtzpVSljiSRL6iMzh
T1Wfb4aAisVLUSY1bo+L3yN+OMOAC7Rin2QAJwdYTD1uorLgtJE+t8Mr2NFuIeB4sFN9KszFARjK
GoGxsFYVldUuRDH+FS2CcKGRfg+PqFpcaTqI9h31fib2cQPk32iWDkdzrep29CDkMYiSz0dJMT0J
Gsv1WBQqS4ty+U3wUm60h80t8r7V++5aGdW4KJyLUfFqRrALOSEZFmAnatwtdMrOCy3jbwc9Kium
0G8EQ6u31rvqjPah9NjTCEVmVbS7kWbe5DpdprJGbjXcfSqrsy8+pIyuv/Pyo71JUhYtzNBVCv5S
D0wXpRnhhyr+9VYfCfqm1s63DkYgnC6rzxPihIctNdasy4sXUQkjLYmN0YLFXUEHSQNl1djpan48
USz0nRsMswSiHEgcsPSdfgDh6p5znbKWAHhTKq6oAiVEft+CKqdspmkarH6JUgO4YJkOM4aUJ9I3
IXzn8qD8ycqXDB8Yd26Y75688WQ6hHFM7T4sDk8WAROtpfSvLKDLVhHOttgCNbGSvBIoH16ueNDp
te1o/0zL7VIbDdzfFkFN6B6LdTi5FHqlf26rS7Y1oyHIl4OEELRHKn4hc3Bt1Oy35bp+kWgthMi7
/GawiijLV6vtHRkIAE1UP7kBgyZOeiH1Ey+uCq04MN0lPVtsv0PmoF5hq8zfj2GIHY54riaP/9Eq
UBxOHj5T1PTmqAppUflg7FB6l4fVH/Qp4ja+e5gz8omd6TuaNIWM+OpOvX1o5uQM38FpZGgVrrii
Kks+ZUglpgQ2igCGMRISCADmyn9vYXzvfM25tHDnxWIFCd5FS59xF5NGZny0Fn6Krcl8xyQ+4C6l
IJ61Qa3/DrprRzQa0TObw0WHWM908DeSIT4YMD301cDESQrgb4ZNsZOyYTZefzRcf+Yc/JNHAaOe
1LmNAWl5+xRhhs3Gz7lNhFK+UZHkdpGdQ4zPvYKrIy0d8r27OPDKXkxLRFAZAXAN6C2IQ6K5dTDS
VpEhIderSZE6Vd2+cLoe2iJ1lrH35pdBtwjh8fhq8wMPXZ4g6tvVwB2uRpe7C3kyNzGdrPYwUqap
3CxcZ86jcKRnxD2p/STDn1ETBuD9fOc2V9RdfrntZKXZDuve5Y3eb0ED764o7NgBOGjr0aVgS/T6
Ly+GrH65gCoS2TpISKIwJf22wpNr98yTyoeO5QMUxuPbQJtXWNEBssklvUnfXOKK3pc4pVAspPAU
p17y+cmw5yf3aE1R5cvcmyEVzh/TEFS48t7wyqtd4aN7A18YcgB/b3SDSY4Wo4ra20duzGmOHg0N
FpveYKrBLEpkQbBdfpJzTbOeADK5Yrtkzde2xn/3vBDQKb7n7HagS6kKLH7KoZ5d6/g10b7wJ15F
A/KPOpd4t1hxf2kbzx+q0WbGP7Y5iAkYpqTdEDvqxjFZG6t9oobmLpjxUqyOfKWezzq4VMvQNS5h
bDAr8jyasVfbq7xxd8zjG6AcCkmJVXHyLxxHloUYSLnV5TmjNZOT8oY4Lp8+7uL8RmzHcsvWs271
P4bYgAPdP9gX/Sz84qNNZv2YBZAmcibXh2eyvkH2qd+Y+4k2lAMt7mzd64TFP/l85BechOkKbfIE
+HGM6oPGkEJpF4Is/lNrNXtsMVjmDjHFMq/xvQFbH80jm7CrLgR3qCklkaUiLGCslGAYacNTInQK
fMU4d7DpiYzeIH8n5tyz3Su1kJxjagMSg/SHMJx6GjejUhMhvVXwAJaG+cecpEcu6skK0TTbSSPQ
wT8P/0lNbg+9ly9WloWMoBOBzRu17/Q49EgKCy3hMcBKGlxtO41iKHDeXtZUPDmnmO1Slu9u8MHC
ZM7tegON1dQyr0rEBsjMC+K/xgEX+7J6pdWAUWU4cD8LCCMN0sQB9SHP+Bk6ieEutu2EGfrps7ei
yhU8UEMvQvkqkL4RBCZQV1d9Gbiz1VA6Xf4Ax3mhz0T+3Qj3G8CLhs3sRzPLXH3yba2j4ToXgKfv
/hMEOyXEOhqn+SBd3Uud8thbZ6DsWwGPjLLl3oKLvJmiAV/Q3xEpCH+Hi9SR7GDANnGqqDsNF17Q
L12/xKQi59HkQe8lZs1ukORod/8Cr79OKf0EdgC65lDUJiXQhYOaJmQAwPM7kcEyluMEnC2YKMxH
3/ZPCfJFUISTjd0vRauKqUo+CPaqkj3uHxmtB78jdXnhGb9xKBxpZj/viHjsnPRcCbhoDEui2UjO
lZC5aPFw7LiPNsbvFduTks7aHLiPN4rEpAEu/MQtPU/34yBfWgoarHQa/vznGlIZTjg/svjpOqH3
PqqPPnmn4k6Q//DRWXSp74j8/Q1TMwUbVkpL8GJ5oqkYRXJ3dwPRvC26rKkInY8eq9GMca8jt3jE
GX9AOqbWeAu/CvYZCc3vA63qIJyfoSj8gdgkVp7st9KF43pGjXDMqOSe7yJre2FRRCGvscXsdll4
Qw6j75pztU+b2PFRUIAjrffJzFPRdkECYX7xawDqkH0V7aGPogJIYdTc2JTBSczF7yUDs3fZH4zp
tPR7qsK9Tz9/xb33xm5zNp1xZnczxPE/LDbf7zT5DwmFABeN5zbzHinzTCa4cgqFWpoPSVtRGvxn
wiPtChxhDRcI0vO5ggvHpM5eaQuH34x+polE9yS7TYPhDVoSKt9rfJbe04n8OzPwdGm24v6adXiN
Roq2LHAoAOpzcwppYti6THZUaZ4eMVKnftyHMfO3vkaAvQERr6xSDFRmZ5iDwWx4PO07phBrsR0h
iBNDn4+BXbaBM78beXgEJyHLX9lvfIoR5Z6mFMZ9joSuAhrJl2QEq2ViPpCdxFWnxOkA/JevInf6
OHVawBTLEsZdS1J2pKY8KB/9yXcpL1U1RfLmbl+DpW9orW6Cr1rxQLSJ6aURPPCXHqH2EZLneE9q
RgPMIZ3oa9z4zS4d0W4lSk2YIzvB3EzxOoKLuEWaf+M7TOOUvMfOwWvVszkIqBpFufHuMkbufbIa
IRRseyx3G3DIcs9KqvuGkzrhoY6kKUSkaVrr0MJsvFs9wdAYgakA/8CcGP57TgnJgiC+4e79al8r
jzwplBvaKiqf5wXoPG8xOsjEwIeHDON1YxyIYfc1/U90qN6gfdzCManBOpGfe5Oxkswh9UqQhPbo
YFjqg0kF1/Ty6+wRIGAE3S2SHd4QzRhrJC5B6dcVfohiibpUidMyNyKEgMnIqeCJJhZNc0MYH8Dz
P6k8t2x0+/NDtMMy2778kzFT7hg2lzo9lvMTjTz2SQyeTYRXeVIPCQzwS7CRZeRZ8eJpaPHKAHQi
FPnkZHbD4PCRVO8bxkgzi/I3C76HMm4wwPIGO21IW6AIAtekTeU0zR0Tb5Ozq5ijS49J+v/HIC/8
GcT0TAkSBNbJt2i6NJX1XeeXg2HaJRFCYQO+lC/YnmrBXXoenoNii4fnRGK1iiuCVf8s9Gixu4Ap
fGtsBU5fsCTl6vpsBzSd/MmAyBGKzl6Camn2saZK1WU8DvUOU1Cj8lh43aySGnQE0x9nRW0CWHe3
x9D27bQ0UAN9X/eT+VbP8pCewfWTHAs1l9NRSWkW8L7fYVN1TwA3Urq5ax5z+uCVQVOS1y/BJGQL
hcLOqYKBTwn2EYUu04xr5PjzO/Z5tiQOTHWNXiN4vfiBNk6Yb5PTf67c3Q/laZtY6+WcmdgV2vIy
FYavw1RdUpu52VHSJJTUAsehxjJaR6BKxFL0BV4TTZP12tYcJl5F9XXgBCOL3fA5bCRhk6enTU81
aaDfcM+/lH3qwQd945phTfMAXZLpdDL5lz2rsnYqGg1qJy6KGuUz9cGxI0/t5o0h3T3xttWVKJtC
ZPAx6io+JdHj80XYp4I01U8vm3xXboAQvXRzq23oB6dBeBr4u/OuCb799r/mq+6GkVTnoteu8CTp
gUcBPplSt32mMqWn4PaXOQaWGphBWaTcFLjxfe0SvJqFoxicM6BkzUoh8EzCsfygVCwrmSZVRJUi
XMFf6fQsl4p66v1N4qv9L4DnqowYTSvHINnI/XCNY6I9mZDUL/TF69gePuShQyijZYZEGBftNLda
ZI7C2gJSQenY2+7b4Sv3tpWGfOgJcvpZDvSMJuUbXGK5/8fkklka9ldoXpV93yTiTZY03yL4TURF
P4Bc0sLc1U30Q4EF9YYH0pSvuAp8Us2leN3nwn53FpJHqtsPwz/fYSMO+ssgh3+EIauVH/gKytH+
qUCsQcfbgAFgSJFDSxEqRfuxItYv806+sk0TOcu4gK+0N92vzra6kV1XK+l9Iie7kZKCJVk0lsYp
D3AbCZUpB+D02OS6kFG35nnFKSKvXMrjXU++UprND6W1J+S1TK7FcO720f7LeaCVMbbGnhIsSzSR
G9mTZCcGO9bUkbesXUuLdF79cr20/95Zjm7kz2eghkia9axnPqYpkWs1odlEBhQcV4OYPxKd0XWi
y0bRTi4gd5psP4QPGVzqzyrPcEg2MsDOaFNJFT/Jm15qHg6Q5ERMyvVZuPex+5SqblKXwEftvQR2
uM1NyKzYZBQDZCX2QtH8CnxyGCpgHm4GszqbhoZae2nDbRK25kcQga30eXPC78WbJcxxhV2zURVA
s1DlbPwyZc/g8XVkhqqecY5n4jJ2v1eERdGbqP56a6Ypno7l1UgyMP6hp1/3MTMW+fwBldQMLxG6
y0JFWxWf4Dbjs/wY4yA1AZ9nW2Hqu7n8W+E7vgAgY9lXwG+qM9x79gd/8PGa6PLXrnrD/N9WFuKU
+nfrytbVjYwUd8rYonD0geuLfM3tSLHpAKhmmVzeML4VeiRt+YvqEpJ1MvxphnIz6/lG6C0rOFXt
VIIJ1x6eLe7NjSOy7cy/k0ZY5ZLlXAK2HV9GEnEBc1KlcHnPhPJtf4Hg2QJ4yk3L2fVOzDW35UMd
jZE4GWuJx/PkCAvKhIY8VcS7bOGqFFfg9pq9mAaWbVlPH+5O9fPMJb8qU7ox03N8xTxzhmozAmAh
QGEj5aOp4RPbvLghcH+M90B3Ny2PDFFpBQjV5mTh7S/15vyVF9mootXmvvZ2w0KCN+ZHt15DOVaK
ItHzFJtg93zFLc8f8saHiUAd6ZiQFMAd5OxzUmmSthujISDcsVK/gqUR5UDXV5/v0SugXxIELKlk
i3j+57qhjk5vzr9CI0qkeeMphfbJCZx3lU0PGk+ANEPciOjPT3Yqk8ErnyMiG+2fLVh2eRP2MHwI
iIogZo78PBu3sETjE7qcIH0FbQKWQqzwaK+Xd0C2RzTfjrDyY5m1/1dxV8oXnB4kLj+YwceKv6ld
B23wrJO/6U/XPKupb+/tTy7cDSq9SUArtAAyMg4xf2rupdlcfD9lrvAxf6EFRzp6YkdQEYk/5t1d
HwmWQyaSzCZTWLTSqII866U6yabct/Z/LZJUPcC+wRt6FosPuv6jYi1oZKI5LY2G0fsPKe7BAEB4
1DuDiEe+NHnfmvc9EOHFLrdTJ+h3/H/Mr0w11jy/nxiICmVOuzxCWd0cb7XYzcQBLEWTIqVrQiFy
lL7bmQOwl8Z1TeXcwUIioKRh+Vl4U57Zvq/B2aLGjxDUpdWmo93nI/qe+OAlKlGYqS3hh0iUUyvf
VJ7SFcATM69ChjdPe/3cB94urmjZiO5Kt7fytDZssHecbzoOcVk9qnYJaPgynWKntynxtASFLFNv
1wavDkSh7Wtq+z1eTY1vIPQDzhkGDLiuNngny8EZszA5A4onvL/Sd816WwihppXHUCFyQHtfQktj
4biDn68gmNGoVKESu7GbyFdYNEOQK/u9Y6W5L/s0nF6k6JUPgOw9RTrBzS1RENH+VDMOWaM19m+1
SITrxFNfqSUisHWEYrj0fJ8qK3UuoouK2rW5+wjto7/SfTZK12G15Mwf5f/J7iyzf1xIEAOB+YMs
ZVMrC3uZF554XRxkQfYXCfpfINRANw7+/VLctvXFMb08ic0JTDr8zStNTUEm2cooVipYjpZnAQKz
w3z07ZRr3qDK9K4JsLFF5c5bA1zOOxly99I6I77vPrgOLfOqXtW+bQUn0MupUqCGw7IgXUEfFize
ZkYmh98LPxD7rLnGv4atUJL5YxfCuWfaN+hRghbmtzyjYGcioJz+wXHHzsOs0lpCs3HJBo1QS70A
2ESCikzKjLcSYGC4l7WIGrCaobQDdsjhSxNl99SxfswexH3qXBASmZUPau7H6vitTPRzrx3Bc1CL
7cTfGZP5tJd8mGi/ktjJnJgRCjkObPtDndUjuStF2lTPG5w6PqJfQSph/LUAg1o27FnJRLAUocNh
R6PfLMcST8CZS+g+9aryxF/1KIb3PK8hx01fiss8u/jKKdA8p9EKBEjLddwT1xO1LLzGU4MEVPkH
dVfeBEnis1UtpglOw1E/JChA/q46/bI7CdijiP9xMrwVxQi1O3sW9d0W9zPErvwUhCTjCJ0kM/9g
/rgimZU+m0iNi1baUW+Bx8KbMeXAGp8ie77TSmKDES7RSZZJvg5nN4yfuqaKD6goK8IlXmmnb8w8
Hjj9RYGghb/uaVH44mn0jjp/+tXjRW+hXXNVCON/gCDu+h6aI+kSaomQqGh+PaEjZWAjbS+NrrKo
7/LnEZiTnuJz+YAJFv0pxLU4FwDvuRFoNLHdiTu/UcIcG+lQU2quxAxMXUWoV9q8urKsP4EwP+wB
EEaN2ixzrAQExiLHHxdd9q0dTixunSrLmxjjvX/yvEJ0sATAGEayf15fylg4Jzc2uaObF9r4HR78
PGIUPVpZ3JNkNSEnKCaeslu9gl86Fug/+noEN42f0chVzp4wG+RVXYZ/BLoEimdqgm50VZUvIgHf
buejR3+aA0kB4Ikq0UaKQUGOrCjjRTNyk+FfyhJYDj+hy+0Je7SmitVVkhEUJC6v2If/SNnmTD78
q0SNviZ6G2Fafb9WVUaSngn462qlD+bZHaVgjR7hInleU7YB3w7VAuRko9cPfQO+afIOZXAZbUNy
9pU0kFlVL1T4sn78ji1jSaV956TKGAsPoQ5veYbXpSDNZl0mkMEvkzVZaptW0yclN0WTPcBdmGWy
I3W71snBRSWrJHnnGEq9Hk8JH8ny2Zx697DP6VH71EXzz+H8VD6p31ikTs/AR2jtQ9dVWAYgZ9q/
/nUQzuo9UHiu3LFS1OtXheLH+0igH9VUOrk7871qlw4EJZ+KqyXUZGUREPJa3j5zHjl1aJZRCX+P
Owg+ZZpziqhdgRFYtaUpy14MNhtpuIc66jVhyD6zoHmM469F133oBmHdoRsiSGustoRwQLK9/Lma
IhOz2t8t4CjVKhhlHZOBrJPSCDQPwuKbcd2xE5n0L8F57MZyjC1qMTjrDNafTdBg/L2Q4wrCchYX
ngncxiqfPUOcs3Eol32XwI59NGzfs4oJZN0S6XLUljT5L6UdU5+HstD6uHVe1Dhw4UTfMBhwBmNt
R5Uo/HPLevx8w0MrQla78wRTdlmueSMyPf6BFEfG3kVCX1MTgDdxU5HSUYnU/NGyWTOc+zX1rNEl
kLWf164fhsL5W9i5h+GCCCgUsidzaYO+gesUONps13Gp0vWYPRvNeN/eZ3vn5eIryJefHD8y8G2U
hn2JY2rVU1RsEQipnH8PeeIjK4x7QCuTfbyJWIdRMlFDlhKcQ50NQcQdm8m218JUdYsZuFrMgriv
VO/rv73hZwpeo7b58g5hpht5/WpP/X77aJcziqOa1hZz0zE6dzvcaIjS65Vj++OuKx5N4zFwbPMk
ua01ci5d51BF9eTvqzfMWFDXoTL1kUmnAtzXdAsUB1T6ZI3+9GBQSeE9DJgAoLd4blbEVFqFmk8Y
uU2r1WshVzYwJv+wlcbYyx3FxowhhRNUt4tVEdIc5vh36fID48RfMAIMMfDBnLJ7IxD8zqqOLdNa
fDlOYyK8OJaG+BzMgCBg/l8/cNNQUC40mzyP9/vj4NVkhz7L8r00XBvYvfltzwFg9jYSSHm3CKH4
d3gkHIYBXgAKvsliUp2/i7I3PQiOzKgUG9TaYL7I2l74EN37wynV2BW0u+2l9X0ALHhDb7l9uACM
yI/6Iqm3B/7I/xwL3InuGxqcgLmHYKLXrRiXQKaKFHgNJ8I3+If2RuCIfjqBxqwjKO5NjPNMnzM0
HXx3d513SPnHbAw9m2+VZYY12LP3JRofbYk2RlVWhhAw/vaOJM78vPBxaSLtDt8pNXZYJC1vDGtw
zk4tF+HblkULW6zyRkFzooHE9cgLEnaFUMdlDGVB2aGTquBTEblnwUtQ7qkp4FE/KhZdHptrEfuI
veA1ftD/0AVwaNstCHNv+v13dvYBsQOX9eAMWZFjtWTLtdyd1oOl+t3D6VmwJ6cxeXkPWWGx3/DQ
N8/+QVN+8FMuCJOEHUI+wd1F5qCIq17IHCn/6ItriPPHnfhDu78sQEtiz5dgLgg6Gi9C1KJFSFzH
R/y1wCYyzBRv0m1+3jIbbJ03EJBeFHciiRzIwcCYLrjpqTTm8NsWUWb7iFIuejeaJVExVkzvIief
HbIA7vTBMGpneVUBYhAYZpaHh/kXh27JLMe/nSX537dxT73cHUjH41byyyZrnGyNl9814J7Hj4uP
TbxbKedMt/HxrHZlrGkq4qDVepb39mxmUx2HsJr8ae3Ico5pLTE5mp0Xxhp45NFh/ntzQMk5/4B2
v7VYjK8iyE9mC0293XTijiaImFYOtcAWZgA+jO/dyttw6r1SGmIfMlWllUdyBxQQCFq8BXxX+lpg
H3WzKgm/NEZNnLwYdRwQ9TVbJmVAISnou23QS1YpSg40HrKuJliJUVwP3jEs4J4sIEcEQi2Rbnm0
FRozBbmX1oQsfTHYJ3TsjMbvgL9NuSsab6ENa/bV0RAxFLhYUs/ax6OW9JYFT1+aCKtobfJY/9+b
apLSnJCmwhfeLpF0qnl7gJ8jxQJjGwJaEI2ecCiIPkhaUKigo3r8X/z/5A0X71Il0ijNbtS96AK3
T9sOJHRQqp4U6G0waMQSciSMUjbmmZuj6Bcjq/eao4lNeLg7zj0L3aer0pGVg7RIL/QYPmmXNz7J
yduEoGU0PM0Zfm859XErthc3brTeExPjoOZ2gPBoeMtVbKbEnl2ADIZ9C+vpFlYedbuu1Nhm3BMd
J80WWxHtSLw0DC87mqJ0tjSOLNUvBMLIIGRJ+JAg7Th0U2EqQQMil2CQc26jcZadaxl3uT/m0Gq+
S2hel6foIfIou7J7DJrml2rnhuID6ZyS1Vg9T8mmXbjmdV39TOl5UMFoxt6zrDS2LqOw1PYQvWr0
vr3Y6bJpiZf289zJJ4BrfPDfDcq3ePHl3oE=
`protect end_protected
