-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HQyHB5qwlNVylYTALJQDl2i5NRe9t2GYW4hhQE14g+R1aDFhGKsoJRIC4bLypAQcnhay/iW56AAS
eiL2lQF6vTYKbtnPYzfj57u2S4C1PFCE2vVu1rIxypyUt/j9X+AG6yAa1kZfp+bxEz8EeZ1zVCIZ
GRWMrl+FtiWLx2eh2iMlXLaRiFhRdHEujo39ElhalL43lsjK2EIS+3ie2T6CW2JSTxVmiKj6WzW2
13Y5WJVYGTFcjyzZKyo2XO8qDsqnEyDq7A7CbiE66jREUYFZhXyQI41DmhNI3WmkAFdN+Bietx9x
vIhe6oTGIB0G8VhAbHNGyv0KLuM612STrqe8Sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
fC0NzwZrvDECXpgVqJUA1krWct1vAktnfy1+ISNQNk8ub1PlEDdiN2DMNTVUiyjJAv3DICmEYahR
eKFc4MzsaThu/gGeK9j2z9QmhOnQWeGz4JfdpaqwTIcJqXQquBAIVFcfSrmx0W66Q2VAolbfNseW
ZsT80LGbT3JdwM23rIe/X+VAYNL1LGX073Vav8Vyc8eSGfk4dUoh8TcBMQwoIomUWMwdb7z4alsD
30R2lZcQYiRqZt7mqh0JmmbCoqc87oipiznM/WPHhSwQhD2ASv+abOJQ+cJwZXARFk1+y1x5KLnF
uKrW/2NjGiDu2E6MjbICPcd/BET99VaQSnb+epeI9P2yqsDkqxWr/G2WwtCMLlCMlS6YPvZFksug
4C6+D0a4jrwk/UfQy4ESBNW1gwpyFk6zpvHD8kV8EHry7LWFaPW7qolsg9hvv7Vj8ePG6ADqW5sw
PatX2PKKnRx2F5Ijq1qynNf5b9LJ8DwsmK7bdT4Z38X3PsgpHutqJqq3ySZePQpLZPe53WiQ1IVA
axAvEf6pC05xHxItOvHGHteohpjazppVQUqOjj5iin9nnmhpDj9qF3HSf4o5Dqkhdp+iCP3wQRoY
w5oTC89SnDt0KzGs/xOHFacMYWVO2l7wIBK0MXaaXarJPH4YxUN/wTXsovL3r8m25CNuVRUAONDk
q0LAWz8H4i4Dq0Zj0fMUFvmKVzrvxFOYqmiR2OM12JkwiSQ/ctuBrgx1xAY0LVysupon+/wihlJM
gMzn2+HhMOBIef7AO+dk4J+R8e3LMgurl3A25y48kyXDQ/ud1+XrVQeR5fpnQfr+RMoGY7kVpkUl
biD/SzbowGPdKLg/7yhNiJX5X5kJ22N4U2Httxa6UIaXPZIciJYQvJqfpNMf/CbWOsHpbUMoXS66
sbZNs/X+K1Q0bO4S+FG93EyYZjwPL+68wggFg7ZZ54gWsPMbf7FUkcHpYR9bpUnImnE14DXnaFIo
BMr+uFCfwI2mYlw1ST5nlT3Xh2ThN6Ch4OZTWgV+RgdHqr8gamhTSJCfunouUGNj4QqQCnY6uh2S
E3Yxk1X8+5RW2GKiYv6LgFmiGuu1raNXtpscLG/k+T4Y0ahaYyubdMK3V5PVULQaL/auArcqwYB8
8BqZ9PdGPuBQv4+5c9C75QblPKKtJafQjYM7xWXZvMY9kn4JumOWBb9SXyKHxtjpnVNf628mOvsN
jJmvIcrPevRF7gnQt0wJf/4x4ZTDV5occ4o1kQiACo/YyzG8nIT8kJ6Xl1r26a98/AgaTf6Y0guv
oP8XdeYwa/K32hFSAQGj6rEZYujehXHIZbm4WWrwJb+JBsd09L+o+3QVyJRjmCiR8WADrGDmQkwD
2Y4g3jko4Jnmi8bhI/u2c75MjyEtgL9r9HbqNsPgqJS13vzEOpVpVae76L7vW1zV0m4Q0Cy6OFst
MfcZCzsKZlCmpUbWdcHJxfHzxPO5k03tmGXpobtExdts15oX85KOPAprZ+1R+FMeQq4wGAYE9ojK
efD0C2u4KBfO3eiMjU4uXIqQTZBWf2ZCsXVfatVsuOYVflF2tJiYxTZI8mluBELUfc+sxrElIKfa
a8o4zyYsO58lYMfdILbzXrd0mlE/mR/BW9HPyBBJjKZ6yF3ojctDtlRjtWdnPnUkp0gvZzwbxgrj
lw4C/xpnuQZ8rxrQaMki3+iVhuxQvrPNPfQ6jV5yfh4DKcDWFp090KdLa4Q3l3Yp+fSWQ8VsY0f+
Zqk7xlUQ1p0AMUZ1ps0cJ37Pdmi9d8cM06E7YCCMBJgfkVY5UXaAU4LMWKwzbVfkDZyqdZG7UUwk
8LGKE5I6rlYObNaxcpykJ5UZDlHGp02swW91kxXZbo2pdvcLYYkFYSWI2CRbyeb7K/bgOcb1KiHU
jQFVWKmLswOChPLlh8fVadF8yWhZSYFUTfBkF9qzCQ6W65fseUCm2o40pfNzvEb8zOzxhSvMuUsC
R+zyitaheg9/AWIZsbG+QkXgjYkiqjTtOMiz9em/+gJmksw8YNZu1eKEtW+Uy1pl5uwgehIZxxds
dKNzw0dBJgGzcp+UwWsWjmjdIrkbTRvDPB6tAhSPmI+J3R3FRUJ3kh8AOh9AzshSaGjaEGsR8JHL
WaqPnwcGgFNV3bdkkPEJjuBJQdCkBfUUVQPKnFGvpDaphaQ8DZfut2yYA8WAlHdVV8AUjAMe9xZM
Tia6k3RIMTQANcFmS9G13AYiRqlS37jNRI4JVVX16MhuqrI8zMi6yMRs2xVTbRWAWpJcjSkTSN5S
yTascz5HFhVXHgxU4rcNEkvVQIMMX1ZR4KezbZhgpJgm80zknVKVMh4AQwrVt/dWBpEWTTECcq+H
HQf6fRz3bua0Z2upbq2j018aLuLTVkUjg+7BKTcm7Bkkmq6PyR4FwZ31GtpGo5umnuy7UlwZjvn0
GMlc0WCA6XiBeoUtU5EuxNRiILLpL/KExLYW9JmULzBXvs7x5hsWZDiFUaj4XN39ci/SxGPulAnp
3AqDmk6VAdCTSmcv1J4l06PuJUmVMwW4ymAzhpZI2bIELLPUTvIc97XJ7kmnivygoPidPJyDMXMK
l7VGW8SEJBhuOhXPcnxKBPwpN0a0ud7lNZ/BokGms+sKMzXoqEJ7U1xHIts/ZzXKAj45m2M1OS6e
EaI/81CLY3uIsVmRHVHmzSPrs6rj0moMAKE++Pi+OROQZ4fyTs+3LMgdZrVeFcrRtepo15z09a3w
eapYe+Qy9h06ZEkCo7kPrsPFKkVZUm8QrFhEcbH7++u3R4uGHT0f20Slf9keaV6oHJFwGQtEYZn9
I90c3poLN81huA0v6HQB5DoEsrOa5boj8bumWUxSXQKRWJo86mkvzujIgHCUasZmYA+qJPSFM9VB
F8/QvkJjUXgOazGDi9R0EclDtkRk3cYRDbDJrdsL2pT0jtwDxzlSwlyLN0UAktCOeZgxx4oEOPuy
WGcFfqUX/wcXEFLImcDct4lLnLBBPWR34NdzFWiUcFoR7exHGuzjrxuFURvo2g3TqHvkDrhNQJWg
3HlSBOIqNWypdqQ/PYGjoMo8sZj/pbyOp8WqhIfw22TK2AG/e+mINRtXfDpd6BI+i5+g50UaOXxX
jnje2/bURmHLmruJlXD4UqBqSV+C8hNHX5ALZ6NCpIkVpEjGdIf+7xiN3suO6DXNdWc6ro/YbVqo
SyYIcN4goF4UDV8tSW+av+nKuEQlg1BLACWLM3pgMh+Uyq+9M/gsTARjjnfonGfTaJrvflbkcGZG
8vTOAbfVI9t33dBegX8umpT6sOIcbvnouKqJM8UaapZiBeo6MqW4fqj5t47FCCrNhrtQU46hZxuV
NKGXmAXlFP2hyJHkFGjFUZq5E6NNA1sDtHL9Qm8UyzQwLGM72JbP/ged6unXw/h18CVo0lpBYTaP
qk3xh2taBcZAeN/FB8DrtiiLzCkRwG7gRIkhPmjJid75iww7GRMJTJUTaPN6dy4eYn9yS02Glvuz
RSaIcb7GbY+7KNDJtEcdh9NE0YY4ZWOdkRJ7Wv4iVFgr2lpQ2C4C5SpTETbUJu5TGM6noCEr4L/P
CiHYwXOW3kiShm2S2YAB0dmNgQ8p7IQNf5a7y2AO6kgKHwTg/hJ7+S0YCkzhzoIcfrCgpYHKmzc7
+s5Ili2gWg7BnDAl7PLI9TLeMOZTIizJHM5J4i3FctQ1h24gDorTQhm5oDt4zKDDI7T10iXtXgcZ
5xrNknuZ4S5vQJqrR5hrEu3qgqTtM5BnoGHxE5nI3WSWGttgLAGzLOiViP1jTHvPuY4/BLHv+gCv
LF0J7nYpkr1jI0pX38Oe6yEPaX4nlpci86AMNSzDVLRYhR17z+D2N+TR868ziWAMDlbNsWn4RVhC
jxReybQOZs9Bv0NW8aN6c37H3C3YMva+kqB1jjFrPfOBEqNxdN3Ou7TJcvoh2WEiUB3IZrpPlEZ1
AEbi9x+m7pmYWfgu9BYdFlxK8ToXHVdrMSpu15eUu1Y2j/Fo4IQYaxycuHB1xNw/WKTNtPayKDCP
iseEsiefobJuuWmRsZcgIhOJmqRvP7DRFIWiAE7rl+6Mol4NSD2T41WP13nCbRF3ziNMIlAzsnxi
4mXeebbVcPgJx8pCc4NYd+hTNy/DOQJW7JnwiCYeur6kavEsklQXTQkyo6UXeocqc4BfkfjZgH93
ToE1cOgIwzQd8YgOjKrG/uJXukcAzbeSMln9rGtQe/V+VdBVflOJfnuUIPwgA2q2HPXCiTmlTUH9
8zjlPRNOpNTJbYrB8DDaqcP4wLFzUjxrflsZAKA5x2ggu2okiJUqlsg3AbkXaLSDEdEuI1mpcG94
/Y7+w+XqQm9Z06USMr0jYni5O4V1ZbcRHKjNwPpKreg3gp1vQNHB01xnHZBjoEk53BqecOxL1vBZ
Qj6YpRK5b+in4l4PZ7PW3pGhIu5+c7TGHUXBVHWiSSSaUYO2/595VbFdQc+RFpyHDA/Uv94EnhTB
aerK//fN53babByh0jsaOYMouPQ1rpPrhal/3OgAyu1/Kn0Z06bDbcRkAhbkwLSnZbL1WDBfZEOn
tFTutW3C6owLnO/kE5t+H8ZkrBC7DXVSXGWKNo71Gf/gZTJ68bVX+oOrW5gW5ftha+KsyxJHyhss
AdFihCjV1hffwxIbV77Lskaz9V6rRibYR00RPBrwIhuDur0zVEwRGByD/IHxzlBuzRYj6Y9ZBXFC
MUUnjHmpr1uV1yzhOUPSF9yOVBWUzDSF5AV8MfagURCnB/4w60Y0C0XRu4/rQ0EkRxAXtIP7IZxm
6xz4FwJFu3bVQgCOi0QatmTi30YIA0pLiZmEO3QjwH7RufaG28FOnb8FI9iffExAfEuLMxvLq3od
VDA1tVDQd6LvgCpAC0McZmZ06KIppG46Cc1ZLe0Fb6X5zCXhq1E+jN2nyfLY86T+NR1MLtzF9U2/
JcQGMZUNkR5SAmiCzQRfjbuLnMPmdMehU0p7c0Q84yw3Eg99Hwz9nQ2fAJVvchk9iYrhCn5eLADy
+NonEzTdoBq9QWuVL6N+F+YvjBAEAtzA9L8vCLST09i2LDkC4eqLlSUAUuYhuZfkChmIJlBMzbxT
xoBrExQ51h7bYqlu2GILgC2PH0zHHvhfc32oGoHHThc1wHZnK3hHlLx72c9UnYGTCOAdj4Fokpxa
yqhv6k6nRniduGC5nQZTr8P+ZO2UCiuC56oq/SV5+b5tMVMiCa+tMAV5hWoG+9pLy7fz00m+NAx2
hXw0SbYZT56sSi/3i5eyU7zxb8v4i8YI0lrzOfjGoi17gkvMPP7rUUp7SjMSgWbBbRjDHFFkDw/V
egWrp1oVrj6DasnFp+ynw5yb97U3YOyg/n75Bhwvg5qYnrjTVrsIQZRbYRT0yauF9VZ2RFs8zEpo
fJEnZx1H3cP4IkXR08ZHsnz7fPVnGF3K0assuwP+lmkAzpUHYus2s008AZpA4URQBIpYnFPp5QN8
MXA6OMlWY78145rYvweJO7G6Dw+Sh7HfZS50tpulOECq0YUKL58ecIO73+QNiR2c3hWfDtuUQrA2
aMq740NzU/9bWJsTaQX5KCOIWVPOek0GG8X5Hii13bUvuPqsy72tSjVT/7BpdzQjQVo7DlGftlwD
gnN+2NwtXn5t0oTxmKKvWhpYGZi7DqWPXyRaXA3xez9kIt9ypwFYHxFgkGlDfGY6zr78LeMMJvN3
6LhDeC5Uz78ZZSNv0sRUmBIelm++93Rc6mpgQxZ5FMS/H/Tuo5zfwu85jEHt9CnlwrTzqBzWVBQq
IINeM/RX1U8Z+bdoCn2cBj0lTmRJ+1RsfOIwyFIk+OrV71hiTCY/N4xXkJ9JxKfdr8zvNLKv60TV
qflNfBrZe0R83OODxZCxoGukdjndBqv6YPGETNEJlFyZxTT8eU8Kw28o9i4XxzlmHiYlWnFZD4AR
pV/Lng6cClj+YYhtgzJMq09B/4MpvO0BvNvKBmOAlkJaAR1FyU/TyG7pa2lQRrBfK/nNZmK1uxwX
HwY5rP02EW2QD1QKX1pbRDiND/xyP3z1cd593l+lN7EAaMah9wcjPBRQh1lonmdpzt/j8nJb9h1q
pzh3Nj4so1jLOndTUOTEtE2Xf/xuWTW17Y65f5MwYaB6y3L3Fhk6xO5SdZQCQqc1+wqMhaminwOV
c1wlVLiE1nLUBhL6r9+KMgWSlAg4KIM+ybOXj3KBc3yYT8wtc2yGUZ2841USf8wPovwNBT6tG6Td
u7Mjpog0WKps++W7sWwzolvpDpH+v59bJgYIhyn7ucNFklbKd+KCFXHJQxE+8KMF4sS7cBUE0pUF
bC2VPasRx79Lot6nSGrwv+koKJy/ctY7wy+Y3ncYU3qGPrV8bSoqAMfxqKKKC2ZGTdH8IVXXw41Q
Jif3t4ldLxUkOPxFTJMpMQfr1ZNIvEyg/C3Eis8J13ZT7iHBg/svBU2Ytk1+nz0WOAjljJuS00aH
46/pGZ0KOHcu1SUL5AmOyJBC0+HzwQEcuAGWjdLF7UQ+QCh1kiaTUpheCiii135+qMXs8lspBqRA
xGnz1A26eXh00swJj3F826wnWFf2cWR26cA43XAsTtJGmMnv7PHIER5KtIihFOYTW/j6s/1yxshS
37zAvAOu7tE/aukMyw1QwDfyyq2214A9+o+V8pkfN6tCq07d+bwffmTX/CCRLYJdqlrNQu3YhZG9
b79K2kCrTSxNcyRSf5UBrNp7mcdf70lX1RuHBnQ2uHxPQqy6ff/uIzZokzRNRGP95OV6vgF2G84i
FS6OXZ5l3lhTrbc/LEhls0wS1/K4o12htoDO+jlTXJHFqqbY/MlS8hv4aJNXpROncypcEEPQW2Pd
NRcKpaQNtfVudt0MPzUhWicpvJ2K/jpF6F9gOysqVhvRBwn8I3EkB4lQaSVx6noYTTIWajlnv5Lj
MHPlWvuFpn1WsI5EfCUnO5gLS398z8Xn0IhwTy8ZWpML2v2QbGPrJlryxMD57+ylkw9ztIUnes2X
BTJeWTsX7l0mNWqCgPM6h8c4lbvygvrbjdwfcA368kKr4sf2CzgmuXah4g/O0DbqajwQFusH0dXs
DJ2KZ+U99zWnYf75hqZulT2wJAdAuiOKZzw7B1yvGZOM6You2+57pFO/s6HxHdwjrm54p5U5az15
8Tbd8ydRABeGYc+U8no3F8Pb7uswUlKfRPBGV9rTJ9n6rw5FGvwnmA1plFmD2nN8MFlMgnd1SeH9
AK1mmwbVWwxWRRfwHcnWLNookfO4Iv11lw9dVAz81f4UCFjFKArplaaXhDN7GjERuVVMRanFINou
RuU7wynVJU0kK7q5NnQcwEmZBBrD+nsD8Iytga4o+qAX5mINToEkdTrnPI5KFaS/ck7VxHz6vVbL
a1DPorigi6RP3dooLhJaknGk8ktgk0erH33AF4pxn1EN6wuMbqhMWqO7eHzZHZ1YMxu9zwaWUlty
56Dn6wVbzVd1fvgsvvuGCYq8odZLZfutA07/Zx+ZNi6skYaznrfvjptvO+U3TaS3ZYNZ8ap9/C/1
W2SxYWrWeXrCYs/uHhkdSIYYJUhUY7XKef9xvSiwul0Sd04zBQIJL3uHeePaYFd1P0q3vunD6/xV
pYCTyzmXfk4XB78TM1A5x5fp3iQROO9aVjs9Aqv5seNkFQWDJPyfLkWng0yDPO/+96JrHuDMXJQO
dNs6xGyGgKcOCz6ZXOYyNL1yqtPdh2N8b9Zg389xJQn6UufXpJIOnGYPK46pmlQsjTJiscKnRIff
SZrfhfZGJBDnnXo9PnYBY723vRSN0wppG0QogOVLHBT5MSkd42vDbezWGDIXjvQRWNWTYvcYZcqS
tRFQXwhwlRn4TcSmHTMVCy2ohHgJgDm8coHIn1u+tzIIbGCtJX5wvMXc+sUGL3erwva1arWJLXWt
1O5pboRA34OSW1USFSOAotC6IdI8tJ627kesr1e8PPoIGS9SddLZontINkq5GA/1BgkiXKKUfD4h
iDBLdK0OWDlr0C2zOfE9Ebnfl1TuWbqswSLrVPfsFFCkMSPAoU3tjb28xedQ/Sn+rr4wtdd4BLim
pJpBAv42QKyariz62VjDwebP0QSIUCpo5EeU/tR7IAt2nVr+L3ypqsfbMpEmSNxUCGNn2PARCv5I
AK9VBLurFjeehHVDOekp3kd+R/5KXjnUuIrjUOE78XNtyec0r68yLTniD29bPPCNZDddJrLw62Xw
fphzMuucC2KWdpzrV2olz4X37TccPxhQtGo2+XFE7tLAhgHpzzJ6+glwEgWx5F/LcgpExp168tK+
kC1jXVOFesACE1E2yK8xGks2BrzdfB7AzQPEOoPItzfgdbm0tL0NTjEhV2WFdhkdWLxp2igFwVK7
FCh8//H/RqCroRPZXt9ArvJZOUlASldn9QSMiK6vmgg3d2SXfpsK+ORzg0R6oDu99rC56tGAUIiz
bexarnWn/TAjqYgqHM06+e8I3vjOpxKiQczWrcn3xvrvMuegApijzZ+ErEZLOrtnu7ECPezIQKJ8
eHK4YYE0METXuaap53413Uz/HAr1Ma7ZInecEdStPEBdWW2LjRez6e2ADAetZinX2jcm46zHNDNC
p2o8fBvK2DpI1v5CF7CEJe3lps5NxxJStxKkgANGacQpwwhhwNmk3n6CN4sl+jY43FF0yk7xqo3b
pyu3RDRxW5phen3Q0Cwh0GiOUne0Wl7Is7Bj8po1VfJnFU6qjMLYaUoGRx0W/B6J130UFg/wEda1
Gj3hMrVUfP2QX78oz4ZxWXZOqGSNtP7VJf2MMRmHQdsZmvNfFkVZaYqyqlEHYMBd0/4hHUxlGBlj
NNhqWPn3qybNUMAS/cPKp3X6dDcZolrRrAaYS6pYTvgTUwa/rHbpNKM24Ivb3OpwGjensQWqgzVo
iC2kJzSSYXZ0ILtjEGlBvMxeY2JkjQ/2SOHR9cBDyKdB16CG3jSarxqZtvAS9bmQplSBpdVvcE+o
yDvQQ9mRTm/0HZXLpQTLIA7cFDoZH8oo4yOPv6uO6UuDaMq7OBWL83McWxxk+ba0sCZmNQZ7bKpK
soLfqbI6H5F1rzOeInSdpslomf7Fh6h08dC0WAPmflEX7snhCLefAIs8K9khsmHXCXQ1VlPah+2J
RzM41KpQP3+Ln2L5+tZaS9wOMZcn0eQlc10EyztcZ/Qvm2c0VsNmlKp9tvBf2CpWEJVKwzkCsJBj
dw1PN0UI2sEUs4SLIdy2aUmavBR4LdVPzpmPbbAKEV73eEbuXrLtZiFfjSAM4AatNd4duwRHRrif
eJIiEhwkwbQizXW+jyC9TaXHVVjdUwUPa668nJ0HL7uoYSA2Ay789doxP70cKkOGRxxvAUIN70nW
a7BW39Xt+ctgHn9lKqmb2iojJ08Ft3HcuNmXXFdGYsbdaslC/NCkvv+u3qS35lgjgR0ZoWGEW/zL
XDoZuNu4altanW1YFzKpzU1+HJ9pPfrrwoRiTl8D2W/GoyznLl6CEK1QAmmOZliksnZATS/xAm/X
Riyg+Tb6yuDq+adrR0EZn7XhevEUs8cw6QIHXl0p+aOhD6GsCQRYgar/l9dWUm17cmDFKOjuh7Gv
LPlKjdwZVKsrCblJ1k7AeA6/g42KyT0LvsoZjHZqH1uEqauBrjg35kp3lakSE1SmYnrU3jXDBn/h
SCk62e6FX30/OuI7VMt0mvBUIu1joasLrD7Rk1D1x8BAoyxMkOpT8kVY2eRwwUayl2YoQBE6QBX9
4tWCmZXno17S09zxVqcPm9AKk5GXApV0LHS/iSWkbp4cgD4nYbgaTOHtX6u2y7W20cn9e6dJBdVi
low1ninBM2TtIgwgQxkcFxi2YSW01Npi1PecQP6yg+u0+Er4C7QWeHEx73pkF/DmZcInI49rfEvt
IJECDExaXUa3uy/iQ900hSnp69vAijgZTh6jtvY1sRMSxPxPYDuKjPBbE/Z9jgOPxZdUMbmTIb1N
p7jgJ1FaxPm9R3qBuNHyAqWuaQWz8G587SMmv+KfBuGoDG6mz8BThcZVNFkG911L05gTqSsAOpvx
kuNXSCznBRTyeFRAbAAcdfgWV0FtoSsq0jm/CJfiVCyMEGBH/8qF3duJkfZfzsyafqu4hveVzDou
RFhJ3JazlHyYTDP0mxyouy+WR4KwXHgEc8xnUNd+CZmVBHl9TDPdR3CQt8+otawXC1k0dq8qiiqc
sf0l40rOmfNcv8tZGfLWg9VqRz6QucXw7chKuMxo8QKAA9EtWR6SgxZvIEJNK+zCy+w1DcxGWLEU
Dy7Yp2rZR0fWF8MVyw1Yj6sgfU4Ow/RcuW3B7GDZ4oFWMNIpm09tg2e8QJpraUIkDvUk4Y6OHLrR
MmRI92tkt6+09KHgfQyT/gQAA8WqDI6+SNRRP+OSoKqnoQ/83tC9pPAUup6Yv6VVsWgb+cVSPhTs
0W/bglTX0SCYa5qfpdP3Xmy/P8NUnfJm1/bCG8H+nFnkF+fkSfkC25c8zQr/aFeVeVjyBS39vjjj
APSXMWuGBUUyyH41lRFnppOGFualRQfXY7kOoawmKogfzR4LWEu7xARI9n9BVM9fyWPKm9MhErIl
KcGeu1yX3ZHT6jjytwlX2eHQOIdjcMP4CG9mdQs2yfoWk2GNPQBis3CydNs1FaefV1EAYUbw499S
LFt6b1LZQ3MXO29LpeijbhsI7p36jydNTLf00Sxf8g5OKHNlEIEvDcgXCHPVrpJr5MygPGJyrfsx
Em1bJIpyvoSM0+qkdlsBOvS7fV/QnCtCx+Rj6QQB68Fb6IpFrFFWwEQeidq7xGk1yBuNg7uR9eYC
7Xc79QLC+abcAfSZN3FHSax+vSPPPShZ6JauxSLjjCRTh37D8OCExkMofTFc29CVSphaSSQQflEX
Tlo5ZLm6uiWpNk6I/iySAdUzSRnQa4lX0mJDi1eXvAvTNuFdB2y+beypRW5eTXABlTRMwY9bBujc
buD03B4pZfli4L3jEx/bT8UQ+l/yKSqA8hfDXQ3Z9OQbxkyf+epFZwuWNLiHbiBFsZb9rhkcWpqL
AuXDeluGVuTXeKgwj1pPpMWWTbvCePYpZyhcjqzJPSwr7sEbmItw6vub7kJIkILDZMSNxRdGuikO
wdHpGVr9CTC5dTX9xP2+OGlCAupXB2noc/0isrGm469gL/TgWh0vGLjOadCvCQx0gbjYbio42rMM
jBBZFDytqHO+v17sWpLQZNE8dL4NOYUU99LVUhnxDfqXo5J0nYALoeTg+2BePlM0kSlLlOg/hIgU
in6QPP6syT92PqefG1OO4HhpLqHzGLm6Q8FQMM19YsILSomEBWVj+q7fcEa8ROp8Symqy8pr8Zd7
mD2Qz7Bln0sBP9yUOlgf1mdTpIdjxybuFdYW1GefzVEcC6vGl4wSJd2pQ+pk1TuIp0C+HGXlm2hV
LZOePnbeXQrspDX3JLMmbXheKtTcfp5TaGeH9vWprFfGpcEjRd/5O1VBzXUOTQE19YHQa4cVM7Hv
PVOncPJTQBkT/WcsRJiSGN9/IRuEJ6T4VgilmgVOFg3iGJ3i3ETHSwV4nFfMyv/ldr+pb+NfZStP
mF7518bfTDjwJEsAxC4gQOlgi8LNH+kYmpnpAptpCVBG0ddAt6T+eJfGq+7LAUVdBPSUxqrKUV/5
ysVreWv08h4+10BHZGWSDN+iCxMUGj6JkN+1JWHlSJTNuYWnksjdRnV6ThIZV8a+pcfzYZehp+wz
TLtvUluZVpGNeks9VjCmjw8yUhpCrJ034+q7aSrp6IvaizSIZ9ubizjbaA5JLEfLSMxQzTO6r7Fi
9tnTpsDHFUKVVdjFRjWsvvfbxy+oFzCYJUPJhntRHbMBtsz73xTBl1M6SJQpQuJxEVV8MgefZk60
B45vJGDYswkx190ptnFea9aRBw2Z7OFjKzOWiT7HzpO3zIh3XB9iJZEpTAnVEdzoufg5xufq43LZ
OWcwSc61Wb6O3VgOVUImlBmaD1WtfHu76gtUxpbFta1oozA6kgC+7gUsVpkYxOxt/Rx9UonXQ+mQ
QJaJpsXfigxm6ouNW8e5Vo4zYDvHbbMhosOFVPuglLJCZ6D4z/T3Hk1P/4LsiN34wP5evyPSmn/R
Otxo7J3k/GUx2nEJyQC8q0I5W4mDIDkhvZehtOjwZR87HOzBo/65X8uMZtrKNIg1eKK45swasD+9
sD1gSRtCa3Li2hWBSh71qGI7+vdI/LPPJ0biKD8Zx+2HvkVJNaK/4Y9kTKtYJpBLYJe3xFL84bwM
HmltIf4w7NKQx86yT2dDvJx8KuucQawpqW9Z5/O+VUKawnd2nSEqcCtfkqfmI6Kjr81lQldrG6gc
fRLCBdyw/J9uZAQ9XPtwbWIapV0eydJheosZsWtfklgiM3UJE5h29VdvWQTPD8aXnxN8vEw59qHO
Muhji6KFVRO2Z8UvAdNqA5bW5KLTuR2S7P/A6g7wCGh7TyI07YP3BXTt8ZXHlKaXsIg0ke8XyXBm
aw30Kbi+6nNm8gMq00kOSdOkIqJ1izEkcPXt8OPuu1Huce1kxJp+V9NQRYwqrXzi6p7Ejp92NUxI
Hdm8BCjRMOjvQuiF+T2ltDFhlPOE52rm39Undq6ju4VtUy7cy8T1OAckbj9QJ7/dyyPU0c/wwCQ3
RbuCBk8B40aqXwPmC+4CkdLhOrGh2QtXXMcUXVF4RP017pj/bNaBc54EsS33KvXjLkpy5b5uaTDH
xdoT/9JBW0ewkC35wxNN20sImLe2AsV8YJgjk066bj5Czvg/M0XEv4+zRk0qCP98AQQ+q//ITsC2
WgGWj6e8S6pW81Zm0/TWpcoSvT1JHvJ4QcqJeOy1i0gfFYZAQwrVoek4HAPNzZ2AQu0PtdsaYB1q
lOU2CqjbQ9Za6qamV5sC1JuE+CjYjZEGr2CbO7wPUwOrUcDyoMthiXh6UVs8uiZS1Vy7NXMBeHt5
b6vWBQ2/rm4+F6uUiTZQ3KmKYjRpaMKLt+nuyC0vln1d7rfhjDUEQmzM2or5bcIwAWveS5RxXbCu
0dgX7w0IEToxvrJAPzmmCgz4GPi4/lUe9wHp2KF1eY/9BHQVNeZ+Skumg5QNfIVeNrOg1QbWMPiG
d8ERd5x+vFNDWQoGhuvrlQpoNKCiCa+QA8owZ2IroADPbEl1YUkni0tIrdF9GwWd0CATEpWo0Bb0
/r/xbTlIkwmyP1Rnt+aKGwcIzzKH7RgWE/xU8R2RBwoNVGGdbqMT5hxo7nRVPO627a8vwo9qDu14
CCQNoEnaKXItET9rWxPgTUbrzqKeiJ6z23KMP52RlbTauq7YMGeZ4PwZYv97C+gvEQv6jklrqeSB
715FFtEPzN5drbWlU8N9G1nK767scMq8yzUk3RkBCIcbLRJjANuJfkPcXJ0qEte7I7xD9j+ckhE+
wOXj0Ouy++05gjvxDztk26FXzz9mO6E50RoztdtXNk2CiSWyA97KTEEW4rvKtG5mv6CcM92IckZS
xu0gJ40mklu14N8pIyJ8Lo+tTeA1x7c7WR445TSLzthII3OVrsqqVlPEytxQEr44J7rKbYn8GH0q
ebg2LCGOyRW18DwmftE+rccz+AXZ6GR1T0iOttKQ+9pfFoVAcn8hmVqwjUgchm1aDtDCSc/Q3sql
r5pgIuzsHa9RCiC+lV0y/bavc7C0V2QzQcYZamrDNf/A4jQih0BW2VQ/PSaF3ZXHKSEZC0ouIbBd
QQeEOW0euclvJl8KV6GBCdb9uwYpW5OZeolLEPuT4bEtJECKEhPldgkrv1WxyXGXQFRHZUtl3GIP
8IGANW1zWoZapr1e0zhRqUZOMu1t/IavZnfkFoBXmHOoma2Onq5OLMxjdGQCIzyyWF9PHrb83Sl6
lHqZ1EWuFZm1f3q4ta6YspgyEhLjZ5aA30WanaC5cQiyMVBjTfno0FMZ28vkZBwh80hUt8FkqqKL
b4bWrLsEbwZFRvezD59bjAaNaH/gWuLj2lIGgx3HH4i947YmBEyIC+bDoYLIO4Kn65gm+99T7vpv
WZUd0xxZDVeDJW9QL2XBf5cPsMXCee4z7e+RvdBRd2I03dwY+jXCk0X2c8glNgYLXUP0PrdKa6S0
wuJSQfAwE8vuhPJZj94wFUHXbThXXN9b8UJeE/ygrXTGcDpVcYsMMON3px+C+jrVzeLw4+1PBKu4
zA4P1XzlYVCKjxW+20UM2rFwar0TuFdFEjFEXiy5Y5vKstsBTt51UsXQ062pqPaVlaru5Oq4L0Cp
1JQruiRzBV7RZZ135cavVUZInGqCagQFrogsqGZ5Ly9r5+jt1TBGqaTlyLDg2AfxQ+2PqaZtmemi
jbU4u34QRZAPjxy+6TZ95/lKEuF/4LYDfDDMW/kdSLM36bpK8Nw+qqc1SLeo8wypc2OpUwiTQBld
/5+EeaZvuRnQMwqN/Zn2wolMmFvPaLUeuwWSseT2FsR6qwh+ku6hwJk1w2eIiyW/kPVpH0YLJos6
A7lZvB/S29MpYRnclmOtzruQL0Tj8aSKprBaSYHWyERYBcQ54PrAKit9HP4syj4+Sslva8+yGLc2
fn+a0l5ZYOGjk+/EL7QUlwvbqZHw066EM5h+cAW9FmvL2VWXdAZ1t9kUv9SwGPfayQBYsnUEt91m
c2cOVMtltMnCIoiDKfTyeAodhZ36R2S4nBdJiTIV43EVdkHUxLY7i6tfrYlRwkHHDtMUZnq877w7
jyLDvQEp3ruPsyIRKXWv74myOYjN3AAqxWQgqK7r2uyd3QZNTo2abM4XYBDTI8m3WfziRztuagMA
I/mYH4mPEJwBNqLYwp8apnPw0LtFfHzEtI+vCqHQBK0zAlAFKkGBhZjzsGl17U4UzIxZsLJxLX/K
/uUPwmTXFIxGiQDrXvKUAY+dcidrJ9KYRqAPE4gGGVBjFZnbGxxxQaYfVH5gAEE/ar+owbBHempu
93JYx1hrALB6Ba7fs84M18Db0xT6oLxKuIrqfi7+6HhPTAWbBVaYSXlaY0U5wfTlObCE6tp1BLJ+
WSZ/O0/im0o0NlwvvXPXndZHKruEmqFY9g51h9Wm5joAWf/oEz5hKH2BbQbTg4Hu+t79T8mOOZCg
xdqutF7u1KW/BHA+q1rT5dLfWg8sduYFHs03xRMkL60h6yaj9vq2az9+eDQBPjEsM1gBRRTDscWr
6f4U/hHrJirIzHya1SQ7ZKm+50HbIPgrngIrHg5qcJYKA0mva529LPReg4PD3i4N9QYk12GeqSxG
gm/ZhYERdd8zimZPud2E9x+9K+tAOsu8EF+ByVDyuuhf1M9xpuU+kB/67EwTfSOYPA8Xp5PFTR1D
6wtfrpXks6I2UtmBW6A4PxS0cPAA814c7sf7N0On6WOZmHFzqcyPiCzhrCrkWj0I9olh7cagCQlC
YfELQk2eSW5U1/ciL2k9w1gMSYQr3y9ErWzICUSdY/B+n+IIGthLnwyPICtKQhDZeSND8+r1g8Oc
FLxO1RNqAQRp0vMFN9eW3AT059LnhTkk3m0IfbDDEzAztzpTH6h1515b+7c0ufvFVzkYbmrqTx3q
waYBEnro/SAQYTG2eLgh1dBDWNAkl3vHXA59968WC69cLdsgfoJWHK2BlPfBhRyB5GLxca8Ge62a
AMcP8r6pwd3mKOPsyfABg8+YmUxkyIQn+WX1ynwK7F9lFpEyuGv23vUzCy0InXsW2P1FK8D1YMmy
55EDCiO7uBm+Y6sYGHLAUy0lUNegrVRvpHdeEe0JoMl0ODExzhBYC5dyawphhV6XVP5hL3d/nchF
CItiyIch3UKR43jfi2ELoebCaGYnKzO/Yi/nk6LW1XqH/nD+z7RthukY3/XhyA2yqvwWpQnVscWy
rlK7I7+ZNMkY4/pFU52mgL/G+U9fF4faSE+DvmbZTvS4G49bfxTC6vJmqF7wi3kt9tyvTdWC3ca+
Zr4qPEnxYtCGpzdWx1TIln7E0Rqvk3kPt0Jv4kHPBfHqUzVAs0fm+jOXk+noKzY4Sgp9TeUKa9Il
Hb5jho0+hzVRooDkk9uFc1GQfSqUvgPH0S2yrhwSYwmkz5GdBNj4zZA8MTklE7Fgwfcq3zVX8ipl
cOii4J0ElPEfrGJ+BMu3RwaDqCbeNX8xQPQhGd1ajJk3UEpdC0OSRRtwaJydl1JYshvagdKd/mCz
U0h5RzWZKKuQbtfvvRp9+7BX7fg0U93i7drButU6xyNjQjzQm5uVqplott+9xqDwWUgQsaKGsrB/
DnuJlwmiO7Pq24M7Hg9AaDzv1Sota051C3x/zDtU+VjpU67SfZ2ELycgv3v2Y9OrgWA2Ct4Oy4aQ
aK2KI/QV0vopmvlS3HC7bjzv8EkFXkX0j0l3nITvWTLk2mjUsSPBraLo4EvCRyzxA7SyNcAn+mt6
JC7kwGgf5QN3AjOXWVOeYDcaOCcr+UoByAj/ryVANdVND9aeMtrW17qfh9jCiNL915+Ix4V4HgGD
J8BsMoQZU+dGA06FhOjYwTyEdmTYi5fnmvmjxigdxpXjUJOegHQy8DXBh7p+SVJ7Go7Ul0sDsWOa
ah64ScrxUT6BHr+G4LdJT/92OB3wksZC4XPK+efNkebm9IAFELwicn9jtZOw4Sjhj831ZLjHCeSI
pO3Hti7AqQScUVnGqiZ8P9FcI1NiahrS99k9fH+CEguhxhRPCKQpJ/ZvOzshEOYE1rewh84MYMA8
EPj05jIXxI4Vky4JBUlwFW21BL4sDKTyKVX4bk5IefsYt9kdvzM/18x/bJUrfQlO6LSkUZorlVUt
ZizThkFchC4BjoCZstwAs6zXv8Y5Nplf8vMxAZVBM7UKKUXgy/WcyRz1P2yCBa5CeMZs65lRd8KU
/DWd5LwXfoH7F+Z02wVl3aB95WFD93f3m6Y4ghe0OPPEbQmJ3SGT7FmlRs+9OBUajD1bV/W5QC1q
Sc//0Xh1yzB32L/qHl+AWhOKeLI5aVO6GG2sVUzlkSDLrvESiGNX5UdVyClLqc5BlMY85n1oIgnJ
PsxatLv3rQudW59DtkXD1obdjuuPB7pW7vqPw8SoalXgF/n4jkqvFWROE2leFIi/W8e2qeSmjqMI
1foglQ8PfNwCLdIZanvBWF29odMTKB7436Yo7t2GVIw/aHxw19C/iu/pumn8/HbDq5HWHA/zTwLo
EE2ulNOgFF3S5bIGa8mcDXhCe0Ben/8kjCBCIEZWBcDSgWTW2GQEOOmFSV2zrK/GuWqWJNLaXdnn
Z5lWRhQRU0Ph0bpVgiDVPdZmOd1hH1hyBWD5H/B+hV8L6HO2z+vNA4GZIafAsy2hqg0q1280n1WZ
k1ZwY4VfDtpd22E/j1p6wvIuI/8V4ZqyyUcHQXer6amvOrXaUFlniXNbhibgVnnqPuX6hwCrgQrH
xcWy640E9pGy1RufbtRpuAbxTz9w/C86Uwa5GzntNQtFds+J38q0JxSagyK4lTDEUyRk2EU0O6zB
mqJoI5WUqfBIdKkqmpJJaxfch7k02ftFgfJvUEXNRjaEOGsp3UcGE2xZnEW66XxBIY+CtaB/WAFE
g02bmsBFrYVP3LbMokoX1IcBfnUHrRgRpJ5i7AKFlXzt1xNlI/eJYRTVhW5OwYFFyT/JDXqKtIYC
UOr/nhmTQBvZAMwlZaTX1t535VAjxs7NbAON24BafLuJSt5TMD3gXktTuOLCkk4X8d+rHKsSG3ls
iDqtwLr0rUx4odbsKcj3HMnIAgFfqAFI4hPRohSY98Q2Xsgbs8AnQCzWZ+TxE26Y2XWVjntu9Mo8
VOMH0HoPySa2migRwBAl7c2QeNzrck+LblZrnsXYjoUY/m3O0d6MkPOQB+NQ1CfF9R1ic2jj8nkX
wQZImUgzEsIRlwCt9VK7qeAsX1aax82KRrVaeALOJR/WARQ5564EcHQsOwJWZzUw328AAfIkm6bw
mVnI1OgGEXOWu+/g2RkPKn1d1uxFV3tF9Xvk8SADEuKIbxsjQq5J1vAhpsMxEPpGlNlXKPScWJUb
UoDtL4dpKShVgOBjYM93ROQXik93sfjj5WFZ0/SPQuvIVc6Xi12Dhm9/F5E6T3mbtBkjYJKeCDUs
Vgtt+ApPxsAmEkPkvY/wJHMueFATFvZu/he3dlhUng85m1ix6Ru7z+n3JgsFznk2lt/EC0l71ORX
Y/uWIRE7LTr52VkwfoAuMB9HUl2OLCPF085/OyPEhI09lhjumfE4bw2TQvwFnBDWWOayJDHF50zL
IKi77P1yPRNgTZCBlznfstv71ChBvSLOZoecGH2B8+8RL4MvaLczlOxgS65ZEUEzgAFuAG/BR7of
zlGmFU2TAoZCmJDSC2SpDoHdjK3o+tNIFsPThAd84Z+0z044wwFpNE6XqC1I+XHmNsOq3ecXT05f
KeQmZ+jivYIlzUdVT5iuUsZNAxE0L02eiyB0q86bTL0XCwP1esqoM3zJ/AWn+BIVj+q1qXp7X/Z2
+hQ1qzt1WXJ1IdxoOtMaAPJWLmUZTRVrvlK/6vWOIa/6BS1rpj3fwahKpV7TmLbPdnifCA5OXi1U
V/0l4FpTjNRDHO/rE+3qrdY415ecOH87p8HgL/uEZhz0esRUVxaJ2PZfy3Z3x/SqHvl5PMp0iSuV
REWJblzezmL5R+KksQo/WDTroAGzcMP1Puvy5qln8fEe7N4AUZPKUBHUx3fzxpsRVLSMavuLXyT7
L9UFrHAFQnIntpS7KWgaQdxlqRGbznsizQ7+TFrWQKo9xyvayRtf8O+JiBbCUyMAlzy8LtSTnVY1
Q6wMcWeFYEeIGtuw/AOA8aV6HLFeWWBnCwEdPw6OgMXI4ZBiTfxoIGxTmKiBZmonzIyopNs0B66b
htkgVOletrFcaufeAo94a6bJzMYEZkfNxJdm55RFeHLjwne5lRfz/udLiOlK2hqUUOoJ0RjjVt0n
5K8nlVcaNR4Y1xwozwwdhlAcnQpN7I5xsoZweRomgwQ2o2/HcnPb8bQ3HBa6330Rw2FOJpiaJIfx
aBtygegKsoekLxSzgM0GdKaRbGAlChJuzv/ptb63Ibr26FVbjKxL8N+p0u6nCOHVy+IuXbcXo0MO
iFjILSlTYN51IZI5I4veRQR5+8qVUfkgJn7XvQsPOxkceTqXreme5xsHYSGUi+ufEF+RdzW9BBqk
sVQC9UqWLthV1fOecPDEJgGEQfTrS9M1HaDZ0tI0NyaAKKXQjIk2otTFHx/qc9irOYXuKrBp2Pnq
vdDQmPr3J64shgLZQQ7va9glIwW7OeVfJKc393W/YBlPlC0Hznv/42+9J42ZO+TJwndETDAOI20Z
p1tiY9pfodLR0IbaaCoQfYnnhA+OoIJz/egdbih5fsUYURyjNS+HFfpfacpm7oiNGId/KEUUcucr
Lg+xTeoabZ8CF3OCm9+oViGBnSlyFDZqTuXtqKgIDFdVyNUT5tDu/kdtPrLg2oIwoA9vRrsrNX52
awnn+6XKX6JdRYJmCNrerqCCKoM4zb28ozPJuSMhvShihiSCwBSMpXygBVXc5TfGkIKUHzpa30fU
RwJcV/dEaX9SjlMRYBB0Dq64pPJHt9RLqerSYl2LlzfSaLxWy0YjUfoQsrn8KuIqh6tBu0a8k4p9
6bz0p8Eglmy53eG6Em7NJXkyNyMYlmDSW27cgJUgwRdRDqfp/CwclK++jShFvjMbht0vBI0Cs5+w
vr5HvWZJst+qUuNGt8vdXILzkIztVeYwX97aiypE+ybxs0ocLOU3nTVkNMo+U4epJTKLQ5XRpheg
S/lM+UdjyM06wZUlPobL0tF7v4O3sloEsBOjv0Tnuo1wKh8N4lyC23vhsrPcppae3vNA9KWIxspI
RlVFNCcu79u8HAnDTk9LxURI36dDTBLt4OXZhRXjd5PAaI0LtjuBxaI6mWg2id1fs7XQfVzHwddl
adCp0qjuMmBW4PIPBMnXzx29VvYTDs1oKAq0lgifVftQW6EB7r2SAiDjqh40NZrPZdaE3xo41RxR
W2cOJDQIqet2K42vZa3n7In7VOf/Pa1kjDPToZc1HXTH9rUMPVMNPNaIZYZQ4MpqUvOEzXqYxWiA
UJ/up3OR8SYd9akLp9aWAWu4vmL0Jj8B9mVOfpP3LJVUH9BjJkpthGwyIOSWzc1PI74DXW2xWomj
xAe/+xZPTwUiw0KpoHY/ibsiEKpYKra181h8UIp9zO2BIuR7RFiIqSX0oBdQdKgaXK316Iy1dMhp
feiLwn+cWcLbgbBQUpkhg77FfGlbMACXefZ3YtYjyIWzBNpa7zmDSrp43Dxr7GvxelZc946YnLUw
UbjGP4zzQebbpge1j2mUhqXy2lqNHZlJu6wyvKccXcghfeYGBs3v/EgkDTrp+oxugRdC8tCy6MoL
DDFrN3fwANQ236fphkqn4oGblsGV2Tj/+Ztb5agnHqQUljoCgguyfOzzBsOnGz6k4h1EDBFQvGon
SxEAEKX70swrc0KQk4s3K3ZrMxBvtrWSZ+U0BJZcOmHfBMl1xEBI/PEbOGWCVf16hTODGehy3Y79
GEoKreC8IGG5mdeX1DN5Tj6LmnAmNmRJYYmGion/N5JJ7UeEgqQ2i73UC5Cp5llTV6nJqbW0NSYm
N7v7lf9UkaC25uHcgEbXk1cs5VXMMQFK+l4q6vsRqF8UsVT6YOtJd7+cYDXdcLK5XcyPlWE/vBJM
5xjbOeNptvwvrdUakb3C/6xHwS0Yp422oxaNthF21viIG/mV9V7WEJIX3hOrlpWWB4Tmcdtvyvp2
8v4B3/+NRbQlNSunnbhLxv95xZDH3P0N8Zzkzn3aB+r6pnP8J9+NUQRAIXZG+dkOdcKX/52/KHfi
ZZMg9KlAogaRiz+dezjFBwAZuWQ8Ie/OLvsOuPr7+304+ipC0eFr/jzqp53KPs2hVL98Mw0VH9d9
AOetQsnC0OGc2sZvsMW1l/vuaZ2cdbMz/RAvCFs0Toxow1rnEqr3zAZcIuDolc404VVrIbTjfwDJ
cUPWhtTcrW0Eg2qwGQVwx9ZvXU0EE6qEKXNSVVsqc2mCBg4jw1Kzmh3Iu2qPAu+jdE9mwkx4Vnbn
h9FwxbREuMzEB6JNYU2qKsDP1t0bEYSKvSkm2Gs1LDAuYMwmEVq7EIvNtxUy0QTOHznIY8W/eziI
TyfOLSHckq+Y/0vWClt2hLuhjmcQdocsCplvBZQQ//X4XQVwmTKWDdVxcvoQcJa6JPYC6hKlMYL1
eldYBPKo8Ke73wvZy8MPaQAySRx4TPWaV6IFg+WdAsGu7k5ysURK8dIHOHbIOXcAVE0AkyUdRgFi
+rFWOVM2IuOIJn4CbJqsOaVxENOAuqYGONts1mWBvHG51haEMKSa8wk2JxP7sTgiZbhOkPXc+Yuh
SwCwxlVPyQOwttJ8APXN9+ehl/yzut/hGz5gLXPEdIBe/DAvHtqE78GY11Ilx86zmbQk6FJ2P4Ja
+z1Wy66icH+beJnvmq95ABhg6paKNQhNOm9XouuL90uJcqe3GpwLm69lMMkexwEjL3jJjHHlSPPQ
YHuydy2CzCGSRu0y/XA8P0CW5lAKf3tiW2cay9n974fa/iJb6+EERAAYW1BBSSXIzqwkR9guUs+5
pVw65J2pX51m1q+SEbRzztHqk4t+B/52P2PqRp9pPHvLQsaHlK1rdieQpiIu07w25aVn6qa4ocgx
Y6aXjDmXdN6kA7e1vhSjTs1YWug47FpID+022uj33gyAq9wer3ewF9oF8vUHwheJ4Z3t4slWwEoY
EBSzfRNdYRCNBBVpMJn8v6++xOy5IjpXzhQPN68G+4phykpRyr3S5bYeeQeO4Jz4RKHGq1WlZKgs
4MduGil+110I3t5I44XQa6chVJztAfkgGG7YRU3BMWpWQKUbwBZ2U11CT+UwsbULBYtYm/cRIHpG
mvAbkQ/sEamiPAwCsOB3FSTtUs5hIibB1OksqFu6ym+vQSWBDE3ASjHEhSYtvZxASbduoooDz/h5
7IxFGROUa0hLNcRUruYjAAQlNGY0ZUDlO6aenfVTnNbdHVh44W8FPrLVYMPLIZj+pzI8AfsH1NJ0
QMnkADA8Kxto6OY1NpaP5BBCR3B19mGK9wTitT1mUXVtsOgDil28NstGrV8Cc3Cz/8bXM1pJ0hXI
lXMRuLHRBNNfxOpeV8viRC2UReie+i8bxh03StVtiIldnEFw4Sg9jXivMIWMk7lzXh8BVoEcnE+O
H3MHhq4ZSWzU+xu62xiyMtARW6NsKTSDoDL5xWlDZE6jhwy/7Tm5xoAVM2YCh2D+8hVHTj5H9aFd
SLOixfU5X5lCjX77hYbf8RfFMnSp92A6tCATWPFrMqQSpuPZER7PrGyvDK/scanSLygBJEeftPN6
CQbnKsDrYWNgSmeYh6JN+jJk6u2J/vm9DS7nu3QWBniBO4Gl+QbXr5Gd65ZNFMNJcDjBKt/xKcPB
l+tW2NRQc5QxaYFulHlr0mCPHeR9/IZhZ21JGTm6/WwaYBFRXf6dUja3Pip+30S8Um0gEV6MYoWu
kvE2jSlxsZer+b9pC665863Kj2JB0TexpBaB7PGLsgtmFtg4ZBqMpWErLLzjVkJz6QMg+p5kaRTU
ylq2zbRsU8A8l73ZsljBRqT79V2f0f3UYJ5cGhNB3Gtfi5Ei7LstE7niggP4JiEzuRZAEBxVL0mC
MAFBZUW3RfmjszV6CvPeTKbqczfVeRI4KaD6jbS8wCGoCSwjoGogPd8v0UorDi/FyQ2ONr15S7Cg
UNrrWikPY0BI2m+h7tMGywLvuaRJ/vSF8EG9sv8yd6Pr8csOQcXLhuVInqWI4jEgurYi7mbF73Ze
pxajWSIjCdY2htGmGgihynfqV5vfnnpLtb0Ax8o86zijo9SAEjBAtseK+/ddN0wA04FZu83JDtep
/LaX3pmeR7F7MDXtDNZx+ORb0VFIGOyTYrAMzGUKU8A1G0Xy1RwL0NeuqWJog5Si6yJutBtYubOs
VXaAs+mG1F+VR72tevAXNY2GKZxUFU/3L8z1ie5LJwGDi3IcdnOwo1x5zT6eCSq6AomwVe8oXV9m
FsSTXYoQMG9rEWvc44w6XtHLSueBNtR7p4vGHSvL8WKlyuFs/Y1LdzZxxnRIUQiT+A8/xxzpT3Aw
pLBdag3WWBEQAolibCaYuepW/ooUdMtTsc9/FCfp6xyrWEhD0WCVhpYGEZ0SG6BOHkhppN6rdCG+
Pi6tZ8o4y13527OIpcL+pJRMa89tuYUDHSaDYKevitDPMMfxhTBTo2T2r2tZtmFIzMrh1nidOk4k
AzrEgahUjEgkPDMLX1Rrysnyw+o4YPFM5xu1DZBHdf6HlOwJ+tcrjfrZRZuzTeEa5Iu4bNcN787V
Lol7mQTf/qcO8vRvea9CyQ94ES0WnMm4yS97Ise2SDx0EB1myvM2mmmF2Ftpd9C6yqXgwNA5tuFy
It3YIJMjxJ/ioWxOtXDgo9jJDgtrWGRevvXGvpDAOskicvxVQZlKn36//kjA/MAlpCz/i9IpaDtT
+nYyuPs/wqQj2S1M2F8aG1dmZzEHa0agh/LWvstV5UxJAA7WzRbRwDcYOyY6CFHuQNhxDH0jeNVM
yXI/C7RPnPTUkz/4kiamSskKnT+SFodPO2gaaCUIvO3XAzvIcG5K0btP+zIAMKEA7MJ2Gu11LPL1
G4eDlcqJPBYrhY83yTrNIJGDbAqLHVwOCw7P+tE33lX7cEbwHO2Fzy7M17eUK1Q3XY4Lie9ZEUpY
x0oq7V+hm7tWS0cd7HkJUvA/THX/ypevl7kp5y09ZmbHhRH7Fe/k2OWbnd1uziu1VDWva5h0fAJJ
PfeO2DRILvCR45VgPiB128UyD6TFq/7KdK6zS5TTE1Kg8gnaQZD2VJCTNHCalA/7y5rscuUTx3Wh
Wyzqg7tOMsD8VkSfE6zFEiglL/s73o98Wcng1srPhOqA8OdffQ4RTsghIW1fH6r/wMP84e0k0r31
2WuTvJyCWjhIGNxxH3Z+DAJaiQWpdIdo+fBi3s8eQhQY/1DeNAls7tW3AdQDm2tA5EP6+zXkvIe/
pPGuvSXjNdN6yoQeTrt7GrQ5hpEgw0J72JUm24WBtZdJHWBlKRrwC7wrPD3g52dSYx/VNZAL12Zu
KTwNHzB+Rzk2JLr9gYx8iGqIJPvXFtb+kGSAMMmQ8l/XR8uthH/6pR7vFxB7IsBrTDR7RAMfT6OQ
9TAv1xLjidj/i90G98sUrQ8qRz9Ou1JqtIXeHeBVrNdIrug7heY8BFUqj39bttMLQeb+9lO0g8Y1
SedlQ3u8OghLNfS2QsmpikSsTWYMTvRrs6hMQiDu7mXTBTbcwuEqad/HGm6y5hfLNQ+lc1zesQIA
CNAhrYlzlTum9RVj8jleErhNDDTEtyAIg6rP7e0rboc13kgHXTnBvE+tj2h2y7eX/msaqB0TCab5
7GUovu4BW/wn6bqIIPoLB29DlVnljSB8I3xz/dxuVwK9KT8vXIx1766h9zW11+ZXcb6n+D0gc75a
wWWTd4W37bxlUcp79oSiV36UK3pGg4pSTmV4BYRxxEsu0EekbtCS/3icVulxeczEGZaySkQSYRP3
tEgpJTWocI4+ZMFyBTFn0tqJDRbcsV//hojTcwND3Qf3pnPYxYL8HpzJCa2IJ6/iNC+HD2M9wft/
5fJznkhSKBBE6FOn7/p225MQLZa+bU6Pf06dLgn07GKw/C3LXj0QVjkaEn5XMQ36P9EwOae3vc/O
VWK+sD1sH0P1CaO0S0kqkCVSPWQrwr208nWb+alW/FRKq7jfAfYuctWPd8uPnhIVTdTp+la0n5Z4
X+79H81NAV0zTSUGTlKsTqkA357GjJZNL6c7rBHAScOLi+gGmFcpzQmogKMAjclGIOz3+bEmyZKm
wvGzlYXtx6n2hHrp6f35W6zjxPKoh587F3czU3AMRbcjSsYos3K+Xcz7yI0QXk7a5C8uo5yNW15X
UtD5CRin94kNjamfGfFQEyFsaFDM+MW1f2FvufIi3h42znWggzh56uAeFM3Q3MT2vST4pg18r/Sn
BS83mzySq7ZOxv0Qk4zxXvpz33qTaJ/s+yE4axriaTdJeQuxJIOE1MymxX7Ekcf9nK2ShsqmkNut
MXyzTPp2jmyAkVzJGADPvN1TSXidsq5I3qNDjf1GZhWzfPBoQi9le9M3FyKh2Pg9qXcqqGwHgbrN
OMew9sukAzmICS9YGTSybm23dvylZz/mIHThFT2Xn/S0MKMkQ57tSmzPWAbvnIbzHssHquFHLUc0
y/EJuFrsiNTjmw8cFe32N17Ez0ecx+hdkQEaQgcGqoQ7aLklzbFtTiUbeghWW6hOkUQQznkSpTiK
sW9PlWSPJPkpyA1jdwm4zN0wR87V1NtWPppzsuO/g6HDLW3XTaEmQCDFinELF4NbY0Hii0CUDw/f
Ss0P0EGksa6oLsSELMxBlcY8CdNihn/tbz59YUA4pfDbWlFR62OlT+KtciJOX48+RbRPWsV1GeN/
IWnoq1ZXo1Md7bw9ggv18QaHUSrgPHdiTyl0iUUImJmzjCaV/Ok1xZmQWvMdsdEuPZlscNWXw9Ud
J/vZoFTgbKY9h+mNZe07Uw45va3QnWt3JyREVpaSkmQX7BnIbJVvGTWHlQ5MT6TWUdo+j8QL7eHW
9Sw1vB8DTH7b4BfDwYDpKStoGYJy+kz/2UphccvoXd0Pm069drwfJWHOMJXm54QyT4dmSGW77v1/
h+gV17MRNMXI+Bg43viN6peWiwsAkKTIHVTNDp5O9JlWPxhvn0qpQn2VZH4JISw0JPR1sAyPXG2f
Jj48VM4otuygTGveI0SnYeNxprOyeoZRTtG005WrRYadxHUxvuL2AGcmOJwcMe0U0dQOIc0sMFQh
RSQCHy6DTQ+lKN7FoNxd6N17RBuawTHkZkgJaId+57pZZNzCk1ItaeCSbgCInMBCVFee5qAkIHmc
DdYxvKvSMlvo49Jjv5r6HKlTWDggtzxJstOAvkLhlv5yO0FoZbZm3GKfg4b7yREDfzWYl29byPvv
WdLv3+BNQ6G9tspczqm2lWSh3MybwEHdnNLbM47fOfKK80Gq7LAgWRed/FAEtuOG++10scOr/DFe
2Ip9N3yyJUFiS7W2fLrP5sKkVPKXOJ4QSF5noypfI2CEJoXq8tFapIuPhUmhDVg2wgnTvVBoNHxo
bDxJ9vmK9G9woka4xSdnariXSgwzRRhrP1jli35H8khYLSQCs7vDIZNaWohjcuIl5CLh1jRXZfoq
hf46e7ixcK7YjmrnqYXRVxxM18oQbGzfJbO8a15Z978x3NDIeOYfbULXTAqwguEeiDLR74kmAAQ5
W/J1RIXdOf2dmATvZYHwvVilES5cNy5s7qTwm6KGU8UtdocRZolUR+eQErFbahiYN86wwJwxN5AV
pXe/n8VpVySpLfQPsa7fySu+tP87MePIUGmG/RKs8c1FCv4U2d73ijbpoUeknUIe+sCxSsxCfHav
GBxsYJCcGM91q7Q247XCC0NKd4uu3Z84ukWT8PsvzJczIFLhRHaeJCUzjjdZlkfCiNZIJxWLLjtb
LIlTo1INgktXsSW2MxnXU90Z4QLeY8lK4N4PUZ9/DS6AqHyXiLA2A3ou/D2Dtmg4oJ6Zutwj4v0x
/lefC8wbb9WaVnnSoS01owfAP1bvueJxH41wtLQqTGp2g/JGqfRPbhN96XyQuq0wDdLMqmimGMpj
2q3BN5YIHEeMWxDm1XX+dADqzcTEwJC10b/sqt79B/L0ddxZScAM59QdWVkIf1U+syS9NwaVp28v
80z/g96nXX9As3cnoy+sOS787apRUgd/xC1n4I86IdMkbUA1YkL0BRBTA7t2gxHisQe2JDT3mhGf
Fz79zfVaGCNPTL670/ug2FeYliQ6F4UZS39Mdw/zSmX63d7YMZbyC1VGe2cO1OUpec+fjA2csuYH
Yifq77VmOQnvzI9GggxoTKPk5qQGqISNsxkAXqi3dAVCVM6YQN1NRX+ssTDErbimvVazYqTTtKst
XqwwVOXEkYM09D3NA5i9fvpPK234cZ30Hpm+V84RXn6dHTJjVVxoTjVzeXGG7ez4x55TVtMlc+xi
v3+Y7nEUnimZHoWFjs9ZRVEiNuzJPWs6aXGfm0W+AAPFI1s0tJ6cj+sEO8CQv9kzlvP2TrDe4EAc
smPuwdptmZi2C5Bnw6yywl/qng1ojjMW0h7SqQ0MR+/FL5FHhASfrkljJg0F2Mu6DjB3HPOOrjuQ
7DATqEGq/vmfrOQSNeFp8Q6Vw0XpD7AkJGJXeXkRKxRYfSCQBABxfaxPWFJd0d0GSPA82NsPOE3+
6ct5kIbj/GeBzA+fwe60JRzshB06Ra9JEaYWUy39VS/zrIUCubxjJXR4wPZwY8HQ8reLSI6/xGjL
xJtRTPQWiHFY2Z2et+HtLpYVYdoY1RdNGLPfcXAhDZiobwb5x/+it4Ydfr27p8wgHuksAtXTkzZw
aQNyDbqJN4sQQGcmBe32SYWNAz37T2quU9wILLZysf4uf0PxB1bcDWfMUr0ex5yTcMNXPTm0yo4k
i6PCgLpCAGeLZ+tyXGN9iMV7Vdvr2l6AVc4GKz1oOlkwJIkTwXi/dZTLqGbAJAYBV/2PqHCC+eOM
VKtSBPQQgnW42IOLSJ9YzOWLKF7mqAR+IPJUfjzZ7j7P9YRlgXx2XQ6ufcJ19qVvnaefCXX9mvxu
7HTv6q4zHJKnpElztU+hxIpQ/KpQn2/+ey6GHtnjPYyGTxvJWiph+tu/fNZmBEytKevQUkI4qiAb
0IDmKFAnMVrVxEwqPO/Akr2AdX5LrO0ltT2/cjNrssg7DpGjaxPG8hIxWmEUCxO950CwCVNxF+/M
kW8lcK713DUIEiQrHNVLDdPb0QdvgBYfPoEC2DrgDcsMzfOY0lTGj2Ed+hCQiHPXAZ/xz+uFGepG
lwOZlDAKg5hqRK3DiV38IBUFFQuedUkKyFLikRGlp0Z2xzzKmhQ1ZQ9UQEZ1vZEsq5VjfPm9MqHI
rb8AXyt+UxiT5Ih4d6SY1jgUWNvZ+KMuyHOWBdWoOSbVXP7UpXPDqPC+EDNnumTmD08a7/kTAh6o
TzByrenmcIGTE77OrPGyFIDd7jAf+AFxBk+VLUMirRAsA1wVVV7iDL7OMaNF7XJ/4PVCEuawN0gz
o20dxzA3uRdXS3PnXsd/hKbSGEEhNoZ6+3dLvyeIn//pfpDrOFI2//8JyeJOPICosCJlAXZLSn5h
k4lG8B/OqpHoAQbektIJRE6uwUACmIrsOhye+bQ1GaajAW/tNT70Ld/yXMlgMbXxLwa4rh6SjNYG
aAiL3YNdklC7VLQJN2AP6xBOMBc2YCDPPXF5OVdOf+wB0kXuWMPV/oYHpbouSJXEAs17OouiElWu
+5w052iWAEJZDKI/L3UeJMgKIhQ75kvmomc3b0w1CtPxMR2zNPE08jypVO0u+BAq3gdufLiGSTvp
LCxApwBxFnWk5t9aVsdDiT1MB7dhpijPsveanuwmnvPHeN7h6tSg/sYicMlps5zlRM2+RJn1vIcP
rKTpqsGs2uDJMqFS0A+A2lnxgVmEOoO2oNqzRgeTXY1VytuKgBETKPQ+HN3k1vC8X84t+ob89Y0Q
wQRxCkxhXmBltP7sJtHNiiOZ4jKkjgYYkZvCDVteMb846x73/vbr+LsCLqGvA+pZ2Iuuc2UvGlDG
mk/HzPnFAgHmKUKBGtA/KED7W9t5TZ+VypbUwCRElscDpVlpNTA+sVYExdBmEfzTpHMRtbM8E3dF
ENXXJ0QyWzw/vJnlqBo8P4DnEWy/rKKVVjqjFubiQjwPSEi8gc0S/tSTANLP3qiSUjILEe9wPsIb
Lavapjy/884tKGpHFxTkQNleMTdrNXaubDs12Stnc/V+fyMYuLI45oQl+t4TvCfrklofVDZuV9a8
94ZM9WeTG6MohwGJJLeCE+Fh7cWQ5svmmGq02zAuL6TeYHl1w3vrYmnv6a52Ht6medqmeyuOhKAZ
Oo6LBD2wG7l63FkjCYy1jid9qzyVCA2KVyJzgcA2R1CB1l4Rl+tHa9lqAD2ICWRyWhwOkVQfaQG3
JYjT4lKnFGbr94ZtvmmYEBvsxufPx43auPIKnlYl15doE3Tr4n15Wigyujimve7k5Z8ODYQL7rqt
lMevb7fCN9ewHagOc4JXDrfKbEDKBwWatGmSJbcifOawTFug7m/f62wDXZpOJjAoE+Xh9rbNKT/u
VMQ2EBZjOg94ATehK63zvrJGA+ULz6Skz8xt1GTgMUGPfZWV09YQDjF7zqozHAEXkFMj5HpDToR9
3TStMMxqE7KNCRbDzT3WMyDz2GGmj3hDLhnLZOmvYNdTcj+G0n8e0dFl/8gibpZMIOKAlyvEkQyP
A0wV+PgMuwv+6FLWlSstcImE/s6x+WQkDsfwK4hZpmxA4eV1+4rMlvDXSJ8xalxyXoaS4uG4+9Vu
50jW4ecbxC6G2S4K0oDnswWhQYZ2uq7BTer5RsWJyvJgPswc4KJ+kixrRq++WVkWRpIzj6Hi8cLv
2+/NmpIYWNoAAgcFvQDeFcvVwQ9OVAgYFWPIudMbEdLsA7F6Z0VR2+sZYJmoPwy8l5vvrmLXpo96
okCREsbE6pks9RXAkxhV3sI1uOq6Lpgp34mm1Glc7kPaqS+Bsl8brOyR0rDXoPmV4MLIx3uB8tTw
AjWE9hwGkN5lsO6xBOXaYrkTYzbXkjo6oT8l+wmhJoQ5KPAyQczNgTKNyQ6LoIqJLvs14u+Z4gM9
d/uvLjvphWaUcJ7KnGCAOuMjRnZi+5JqQws9G74o6WiHImYSiyf1it3PrBLSI0QK8PJukBlHp4w0
4prUhldDBSOZJQNnIA3UBVX+okYhwbEw0U2OqUYqzlHehH7Ug5NJ4vtiYrim7nN4OqPRWk7V72q8
duuXBR5exKQXHGwKR9HTIaNaC1BVcWhMnpndXsBTBHR4+ezew9o19X/K7DJsQPCf5BOWpHQA+fxd
t+UD7tIloOPlSh4ESwOr7PAqYEfDAQMm97FmiiZYX/a2vO9XNvQRkCC4Fl1EA+EyO7bGwrNQZc6f
cL0GgrRKqDQyTGpE8/b3QiJKufyNLsUDYoGtVfCYRIHvkHyghx8z7pCS9d3dDW+yaliOhaBT46DK
lxjHVJF9cpdNFP4RsCfsDY/qWIrVJ6KWYvNBDJ3W2lvB2kAPOYFHsU/wv2OewJgwJQmCn2/2aE5s
RNs1mXo6dqmIVhnPAL85naSt0pC1IHpZ+eIQx2fZe5CJPQgkNVCo/Z+n7ajuwgEPCzWjMKnKLln0
DunenlMqQLq/EGE1p2GpOPtpGfhanjD3dTh0MztX+wlqM4n87l4puRDSpK0+GH1oKD8bxsMPoPH3
ty2I3VdBaDUMSBG1b1ha5mSDsCUWR5Mt+uB27VRYf8jjsOW+G84aT4xvW9aq8j2FXC4AUhAX4+0R
0eGhiObMbHIefFvHvlJmY8PEaUHtmWfGb9WU4KIV8/pl5NyVD4EeEMWYQHS/BpF68COiYgoQ/I1q
aGe4FzrKDDaF9mj2+AogHjPCia795fQGAJ9G/sv4q5H31fw6fEu5Sa5GwttLmN8XzPrMFc2IuONG
B0VxlaJDKP0y9BCzIQJL3FbE+0HAkXXnFvm8A/J9U+em/frfB+5frj6svHNXIgLjk/NbCAF193UJ
lOTckBkTnQbMvBn8CAt5wnhNs/0ZQaeIQtbBNZtR5C+cUQz5q+7SVIMk+17O/kSxHhNHT8fXS4za
Fy2bbqXsIXQ5xV3UQXjgazBnU9vtwdX5Y2Kv2j3L+yqX1gCBIi80jcvoI5AunDHW8vjcJ5RbcwJ/
DEf/S6tfhZAhtIx6J00QNKrr+4iyJRghDLSSKEmny1NNsUgvWUcd2BaKc9lZKWpt05OeH4zTwfSX
kyIWowMUo6fvkxSwn7f/WedY3TJXzSfd4uImbHAMSp2HVpkjYIlBcBGTXfEoLJDq+jKtS0OyoW2l
vKxaG9GjMz6Sr0of4t6ZUeo1ZcjVMpBUCyyTJCehvAGRJG2prP0Zx+/8pqKoSeC/REV5h5qvTdCB
Q/WhsGy/KErCj21+i/qSJLiI7oZ60mn3ukRkk70v4S76CxNHNclcNg3FkfAl6sidaXz2GDn+Xn++
GvK8/RWeuPNFzxLsutnGVdpZC6bgKyc5T1cVWD11eQQ6T4hfL7Yk9yWjgvNXwHqfkxHKWLIlW4c3
li1lcszsP0w3K5Bb2BnwolbYxsMzrlXelotHchmj2uedIwdrMybtUjHnpFNtHBQJ1iQ21qYNcpnA
B0+CqG5W5agzzfNrQxKGYvI1jwc1JtQmf45OtBGECdHYZKBGDIbDMw0461IRszBd6yUFzioUtx+d
5/yY0THA9g/gPrQwWSbfqHNtEq0Scwtb43rzUYst4RZw2EXtOn69/1vFJJEjnGfqCY5DMa5TTgzN
tyrNrcnnSMcBmIk+5/DCKccbcqmawH9AhkLQ8E7YnxlQvVMzeER4aZW8GEdcFe4sT2So6obtZcZr
lPksp3lUD6RUOJpMLFCTE05UqGKM9kiDSUUAMqrz5oOCziGdu8TctrdmlEThFSNPZ/xKryHDijmk
YbGGvKlA4tVRtxYfAl9EmJE4DPWhmDH/XIAa/+JA2UDqdNhF9zGXGFm/NyWFSRiEl96uoiwy1tV6
YOVbXbjkExX51lPuF71yKBolYDqFQAipR0M0Esy/EoXiiukbtHgEAWXpsxXO9MIqHCn1thX7DzcX
x132HSSYZW+MgxmV5MetCRm26ySKyet1E0gjxL0KxuyFvLVqz6WG3v1o1ZWLyRDDc/MXrmU28XEf
VLi0z/l/oHxb4n2melU+P4XnFcGs+Nn8XRDJUZk8zJ/Gvb6LFyRAFfWX5mxxDxfzQnKdMvopSw3v
zflPNWnSARRYV1P1JV2xMLzMCgTIziH01n9xLiro83tImw1weBElWr1XrN8klre4yx2++47YLVZJ
1ggsovUrk4QeLyB+k5sXr80i9Mt1rM9Fc5eyqNNloYsYy/ALPJ6wCNtojASJa+tV3FLcpCqJM+Cw
eeGD7+1sPKQ92uTBbr3kwfBDREXWfMEFkWoa5BBrhKS5+uKBpYkDanm/xsWheSWSkz7WytjQ0c4a
LFtoK9uTWyIqwyjtM+KNrKS5A+GDPH7+8L6vufp+mpdDKAQ2u7ZEdQnWZaL7PtV1hqoXCuLlbKt7
mEuHY60NKM2hDS6ITJfYXgv0iLrhoW+4nvdMGs2MBe4Y3+Ybzx5Sb3nVpGpBCRypPNw3sRkV21Tk
Tkfg7JHJcIwizXdX0ocwVFXMaFvGO0siWRSpnEfxYpkSEgXsvoe0U+jeghIgf51K42wUlhASftM7
yHxpi1lCnFNEUc1b+5hTMo46jasU3agByqS/kQz/7kKVEhSW3hbXCNGm5me43DfDHEEHIQ75I1G8
9kaP+BBhkuW0qFW8TW6GJApFKi3H31YcllK0ilS7/v/uJtsFWcdsxi2djItCxHUg/pMX5IKKnnXX
cuNfiSiT5VR2b6RJHV1pwesiEpdXYtXjYV+kXMW9XDULZ23AWMwaAJG8xtv8gkhc4ty5uudmEIGM
9rrlrfKAPRy+znpA8BVEHraSTtrhEDM8Cg4aV8UK1oD5q2zJPzzCtS6XVLRl0+Tg0ixPDAbeLsrg
ZpQiSzr6JcudF1VRNa3dNIGQ+xiToPm25hXxwKA5KZBBv/G47UcR8NiJ5ylKSCQeiOA6XsqthOCI
d5HiB1CaZgFyUHGen4yQLU7Wa5IcO9Ecs8p/0MFzGwUwnznZ0oEoldNYUYqVRB5FbvIISSjzO54N
upwlPGJCKaKEqwhzjt3SAliuVgHvzxzVJPlODinpYc+tc9yIPryKzIzG9EZAWZA/P1xtlncBZika
QyXX9WlDRJQfZ5y3sNl4kB319JEwVQ98UHjeBd7KtmQ6O/xXHoY2jxWqs6v6NOEmQHAb/SS0/6p7
6NfcfO/g37E5y5edNgMxFbEdmPGGr6wwRd64sSyZJncLTyZcs6L0hXm81vr7+055woKlaFGxmQeJ
hU9RIT6ipMNTUFFpDIAPompPGgz5kBdfTmL3qJ6g/C8phv4xoHxEVRstO2sHY7gFj5h1K9vK4opl
3N+LSqOQUaacoH2KB9wJMyEGR6qDuwa4QVO08dhqawrsNWOgp+Cbl0UcVfY4FKx/+h+3RT2PkEBv
Oii5RanGm05I9+i7M7tzDJ++dwltQwtTr0VyvbPIagJr36O0awez9cFYwXHcU20/JpZHEB0v5ziF
1m9Br+uySXAE4LRSqfs1OT+It9AbTavz31k0gCjATYoZSf/XfWnlLBydmNGD19saAE2LwGzsImgG
Zl5Zuo+P6djY5WfcOpMpt3yybwoCj0gRGMmcCQzGuu+AYxu0qE+SxFUJ3TL5OT9/3B+IJ+OPTqnG
FIhD5qhIl35ZBD5/8mBpHNO5SJ8qraYmXmlRAEXeRthOuXIeBqBRb9DEbQXCAwXEo4/hVbX25TaN
5Yi5a28jiKGS9owTjSy0C8AnEnDbOIvdks5s63I/3eRkz2+vfXYWcu+qDdWObsiEjjEbxR6zZHvy
nP+Ub+/2JBoWNlbmlduOsAenpxQoZptRvKKMMDQTiVwNUN1Md2o00tscMZf6pP9Jdi/GozUkM2VT
XUpmqZcxTcvJqb1YkZW+CI4R+GHdl5gZ6+JpewVbDm81WuB36S/VTP0+WQeHAHACPKuzuCiwSgCm
Iyig5QSYr+JoYwEzIIF3gFlNJUZiLoDJHPEr/viPupWo5Nxvev3v8oJU3l+umH/OIeJZUUW/73Gk
7ALnQEeGzXtzG9eyWhkK6xuHJfkNBOSW70lNUYcg/qUeLqR20S1Dsvc2KZXPPx7qpf/BMRQ7KpIg
4QwNfUBavVV0Jx7hap9V0649YGmb7aa+Axzt9JK39FALBKubAl7NtvW17d4nOfzUzOG+mVr6+x+4
IC2wCRNbpgpuqtR0mTtpqHFT5PToCUSdrvOAHCyns/B2ysqANxCsWGHPgAVB1QzmIX/LMfDbbIAp
52DU4dEXDX8PQNs1HGC9HeJpAH+8p3Lir0WOaYRZdClJT+nzZy69w/KvO0VnjcTGVI1NZ2P4r9m1
z1TLTLtl/Rzd3KFsA6L9QqKsr50/bS7jlABglTPC6ob5S1IUxciv6w+fre2THOvshNygb9ZDRuwx
i7JF6GcOuSqbzkog05JureQh8sIm84Xg+yQCSoV4DIAfaDf0yeZ9yCpelLI51OwuzjtZWymJCHK5
I8Ywhvx2u+1o9ynpS+/XDYLNHUcYZT+hmbSsDZ9t7S6weZuCnCNHmYL/Sh5n4H71pZ4nDmtlvs5+
u+zmuYPDSmBRVcXPJK9XsEl4J+avJdy00/KALTc5sGSzhmCCrz0kB0acguhSkA1YTYC7kdoY0vKV
CrBQNCcETphEYDpj8lGdHnyOVqwEksiP7GdQaHDNDJEQW95rjWjeKhIWiXzHP4NF26XA+T/+ixm4
T4bFsfhGYkyMeJ18ecUBSlLULHa25cq5nRiwJSsMQIglRMYi0+vFphutbylVRqoddV9pwZgeZW5J
6IFOcdg1NZoo5Z1dMtiOkC5I0MNz6CgvOt55FNDnPbpALJIGiVuZvnZHoFYCIZ6CqEJgs53kPvyw
nslweIzXvB5B4CbsV4if5oF+fZvwoY8ZQ5xYfVmdLvC8EqNnrSAlbfZWWm6ta/Tyu/BGhZxsOSk9
w/bPBZcd2mJSLdQxL16Uu9eHcpxnALVqJWAP3qMymNBcsT6pUDfpJlPvR6z6wXUTtQY424bXED3R
hWR7HJGjTlUkP7sS0O4vXhpPQnari7kVAo2uwux1K3oYYqTQfCEtFTsKg2PQJmffR4gHvQoZCrPj
44xlx6eHnN9c1B93G/drbmbpnbZaScCqWX5d1qdWGzpOYh0LGEteev1YIUz0Y8coSGu06pl0vA7a
53qTa/54F5AbPTfQqO1Fc4gl9leWzweOGMckvMKfPTwrFPPm1SpLqeqT/Q3Gzlvjtjs+L0OMzmko
q2V0vyD1EXtdKS4KX5Fa+0ka/1YyuIChzDGMwOJS5mAAHZ2UKA0oa7F8wAbLhcv6094ZqXyPwZij
upZ9rF9OVS+jme68vkuQzxviezCy8ihYF+CC+PB8z0xPyp0N4zYvXGVGd5hS5jeVUzKOsBiB5CoW
ERBfV/OBjU0HH2Pyc7kTUNAMDQAGGVFHumLJMvaDPQMxJsIa0O7i5HVgdtkiScJLw2KeqwZazA0G
e7srr1E/RAXqiBZva01mzHlzmOSxIWjZYqq6/DOPx/jh13SC/Vp2/HpS7U190PFlwiYNJYBXDVur
dJf8dadq4dc7sy9gB/u1CIHJYNVaoXiMdeUK9gnOdpjlMQ1wjZrdH43G3AtkcgU4rckTLKEdqBeL
Z9rw1APqS/020riaP7qGOKgiIBZdCsd0+gWRLPBOrLeJFm3AsoLK6Rwi7wI7p8lBrv4TNYAW6/rR
ZV25Ho6u18CHqWmYyWzJAfW6ix7d0JQ8xw2ytoXo2RtY6sd2AwnMPJVCd4a77ZK5zfCvSLua+H6I
QHbxezNo9NlWSlxogSZpUtHlly7OVIVBA0Tm6P+euEG5nddgoRHaBfUz417I3R6NgRvdaMYEQKu+
ymmEmEsKX2NElENPfDvT2GMW2UuhWBzOyhvY4altqPTg5NGVUVQ1R3pQHPNjR2tSjR9O/CvFToLQ
VUMqdQhVna+nzBYu9J8+o65Y5Db605YG4o5ZfN37hz8m2NMYiCO0uQrftPrhUAGF2rc59dnRiCK4
HCB4gJY+Ug6XPE4h48qRBe/v9gJ7M4UFpPQPMUecFluitRXOgmz398RuHWo8W+ajlU0bppe/a2cl
UIEX/CwuVRHtNAJV9ZIsYKaDk5iZ5ARamqQHrZLfAH4Gb7i2Cn1jFg76sKSvYPFFN37SD+yOAFBx
ftVx2LHyBqWudkfCZqKDgTLdIIESmmd5cg4bi61ZMVjXgkSuzDCRl/HPAd/c/DyNoZvSUBwidO3n
XuZPTSFxJLdrYu+0BnemmxwbgW18YqH5FHsccQU9T9xuva7qFn5E1q0VzxUwkfCXrD9FWh1mv6IM
Ch3DOnDq/hidykP8GwjfXJ34+aWihpnJHoOvRB4xA2/ssl8rShLdSjnix5lbbFDFGG71WLLC/xxW
heYzeB12Mg30TkY+oQ7tOX4sb0Sc34RCNT+RcitymcMxZAGvYHUvaF6jXqyNAq9fwHsRELytFvke
rvwX3uLfLSOMS1VONiDuxtV+VlzIXtrhv/nQGKjNBh6r1Hr86/SRpac3V8Etu5cWaE3MdIwZmlM1
20pk22cRO+0a02ULOlACT7DRmuGjVbC1lL2nulAgzzS1iqgpQUjiqJAy5lfkEZJVoUC8syIZQIwl
GteUR04YD2fJQaioe/lCRVvJ+Bm0I0ViFHIyfLxhqFxXan3PiUyc/Hd1uro+CGUd6s5E6D17Ty4J
r6mzzhdKNL43a5oNMSzgYU9a07JCEt0DUTNZhLTd74CxhqiYSN0gHZvTtgpDChcLZDBlDhBZcYqa
SLgFz+Gj2mk2sZW/3hJ38kd8RCt1KUxFPlIUEVOl8G1VvZc9SVIFW6OkIFj8LOs0VWCoCY4VmX/e
zMvFFXUW/Dar5AbEBMIoOZB8RmtV/55IhmCsudaFMMCB+17YvB8AB7xV6LBTMLvZInaOJrlWO4xL
ZFjJOOoiiyW//UonrYtCDKWHKlDTgQ/D2DLTMAOyVV2wIYBbLUbZBiviK3TZOf19YJGBUE3tQ3zl
QQsS2i3P7UYi7IUM0/5QePqAuGHmSTbKkP/PNrR36kiv9jkKlMhklh0KcBZm+gOV8ZjJ2ntzMaJL
p1AgqqZIjfYnRCj5qOriJ3RitX/pVKsp+IubnekKjnQpSd67dVo8Nj6ffmKWq9MJbAzK3XMD+E4m
qOzUBX9ezN0S8AGfpLwTJjkNmuY+FfUHG9qdK/hYxkGUWhpog3FA+LjFU8zPbOeGX5uS9ZofELVh
pA5VnMt8/JeRq6AKtlUBZTt3vHjMc7Ft2UTFKQhqBsISZV+uG1DLc4ZiuzompZ5pupSR0S5nuW6S
wUEDaw1ZL5K0s3z1tfUVgY5/wbmhpD0QEmAl67NAabP+Jo7J4bBzKeSxJCn2Hyg1vMrLWsutPFps
Li6Wp/yf1KwuzG2QphlPd23SlhfSEnAt6fuSIhIGYY2XzeU0yOnX+t2mZvVGyhW6b6nWunzcR/YU
yiYzhbvcDtQ3Pp87jM+Hu3v8xkLUAPD/2/FsZ7pZ3z6SitpPECwb5Cut6Z/bcPR1AOaqKh30jGXd
cyjINWaJHQI8q6aqgSZn5uvbjBMJHgQ2lHlTkDP3VTGADlClPzAZRMtryp+ee6FWPG8uyIReHV0o
3n4+MzDiFQMbFLJ7+i2wiOBGD0KJIBPcRIYF7dgKmgZC/4lf7bLrb7Q7IphwnPF06zyORCAujRou
vAcd2JlnUByXkl8KkqQPqq4DY28Gzhs3kDBQw3ezSbos0rezswLiMYpYKEdOCnlnICVzShdlVRk2
rIeplIZoPVEx2P67PS+4aFGD8oQKsz8Lz3ic1n9sEl0ExOlyvdV4No+6jkht4qr4z+iyM+Zvk1Lk
IMqRulhu50XexC+rBTzxwcyBNkbE2DQ2zs3DEGkHtNdUKW3hFoiJKDsdry2+dTydYxE95GcZ2Npo
HdoOnSfuXkyGlbxB9KVzacUojCm18Kvn555yyw5qQSq770FHmNo0Lr2cRODFQyel+jhTJg9MLjPg
Kl2fqrd/8Q9rJhkaMLZ50lSatzm2sZbgChl5YYrVX627aad2twA8jtIhCJoOv2Dwy7/1eM0zsT3E
viNBsK5cWrwYNzEghCnFDj+YebpmROTecqTlNQ7Db3KnJgldIdz89H8C48/tSJ+CrfnZccNpkZkO
UFTUw/cbmp+oOotas51DQCNao9U4EbnbS3sNzY+1kL6vXMdkC6xpeeg9FQxxOmh1v4Z6UGQI7Vk6
pvk1pgPKy5TVm0dmWTg08JzQKgJfI/u+OVRfEjuR/NtGDejs/Y0Zn+plfUzR+ByGdHDu5Bw7zilt
IVtuWmzonLBPJODVztGOL8fYgmfG8n0F/Q2uIh3CXCphTxvU+H+9ho6Y9YR70rgATboRRI1nwSFW
Zb4r5WYKbFZc7tRaAZya0B+C25nQrtmjxAWQMb2tW0Xok2tkEkq5KpMIm1RJtReTukZdiRUE7boQ
kEY9LeN3U3KlRpxDTH+i/ufMXS74TfgjYWOFVB8JQD4QaZXGEQAGKrRBu+H199v/nnVGH4sLp6uA
ioEPZmJqNqIgbPlUc8efg4oC5Ax6io0tt8lSuDYG9TlPdth5MyTv+wlfGDWYKaRF9fY1iK0Cy7dr
nT8TAROVy4wc+DyTEG34dMG9EzyRyaCMxsl3g9oQIAdt35K8I5RcqZ4YNjgG3MeaHEe2Mp3pt66p
8t8Apz3YAroi8SlW/N6XL5tE9dr5ep+QVQqfFtdis+Q53gC1rvGWelPlZ7hg1C5seP6YMv5lULWq
M386mxAtqPMCe3f4yPH7OiorYRkFrGAJNxBhFYpexyrNr41tbTsKRA4Dok9GrRqBX0DTR4IZb0dr
X4KrQKFipmZ77h7BphEhdFvFoZfpOC6MRkkEePbJuYgPFr75JLOkGt397JnFD1aHntIYFogiVNsZ
hyXP4JwBt5/3vaVETvPfzIOxHaoGDP1vlZS9PHMlgURdycCH1SsMHzyZq3KVc4Zgpj7xDb1t3mKH
EwB4f94pjs3w12SwKK/Ljd5c3Xwktuv53e0KWcTTY+DKBRSUzx3SeoFeRdn4dHofHpN3KPrngNZs
erf9s+OHVwasMoyoyN5/62S9Uu9sSA4DNWCS17eFTXiTNrsyMS9561UL7SaQ+lRjw1DfOufHYUPV
+T4StCj15+mE5++m5tObksfLWgblwDFCpgtwWoBy7Z+6WjVD4T5P1nrr+81DCnH5XSu5WEzrPkTN
IXvniKdO4jmNYWxQzdLepcAZeg6NLCRqqeXFJ22mip6nTWqU8r3PCDjiQO3zcSzQKrq5Pll0HkyL
JRX2MFYdBH3dPCcS43dy96cSvbTfs2Wye5+eCVFP64YWhr8JkH7kKvy4Sh3yI08komQ2HcfH1ab9
Vj2KNwQkgRReRDHY2FDoZbmqEPqi73KKC7/oVGUERG11F3/E/h7nL0K8N7CzE+5C6W5rJoB2b1nV
bx8+92Wz4THwRyhL183M/jKfKbzvWoqUMJkg3qArXK8cH7dYhYN6WRy2zd6kEmPN5juMLu/sPwuF
Q4k7azdne8L8quBxiu7nx8hdkjv1u0ZoetchdIjT30Wi8E/NbTo9tRWYSz/vjmeYwRot1ELYluoX
igNA/P9wxDG2EkAHPmD4+A2CmeTTJo1spnzjiUzm5M5Wx7WiaO7J/nV6MEExFDm5lF3nLu7dkQ8u
n8B8XYMnkXzz3PA7ZdcFp5DPRmdeb3Tz5aPEIZ8NNwOlB1vWEQIxtPNSWDvvK5liH86V+XnZGusE
RcIcITyDLNJt/NDXr/QrgwSpJeANWxZEoWmkaULmAu1gAOIjuCaisJf1fbuBO7louuBvTq0r3FuQ
J3qfRRkQuHTvQ6G6IglkZ1JlfuhfQ/7tZYWPLz/Av0G9A8V1raziYnfGVuKbJVJ+Qv8Fqp12zTDR
8vKytr/EwXKNGsKPWY+XEdmSb757cqsvw83gt1DXZcw5FGxvCP4Yo41m5cuBzWc2WB3mh4nEo+vK
Q6CPTL3UU74LfWSUynStmX34Q/8x6dxStAt+hIXpCsKTv90fAEg1doTOEXmqWcwXK7Rbtr2IzG7h
Nrj8nEm/zdljhpOYqq8N7asK+dX5vXj6i/hF2tS2RaMM/Gj4l/tQgW6Q++/qFXgV2YL8y5LZBRdu
6Fql2/9Hh3eMap4cE08YIKjvr8nZRc2Ypxvtr8ob7eKmcrptnwKPN+1HJNX98b30qt00x1lwzJ1b
RKX987MJ7lL2T2bBrV1sHQxMuDTRbGwoEh1jSg/7J0zza50TJ9jM2+tv32CddE/gLZEDnKR8gcHj
zXGRCDuIzfDVbwfVRwjKy2AgmMMjpIYn4vakIC0wwUdXEQPFWoK93ZrWNWjl6kTqdghwOvwcCt3M
2SAqW6mYd2x7fVa0T+Bto4J36EHCvyVPg251FI9mX2dtNHk8HOA1Azt+LjJMjlCtnTf58rsxNGlu
SNJjDz0diUvnNfjt8ckl20epeqFnQnQu59xhtXU6NEq9RmRKlzJ6ekDMrHdlurTluc6a7G61vdha
h2sUO+Ip0Dj6jWfJjMajbYSo5RmNhKpl5PuRbC4WgJLjyEvuMDW9B5Et4ODKzEVuJyoPsdi0pZJF
ni+k3OMiTIl4FI8jWpTGDDPgsic+vR4pYLI6RMku6Nn1bKqxadFM/JJUkz2IkaU5Cvs4sJlrwqVP
JDjWb1yYlqRj+VY/XDtuGj7+FGeixyJTd2SwfDfX6wFMW0stHvvcGdONDXJpgkwG1r4glr8ByvRv
NwFf//DTD2ePUjmg9XD4pFjmvLYyq3yPhYRH1te/2jsQq5W0x+MI4C4q8zDFkI1kCISrtKYes1lm
ZQK3YRMQGzAPwmB1/w7gntZ8jfvL4AxGm1PMZt0gaKh7ZpfiqXUTAgIXZMeOvnz+QQoQiGdbwEoM
ZRJIdANU+0+wlV3OhzkxJLZTGnl4aiNxnAXwxeUjwylgRISnUPa4UgzZE8zXXTczeHv39sbO1FQd
gSKFucB/kullSh/dY5bhizBiNGk78kNOGVOd2u4Zjc70yPEeQhLFYcEw8oksNs2yldk6PIvvve9m
0As7DB9X2W2k6yFJMlLpBYfI0hmpiiy6j9FQyAn8cgQ+AG/YgpjWaromdKCglZmfaJSuOaZdKTQy
ZyLsiH7pul5odEdyIz0I9VL0tfBLejOs7oPX49dz6Umq+XmcnsMwlCsT5uYcx5HmoMUpNAvuEShf
PLDerVR+4meE8ER1qyb+t3/lXnkdLxYzx5meopQWyWtjq5KkbzdkYSP1Ycuw1vXi1qYzsdKM5ij1
E/WbW+Ch9kmUBktKRg/Q2TlAprYe5dx8yB5MrapsU1NT3a9Sb+K0feoj0Ra4/InoZjrrqBzV0lVP
P9a+XSW4J+ceTtt3HhZ+udG3cZ7if6IZaUnJsQdqKW4sHkmJ87cDvYmkH0+Ql/LS6z5dLYpRyTJx
AKgMW2jfzftWDw+Qdmb/Tocf3Er/SdB1eprcp0s+xRcXQmoiEkOA8A8Ks01+2K4SvtwQZiPzSYzp
1jxqcI+QYcjPrHgp7FemVDV4mthMjnxJCSQBq5ZsYIVctDcA4v0NrHzko1k/CaaILvr5Hd2xbvYI
5WMOB2MABqekr5/IW35W6F2Yaw5M4vZRwJVq3OiLLuNj/PwEN0tCWfWD/Fp6Qi0cEcNpaR/5+q6R
DznIpMamTvMSh7YRMy/x5L254QzHwl7OuKx4oewAa2kFb8xUsezDCYAr2n2pX0gHwLcBwwBZNcx+
+c/7Qs1DhZX3jF9hzTCgQNfPhjeoPU0hxQ6/tWYevevJayVb82s7g2SFgD2eXN7+67CDXvkZulyt
LeZxFzTJUliUyeqw+CIDySuAvXgtzyWkfRCi5W1WBsfuT3xtGzTxLIoMwdxYOf4n9z7Wfyj4lFRK
G8Hrm1CvK8Lq5vHGNlv2Wf+tN7KTWI1anlLuPKkkgci4+rg69ntlHLl8Gw7hlW0Hymh2iAo84ImU
CFnlZOjJsqim5fPJbp831TL4VZazHjGIr46sGRCCmIjhrJfwJ6EIi1idJAof6C2/EAwXXu9pMdNe
Gp/VYwIU4pSnTQ23/hlaCgJ62EVXO4DPfuKPXSlFMiVjNce9QumugBPF0bf/EdDlesT8W6Ei2mpF
48UmurCo0KHDf04rgzYkamTmu9zo0GPvrCaYOkONvu8urWrrXUz/Wm9+GoFUwRoKQkzrTzl+aAqo
skSE62lNVCc10mBaYc6FnrLZuVW5nBTe7ehIgJyHXWnoEmwl5NX1ZvGc0ttH1mb+5Nsd5nGphVvg
X1SIIOiPhBywj9xWA11Hvi/Iztl58jd1sb4gSmPxqygVUCbQmdfqGdhzZKecJ3H4C6i769okfPpJ
H8Fdf1ybArXAHFVubUlTwnhQfHEKifGZcAELNsh1AqXQpDK3OTY7V3C/UoJPMc7cPtcxxPNw+SyQ
KBg7GZIaliHOoqODsWu49bxoFDspT40gfaAlCjQEzb3IwnCMR2p6XGXWT9dt+jigWE9/Xbjgc2g+
JqN2qBROmTLcLmX8wZG5oClYWyPZWjVBzoE0qKyXMKaDJJhVP2p/PUZAvQKnhg01L/3J9O2ABW81
6UF1V0fiEm/UAfwMPayOkEcGPHHX5HsNsKbVSKxOfHzHt8EaiU8244VAUFZlCvaoGV4Oi6V9DTZe
BDvooq5JuZaJWyiXUbz9b5W+XbOv0rUM69WFe57RZfOoB6u7P46gD4FtDCJkFz4mQB6qPdMV7Nl0
A4cpQ/IGmjAa/Ya8iV7mXNWime7aWiGBW0SoEwdS0fiaB7g+cWNcTvfg7ltMj1YfdSin31pt3WNJ
OhfFrRWZxH84QwOGuVbEFMam09q5r8ULyTvsJdCn6E5qbP8xUIkxkQ3PiEUllY3dMaDyJJI2R3j3
rnJYj0+iLinZZERxLd5UAJAC3qQtU15y/5DbXbq5R8iNLQoXUaxL0cRs4IZBRY2RwkpIz4LNgFlU
rG/2ejIZvrKJ/hRtFwJ99TszS5Xe61L/SzIizn/3HEVQKEbmtBWJOn9NGhxdObU3939CRh+63k4P
PJElukrrS0YV9dBaU//i9XkCpevtFLf1d9tS7uPXI2yRWVmKKMmDE03X42VRlSML2uTYJdtF8eN2
xMBI591fcQGx3dRecyW2bnt5xpaXnP8F0mTp0wiMhkeZQe9eh9wjCX91dW+lauX5tqL3OtEPjoa2
rCa2lViIbv+ONp2GIXBt3XzRJQgGe2ZhFE/DazqUlAwuxUNsYth8zTv4VS0R206IrpRe0Eks03PN
tOnLcmEaUpOAmaaydTPFms2eE0+NUu1Dk768k3PTPSwj5NHcY1AjRTmbZ3L0dDSQcS0D49AQ/SJ+
xfiSGLPKIgaMpBGQEo8SpUzKVf94H+WaybyIz2ghXkrxZFq+XLrh6YH5NJXAd9+/+Al3r8r57quA
NHcSIKodSTPWsDt17guwMBC8GWHsoj/3v9AK5huh54RTbR3E8IeWuCeJJO0eMqJ8GoktxIrwSIMH
wpEAYPrhb1LUXrbrJlKe1OJWJeJxaIV/fxnsRI7AvIcU4RzWpDB86W0hrUc1uLTUxKLSIy+M+rT4
+IQDqoOup686Hv5cRDJbI8IPjhCJUCbVK5Z+lLcHLSS1umGrzpQqkaDZQwh2Ejo0k/HFMTovJazX
57mAT+ZrcSG0mE1J/eNxBMHFISEqBjyKZP4R8zBRVuuum5ytJ2MGhxX7jXe0DCw3SWlUDQEe2O61
s9FJXm6rOmaeEvJkcGYK4Zi9AKb1RK5ZM6uX2FLH50XQ7yAPKGE84Uw0L+vzxKqmgbriU9UR90A0
NQsQ06kNUL19xIePGeiRoClaRWNb/uJrVrF9b+blIUh7xUd7njM77gX1EwLkXlwYJ8Xq6RbZBXqY
TLu/Tg6FlczaM7KAVa+YA/TNJpB1aSWWhi9vPNz3GdeuftCrtpx9VN7/lGNZpCJCLNX3Xc800TRt
WElJfVzlGEa8D7ynLAaFKd5O7ElxVbr/UJjg+IJl9w+c/AXUCo4oSYNyZQct713hlvZXDLFerzUt
/7bMFzYHs3Clnj1iNcATB9WPIo10+Fu8aemF37nwS9fWJW4kJjkaat7bYDAkyfVNnRp9o1GSEbO8
mzZbfQuVdDYFU4TLOeXmR4na4IK86TKmcbqsjkbil3FQoaoiBIddDNhnq4268sHMH+bZRMj6/ynF
e4dANiuYFEGQ1VEeyGVnEUj8cvwAPoYk+RdHUmduSdSteZHgEk0JFzbZ01J2uV3NhdPYSSLeXR3D
qYnJeeI+Ny1LMG4FXgpEGwK5SioCwlfY6jynADOlFXr025bj7flXkROP9pUOM6gLibS+vVJGH8bE
EK50p5UsUeCU403tFhzwZYviSWwBmuly4qr/j3Q9LEd0bYd0aGbQCEYBfyP6IVI1bNRpHU4sfQoX
9bu10WL5x6KeaoJ3XudlIgz5SZ6AQrmHLqPrcBMy7li73+jhdbSQCENiu/hTyUVaf9lnuvMMFYVo
BCByokefSx3pVeE8fgj0Z54+s7EE0lYyZlw6dlpLnmQeqRdQp4cX/ViTzW4CfoLYtlcxyc6KvhRW
BVik5EiRyvz9EMi7j1kyx2NGD7CP4/WTFm2inntgkxm+QbXv+ASBFdVNQiAskga1OdaTSDLhTKQc
ZFZtXkAwS7sHAgn7mdkFFHylzVt7Il1UHnqpN3ZSfQgikT1P32Q2oLHWkTJ3YJFHoi0eOttw+xAI
OvPVCapKAZXpvDzqinVw7NnEPWZCpvvxS7JNB43jolvZhIUq7BcWMaA5p+AJukAiEOhBDhMPczHH
ddTuiZ/w5ZoCZm4GWjQYwYPanGCqQBhWGayBushCO/YYqJ62nlMLJN3Xbn2I/aihhXnF3osk/4oq
o5vTX4+5Lliyk/iiKp+GSqj6AsuEt85iafTW2LjpZDhXz3lPgUPHWtbkFkw+xORsFOV5YUpNCRfh
gNdDi8iMGpOrJOh2skXabNNxqE7Qv1TDizAvSL5gMsUzGMO68+Au5G4sBLon6mBIZ49/J2KQ5SC/
hnlT+vexDYHu9yNriKxwKxHIZMdLys7evSEagjOIcn+fXZxXkjWVo1OthP5zzRBPBXkBZTGy0XG2
h2ofZKqFPOlwWv+vFc4GaBWRyZDC/llKSUcKhKMx4iWQQue+rcxojw8U6y+tThLR3n/dCsTdO8Zt
rEGwyutwlCJNob4AiAtESAgvtQ+Qx7SZ1aaoCvtweBXauQgUtDMRDbMVsxVRMqXABGrmIm/QPCzz
vQMFXV8DZtBxq7sG+sMS2N+D6755yH4atDwcWQDCmP53W+p9uMTLhqkPv90tInqdDmLFhjkDRuwM
M9plTmDK0Dba5ACgQqPOcnNnfLa6e1cpwd7yocC4YWveSTeCiuw/C8pR0Lb4JZ/AbodclK4EFo50
jHdbmAz04r9hIuqGMpfQBljBywjXorS5xr5H5DQaocGMLATgLuAcrTCDaVdYp3knemqqtvoIwafG
QYMTf/yGcdeRAiWn1qySmMABdnv16Nu9Pm4ffInLXdw8LDUP9PJxg0x+8EV3rsG6z59Ql70hcE2B
HcJ79F0btEBAjSRz2h3G/XQLo+IgVBOzF/ioV1iXX860zjdug6Po8mM3RFlz6X0CoQkcjh0vvON4
Y1RkNEeyvmLNuRCMeJm37iG2OxtMWYnLZO8OKOSm3zzhYOeImgpROLHy3uWycRB17q8F545dQOuG
jAf9zF7bXC55qqsgwMhsBlB8emDJt0VkoLJ0OmrjzSUqC07RkMMtN23N/fgjUn8ZDPFca4Mx3tAi
tB94Z51KatLqMEu7IICO4Naj7AOBTNMLKAjoCn14TvCJSBVjfQhb05/xDskO+HhsfHVicwnL0Inw
E3lFH1KLEflzzurZYToMW3kParxysqnOROtpNdq/+vPpOApnAtvURDzw1dkh4v73afcr5TVKFrhx
kwh9rUVIEYvdL31bx2W0voodmznyABFXrnPhzCmvUkjRbFdCUD3MWTMLGxbI8xktknIbiS3DxHEx
yRfNGLZ2A+pU+V2hjQct8//Pr5npJgyShbETvnEi6LsrsN0f5qwuLaCFSAbqThvk2PFLxEs5PNAZ
x1PtLv1yqUutsQrxc14ceyTMv0eVvegFN3cB0/6WYC4gBsDTGEIacenSi/mVFORxkBKW+ZFhvi4E
cnUvWKBU89SUATnQSI4R2oHX2qkzJcezZzoDBKnPwC+AvO8nv4cQ3kztxesAuR4tX5GyLFm7qpf1
0Q7BgF1Qjl6p2jULt2PYr2kbIG3V/dwfzIZ/Y08HJHtZEONF3vmdSNmqdSRip9G+qGTRTvnRTPdO
3GP09MmmPudq/dunYW3CqYl1Q6KrN0aXG5O5I/pw2PCJFLJJlA9nuWYVFJr9eCGp3E59jjp1DpLw
GIsG8WS9Da+enHwfJCWkC+ExwVVFCMCUMy2VWan43uMijpk27bJ/WtckaUrwrSn6O0Q5diI3a4CA
WcArFgaFWARTViqt3nQ+9nQc8E8HtysPtBWSP3FiStFi5Lb1NbeFs6JVuaYt/FDNzWRAn8WlyIGB
5DcFLWV3qGr5z5B2AUFW54KHESf75s+KvgBFF0nI/EXphEt6jPu46+4oClJkfzAGKYAZG/VgtF/3
CnYuyqEiU04FUgwiEu+xgfIA+XRByYNGmHiTSD+3Q9fNtdKm1NAsSZOLr5PqIqTiCndsRszy5Qli
G4RIAiL5lFTNd08Q0fWjAWD7WpSsJ5u25Lec9eQI0qwmLpeZoX28Kj8+akUWhYULHmY46Pk+oUrQ
nxwX51/Xaegnx4zaZcDJ3koTWh7LMDC3N/tOQlu0MHrFXyyVNDbKrQTa7wNLt4BbIzz/m5EmDXUs
kipY7TXEUWo91TprvOdNrJc4yFcKcR4hjV7GbUBMn7mrPaAG+Q2rVS3TSBUsENVcicBmxxKPfaML
3KeQskEPJ2seuoTlcgba2qf2XtDz8ilsKBEbHvCqYQEwo9dugQqQZ+/whN7BPFbX1iJcflO8Cj4S
yEGaQXT8Hkj1quaeREfMtlhB7CxuPHAdx8tJJP+Q+BYoVcj03aK9gnkbXbARyF0+M9BvEumYsPKM
UERk9H0Y/wiV6V9Aj9F9nKLTWBTCJEorNZKFeAgiJUkMlanjQmJhojz1xEd8wj63qOgJxsCkOliU
udkIX629nV9eFCDi69JHtl4UXB7uboI6xU4fC8+KpiqsYSC1iTyiNb1y4JmHYm5LgQEmjk3qax2O
SzgS3Vlj9GlaqQHZaQkPwUl8TDXmTKU0TUImU9vT7A0NO1I10eF7deexz+YiRMeOUo5tw2K7KMP0
sh6K2p03UZwWy8UTJ0cxH7AqdEIl/kq70PMQquWu7Jc3LGl0MQSBErpZ6yfj3z8tDNl1mI3zTD55
5vvbJvLnai1EOJ1DGP2fmx0xPRzG9dsSapuFWM8xTS3NnE1/jWTVwjAmQsSPF6efzncvNq3+iOoi
o2BKQ153KItlrO6ngJy96Z5aVeDyiPoDv06/GHe85Od7AuY2oFavcWloNLAi1np03KM1dZR1wsm9
FYm+CTPIZa4MuIWTIH3EVrfkiBHp7wAuFZNwXT/9OT2scgnl2A7Sg2pIQF8MaMVnucAtOHMK2Nft
zeq1HpCbcK9f3/4+8gLa/A6x6uFHaQi2JhovNlyQNDocucR4z4wsDBB89CSpOKCJTN64Eu1dm//s
ibPnTLk+mg2dhxDiQJc2uf2ZClOACOVnEmqV+NlyZ+LQeqO9sU345tpX2fTCAKZnCxi5vM/zxIJ6
BpSlUksGiqYglJdz9HFERVDa/d9ZrY4YbgAEh3gFBoD8DkpGi5GUWppjnPYVWPwxR2FY3ktSPrhc
ZqpzjALF5y2hWTstS7M1+Lw7eUmP7cLMrRl71CODeZ1LwFcQsqi4JiVhlt7WKgUjZltY1kUWbRWP
eEJIwMhJdpjhRb3PYv1M3EDtNYyBXelbC8qMNZLNNe0VGMYbWuD1JoggngD9z3gsLdqa1ugENHHI
uP7cQztOO8QkWxtikji9G7g9nwLuOjUbktklHTsD4E72DOvFbNW9tL6gYYD7P77T3HFrEA9XzIM+
BOpX81EAUxaO6/0nfoWVY/xujHl9pfzFYN9FX4axYvCfpTK3ZIpSfuFSag2LwibRROZNbPUejmZx
Qc7ZozDVnXFIWP2iL8+CjBD/CkHN0L8RN91RLU7uGdJc7ZJCESoDDp2q7hPy1x2J8aeeMydxiS+7
lh5crRjSDKYWtTFZxRDGSXVnieaF75ggMprtmsc7CsCr4eUewwuOFPpZVK5ZkR3KF7Yt2DO78Ql6
0C0zkf7Yts/TGHazkOqG51WyPZVp0odTm/4iEEu4dsbHBjATxiq2WNIloFW7EuqCkvY1etYT9REJ
1O+wWQ6PVh7hRaqJYVVXCL7f4rCgiGe/XOVHuACXAjksYkBSCTa0kSF2U6iwP9oVC/QB94bo/Lpp
05gSk5iyENuvnHtdFqtzLBkTFUEYhpgHjlRlGUPgk65chnAffZ7VIgUMj459vQ8Ixu0j8xywP1cX
z6AK6waUIVgzaX9LB0jqAeHVMKk2IpKkq/7PleuohfRmCQGKQpaH9bRBmtY5UGfAzIW30/eyPz4h
opJk/hKx6Qwk3f5bFC1TSK4xDMJ+0nv3K07PXVE1o1NeIYbJ1k05kNPTwBYWt0YBJUkAnRIvT9Uy
QWXPVL1BupEb/97vs22PouN0PP9KwPMF9J/BMXWpS4ZEDJ7P7hpbLiuVN4iF9Zco2E19RHv2XbkW
gYfifLIu21Uaprp5y6MJMGGkhhEF3ayQUn4b5qHimmRQM/aBGrNH3Kj7ghEGNHalx8Li5BGWjtlc
rNbgtUL1A8///X+WyZyHOpS/LxVw20UYtSf184TSfmvtnvcmOtJDWP6cmY3GE1o4rLLYEljCxbVH
WwgKZ2YLCP3C/wkxK8Zko52IFfcpdGmUTxGT2VFeer/NYkXhUg2xaAVZhzPAZmq4reupSdaRgV6C
10BCdhA0hJh6d/YmtMs+oUd/+2gxdz3RQY8PO3LoLnDGmnARBH1+PESkJzRYvYnawOgYwYzgK/JX
PSG4aR8nvXPxoCUToCtjlFUThn+d8MeXr1GhV2URL17ZZY76IgAd46bEWIhkpPbP54NA0xsCWvsw
hxTyE50U0APq4ZzxXw9fisBXbEaWqaF0KkRE7D8PzNLRYoRxjaACrexOOYMOOW9HdSQiBEOM2IDu
Z+lAW8K6RoO9XaZudhnbPsFsugYjW05KPLwE5V9aWI0ia5fJNDxCGJajQix9jEfowYOO0idATRqd
tj3UmhwtxwSkA+ewFXpBAThiMv5fjRupYf3vDZIKTUVxGOp1/iijJ0j1MD4WiHZ/BQ4LZ/66v+2k
4n4Atfhzbt5LMyQlFsIjTobUV0ZYLLZLQTJ8UoRRZbuCoDi6o+z7cBWZOCNX6DPatOwTyBZoxIZq
VHOml/+8HFxA16YgyFDymElY+b31yYbhrsqUgzvFY8VShnPSU5qVQcoUdJX7n6aeCcshpeVZQQR7
Y7xpzC8Wkoo8B/8vxIAYVV2rKlPy00w1MPXhZkDxfwV6U2dI4vyqAXWYwliqKof+Tbsn88WGzqOh
wirdsWe21Ogf5yA/cFrtpQ+wjEcWSIIvXuD+MkRRll04r2kITj11BE3G5f6GWGGv6sPfoCY6kuxs
eXb56TcwjskJcHZn1oRZkLJzcgf63tTDHhkIzeVjOe/I7c9OWKy02h52qypONbKV2YIRyfmXUeqG
IUEkulklmWhRSKaXhbNll57WCH+6LFp4wU6VerFKsq0BDCh4RHP1D71viJhIebDyGydrAFOdyLPK
lMu/YhOqX5cTxX6+4aBZG5165F5NIIeXIb+SlPWy8rGqpdUitaj2FhIE7zWDEF/U5YkMPkjO0RGR
1tLkO3nAwZjJoNNc1OVchYT9OqWT8EQPL6X5AzjbSBoWDr/5H/yduTSHjTi5n1M5ZHtaojgUO5qS
7COsPTSMcypIOS9+5fNmsBY1rW6SeBoImNvdTtpu+TpcFMbgkegcxdQm3jMnpE3bfcwwKlI8r+WV
LtQk6vYD/rzGoywx+wveV+x5nBN2alo1s9ZaHvJLdY6ywjtWhIiIKR60GxJ1qbyf/320X9lGzFXw
lp6KBndn7zcPj3gyhgPFMhAkag4mQwFDsnxJ0yVjORRXaq2/+KgdQKYndDiYwY5xCMT5VoHSiBXE
YDcZJaBjFhV3qm1SjJZm3z3ihHRm5KvnY42bY7FsHE9pvT8ieBeyOES6Elidr89T+HenOOiNti8z
v3pGPz7xOJtp/3FaawVHkAdnW6n0Jr906nT+avzD+RQfFFcJum2oSRcIwxpTPg49afFOd07A9gxR
usYSI/JGQRq74c9mcNmGtg1XmZARdx2i4U0NLTwq6LCrJDE3jm5hIaLxMKdDYXDVdfv++0iX+2hF
zJC9aZkC4DgtqwLfH4SWJHkumIrsFck2b/ZwkoHbgND2bnQ+2PVWY6gf9dFRXx6XdrNP+Zz9Ub0f
3iVH3AwA5zpsY6ENg87DTGkQKmBfyuk/oROp1gEJuE8YHN55yfVOn40yV8VG8yYvUv1v96ZZ3/QI
Tl5U546X4q/yQY+jLWj6ONnWrI7donGUNempQTntpL3tRpa0lwAblTIbQ80E4u+KSa4NipnXn2Ej
O+fGVBB3YXWvYpsefGwhyM5IVxXqR25oAOtirdQk6luEVbd4xYhu7byH1QyG95+2LsCWi6BUBvjB
KthlrhzWTVFEDHbJDKV+a3QeU6Sfvy0bKe8Y7p4yNJW5sw2tZm001lWE1eKO8nQx/kjFQE9Tpqxc
z4j+a9Zyjpk+ynU11P4ch47ncCZ1A4ys9pR6ybPiBg08RoRUbY72SjpFJPmzu4ZPjiPcdrzrq9mF
qXDjQrO0OcBOwa9E6UPQ7749aq35xCcwbt11Ts+4ZsAwheg3RqohuOaKsLHmnCgX+pbPtfNVXtbh
mMOHESE4sjI6Z/PyzMolg/HLm6SfBFwoIo8xUdBg5KVolIioPcX0zRKm6xdlxoAmcem2gL84HNoe
wTJ+x+0vl4JPkHssfK3/hBa88O9UWTmHQMi0+uOynya3+HiyXi+CxmWhZeonBvq2c2D0mhWwVcmR
KG4PKyE8DOPqze/ard+JBmQpr90j1I8qV3qg2bxAy3lTcaZWjF21vkgSdvN1QhmRM/O9hynR3JWJ
RT0bivZstoum/xQmET2J5FQgaFv9Jn5kVJUXP4L6/oBAJC7RYIxMGQz23Q8hyiyNdeIl4Vynrkb+
yWktcaWcVUCTvw0B3wYdjJHmiCxDz3dSAeck4+R+OfjTTe9cwQEDNeXYillJGvG4SrENdDyPW86b
8izVHJ1PekYHyuXvwc0zUZoLphWksEBFQxRPjdXo5Wo0YWjMXQ8yZY+o5Y2R/eXZvjOdiXMOhgiJ
KMyw3eMxkNLHX9XyQYkqefMwIUhy8yf/cqTfAlTvCDMWxLjPu7RicxhKfOw2gBuujwcMwfaq1T2D
R5zvVsCXkdlfOy0Y+nM8TbRufnizDUmUh6JmMiylqIO9xcA5UH9qUfLG+F/GmR6gu8I2X4xx3Djx
jA9GBHq1NK01G1L5P0r0YjiDWmh1vtdy/54D+t7NJX34CFpAVFjDMtIV4fyD/QZFJqFfnQbHfGoY
Y3Lf29pWHoBtnwuGQK+QTQAxMpa4L15VzsXodJM6lHQz4K8olRi0k330kvj1KCghW1ZaOpFm2LCX
jp4bQrdxvFnoWNvL9q5Kt8ZYXvLgpfDIzu1yrl9hccK4oxs7qEfma1u0wq2hH6NaQwKGoAUcK+HE
cg3LD2GJVdAjZ87g9q6KlkC3Y2A4E0m3T3ORtHxeljnlTYanK9ISsr1gk03euqYoCjwA/fG1JtJ4
lijv6K8x2IXUP2X7mgILIXKnS5DCF8GbK8zz6jzFTvoNlz1W6HiXE8kHqqnx75LwLYa+V+Y98A8g
m+XdVuknHYhmpPEWmG36MrwaL80oMDGjYTlItCZN7GF38BEkUpgsl5X3gmJ0rRgZLmrpMrTIqQFt
4ImFriuONvBEFNkk0JiFDjxLgKZnwilBMgbWtnKYKLeT/UXjfEvOHArpU1E7UDmTiW9AeVspt7Do
Si5+NM14p0JECDimt2bYdrF0hXTx/8qLnlsw+3xcq3ZhDRZpqQ9eRptzcO6wnJcPXUluQxo2khT3
8ocvKYopLdtA1/meZ071hh06yN0KiIxmgjyRLDnnT6gdN5EbqQfchKr/96W+V5xBZpjyBnE1JpMe
Hketa6INdnb0AwUn30DmNz2pY/gEBtlnnUfy25OWie54fnEHYSebFJCQAVX2mjDxR38MVRBZ6RfU
B6xX6hjWAp4Y9Bfyn8mCFxeGzLoXccsZDmLBabDOW7VDBq2J+jrZQ7yxuPeLSGpTuAl836klksuH
PakbHK9h/4la37PBAuK+B9GgIVs2pe4rCxsDrAzENuJxLf9cYNSmCLJQSfjsTijmUt7C5w9Zogo8
XMQxRNXN8TczEEhRvR41cTNgkt/RZ69ouq+gMJ+VRCKLBElVjXfh2deHCFiPzgIzi2d8r6wEddBT
4VGbsdsZPXxJsXt9g1K2B+nCyj/GtQlgIExHPYVckR7coFgHqwN7c0CJ/UogXscn01h/4KO9jPCL
gJXvPox+4Th8R90oK2xLrCpr9FFcI8D+6r8xfXvLdIkIT2Uw72Mvaq6cyEN4OlofohgtjpkUI61M
4Ic2LRFnzhV+/hvfCkGqZq1cqYP6EX2vEoSmZAl72plwTE6R7MWiNXilJjP5xk2Jhng+gLZCXwvO
zJnI1RCsr+/Hw491iJzyhFYdSZ6RQKnlQZ0pFOzrC/oAIcxqEzsGhC5bVDn+NzLBiL/2raKdUhWz
qgnYFr0lUCapbNp7H4Hz+UYtNJJUgdi4JRQqiOIgSRu83UmbPhTlXtytkRsrSPKTRU/Lo07sa3+9
/Igdj3Ea3tnagrh0ZtZu2DzVmFZ60TGxTpnqE/Lk7kvcFuzNN/r+tExqNGJCyCQ3O1LD5+rxEorc
Y/rfS2QuzMregrOZooO9qacb9zRdZtk0OXn9RdB1O6QxO6goocV0QyRqpLjba96+NyTmdwAU+Yw2
kQl3So31xc/b6Z61EpK1XmOh1lyLQt+MD5CbA4NGhbbpt3DScy9bgTi3dCBfm63MXTg+J5Ttg4Pm
ftQBd9/gKGkOOTc2lMeo/pKDILdzp6hvxLapgAn34fRuZI84WGrW1Pn0zAW6zb3BfeHJlRhb6b4W
gq4NF0e3SddejZaK8y79c562L4JbquQy6yXD7T7dLOCd+ZjRH+JmWaEFrkDjHcl4CoNNfGKIlWjv
eIwgmyqiLd4JLOXzXmGC/Q0vCZPzNii3xc/GbTnU3GN3WB78usQYQmD9QS06Sl0GaZQ5CTuRjuEJ
xO4tRT32vzPAyf2dcaoVA8IME4QXCK81Qbz05XH66LP5lFEpbWnYjVbnm1oNJxSH63UJs0wmhtrS
ayVc6af3tRAbuixEw8OTCSvvd91RADi8CZ5/2sC/g64S0O036VlXsHj0RDbJaHqdq/WMvCNYYoRg
E/GoY1/cS9Pz8Io6qKmwq5nW6qILnPsD5SbijO8UR2ErV1znEcrFWmA6+m/5VuYgtStohNxSakIX
NqI6VntqCSc0G0b9SQKPQcT56onmS8ep3z7ll3WSkeOO0z5wsMjZM1Metm0JOcDA2ZttRv4DaK60
HYwVV1DMu0fNZ0ywYZYOF7KKc4D13xEJyjYLrrfk1biJt1yNdiEYs3n91r1ZY9LyOCvprh8Xmihn
yWmDU6cKS8y8K936+tHZ5KqQsxSLO8IOHM73JEC8AMg4IseJTx4sk8Qx/Q7R4PHWWgv3DO3FD/y4
vM0t/3URiFBGqv+dFRnpYcfJ8nrJ8kMO6gHzdBHAPYaXg0QY0eVhYGKwUU+nJeB9h5UAnPj9NH4C
mvnCCPjm7k/lUE/Z9uccjlIS1eLN4oSElyZNyymWvI5GUpEv3Ste9wM5eKKp5aZ3Bfh5R/V4Jtfa
9hqGaqXFHjxNUT5ZeMYAE0HX8IQT+E3gR1fj/4C0/uXQDp01Vlkf+SM8VOuDCmlWyLayKw3xFzwN
imVOy5kK24gKK5HxQAqLsYlOzOCFUCcXL4ongyRLY1zFOXOX6lR30B2zMBZXtIiWgXlPIRfcZONk
3Rd+/LFlQcC+z8CFr7m/5I1GfWQvJAx4CPQlaK1kILlDUlWMuJA1mGXsMyWgcBkH3CJyzeoGS2Ub
2fiHcqUXM0r5Z7dZqCtnK/suPX3ln481OwyjN7yJTOuAtj14rorz1FbFlPKR2a5hSwR5GB17XEjH
dNYbAfB8KXgMfa9cF8oDJQKKh1rSk5zjunq6BbRgo70LRRCorPYhEk/Y/YPZDzeJykvuVYHQ9VLI
Z9h+G8HPkDpnoRuJgU/5313JXr8FPMDlO/97NwWQry+8YHEdTvs/bmftQsiWeMdCsVy7MmrZ8QxW
t0UROa96sL98vVKGWSbsQbyE6l5lnQHlBTWQEIN+vfKZfiS6kMm2Pv1Kiwwmj1SHand7aG4CDZoX
bn4FNyJ5hHqHtmhXnfDhr/XBQO6LOvmKrKkxiVCpdk3UdK5HS+vIdodUco/OcLWXsRnxka1SowpP
0jIHfgxLtDuYpIYsuC+Bui2N/rf+B7gnsJBitGDwbNYvYz/WthnN/HQfDmbUaVP10xI1tJqlO5o2
QIMh5T24b2lM5h2qQHx1oSN7857ATuaJYtH2k3hmQ/L0Wm9gbhqAxchkAd+ggjkdWlFwooZma1r3
DTqbeaW2HtTBtzS9egu/wiqcQR/TzO4e72wpMxzxE7mcVniYceUUDGXrityF5t8M3yeDeiWpdqo9
LHUW1LDWpNrclg7uk3Z8+u2dQXG/ktRn0/fqCyFobayEZeL9lzZR/LcCYe/qc2WpSYlPiP0R8tch
iQr8GnyOzgnwPg8u5MD4IFjHOae0Vuu0aRP1cGQBeIOe7967AglTKSKaJBXcd2gMZDCzuI0k29VA
eVytbwNWDm8BJ5YZcg9PDBYt6EfkqjJwnoX0asgqVZV1aO2eOJvzUoUex8iGVYk7hoKfssGP/5bo
TMLGxFK1YC4dibP07b4e/of0z+A6OmIt8iGLFK5UT/1wSrwuLO/11eWmZ1RaeJt/nGQqpqigV0o+
jMRosSCf+DTAnu0t3JWfyEb+FgUUnCnOQsF9HbUrCOAzPWTcHOcPosjj8v5fbeIdJBpgEq9UXdOT
UaONIV0QdHJVuD3QvZYSTfC8SjAy14Sm8zbNK/4CieRBEqkvwtxV19BvXUPhhvvregg1kL3jeM/p
ybMGVRVfcXVvAN/tBFQ4XvEluUUjugsdHVxoiogX8uyC2vESdAwyfb2CKX80tqsgoyzIyblAOd+v
O+lBioDdNttKz2IleIya6Cs2qV83fdGGuKg4re7VV9v5fndk5pGN+puKKLN9V3QTTHzATPsU9EVQ
A1ICJ7x44drtwDLJEDLSp7lPx7QdzCcMtiWjwSnrGI2qc+HuwvVX3d4SDFRW+4UrbIYIztwoZjWn
Lyc9JaM4nZeRU4CxdutQ6MGmamAYjgN7FxmK0Ei2XVud0EwO8WEKndFePUCG58i1kwWTg6jVkfic
GiisyS14RoHjfpkJtHoOh/tsNezprrXbDx9n4ql1ymYfeiB0xKyVfRJn8C799KsYmACanuZhfySO
oJ6hPR9tTfAs4EvL864Xs9RmAzFkxoVa07p68W4jJbqXBAOFF2z9lQokRr5Lb9fTOvrrfe2Bz/7y
r+H2Z/YvVsxIM5x6KYj5k37z7iNdSGTKwFQVFMH/Vvxe13XhyYamWgCQ1+ZcDjUwxGwuwbieoqiD
eIlAFLt0w+UmQHkj/2JtruiAc6V/lDS7sRaQmgOXJIyE9h+yQynGJ7ydeC9Jivwe52Ztyna6YLlN
FE8yaAt3H0UpQgQ2/tFKacvR26lQj+q5dZaYOmwb4xPz9SwNqhuYCj12uqgBD5mAqX6sAjszb9AN
Pzm7A5x9l9B00SgNNew4RxT3bArnaTG+p4eUI4cNbSJKHu5/7SzgLHFpXss3iVzXAfUbzTYL7n4a
pjfbrX8zWwwERwMPMFXCjBIE+VUT0ueKgQAIoTDrEv3uKOzneKtckPdGSFNy0IdBo3QvkYG/4zwb
kW2PW62+FiI0ZkkQ6uh6nMrl2Wmr7gwkSu9BQcrUfnnROcWfsTmYm9PhqKuqMgNSoEVf8Jy76DVT
OwZQjVRKMr2HdaDxscBszLESyRbleJ/Y1g/QNnzDwm0Lm2yhxdiKNi7B9chuECb9TKeTlFDV4KrK
SD91ce7DjxpE4Mzn8Fl1BqpWrgTjvi3H8Xsjbf8eoyF4o08k0iU0HEU78x/ZNZGWtRvTghxnDpXt
r20ZH1op8IBLnmHpNYA17DoHztfSnY7FAQgGL9Kup6YQ7jMGVORKl1sQwYgnGcveftxqEp0dmF47
mr4wxL+UHHa1FOq9vnYbgH+McEDbRP1Xho63xnX7wdhh0OqI+yXKNJHPm8QuZ2z75GK+7c8n5Q1F
/q9Ry2zQLGf3BxH2YZ0Lf6wgW2hT0fIAgsBqM5zD/DxAUIPThBJIK/Twi0OEy6iMqYKQG84N2V3d
TpWvzzdAQHXAtBMPqvg3bKNGZeHyISpr2ZZkWUOIL5P2d+Sf+pwM9/+M0zCktZKQsmiLMCTKnCrN
cfVAgdLVnSIma7W88C9UW/e+6xIpJ5xsBJp+mZmUyJIQsS3VLcT1NVzQROlZ14Zx1QLLk29ndC8+
zTPWH8QTKHhrYr0V6R2H2GApBBm4ipJf8cJBee2SmzvR9LmGvrElEVBysRqGb58hXk6xex4LVpxl
atrzXXx8SMiFoThSVL7mNlagcPaVvwaAI2rsYbbEekDUAf7nbnd9TIPxjWg8QdJt49hp9EtO/+ct
I0uggXfc5cX33da8TBcCZdgpWx75JvA9Iw6RIa+ut4QvipOfGrY8XBmloryLot9wbTwDHXrwMTwp
s7pVWJyVN7Lv8+i7TtHv5mLfQnyTwgcw7JyHk0AcUjRcvy5Vw8IHE/LccrQcVs7QEk4GgLYQidbQ
WBKqtURt+x4Ype8kRz0I8YAswTdyXYSzeAoucg0K7EF+O7GnC4MPv4TQdW+IMOqudAZCEkqMGe3s
xq7VbZNodSk2BV/kNaCHEe94ylGESr6hcRzf3wx2DHx7nU6N2cvihM+F6AdH3lFrQF9KjCjjpkyk
cYK/WhltTn1e4Xld/oLYdkfzPfGyE5wYrL5Bio6iaHf3N/ZJWEW+9rkJC6WfYBDuEOOEtn3fAW8w
7T+xfOb89ZO4U3pGs3N26p/TBwhLJMe29SktgOtwBwQbdvdhVSt7Fczke8fyLD1zGpcQr15DATYD
bwui5koYCtGLtFK3fLeUHXnac7hqKTFnq3wWWN0FKgZ2HVmNgJzyBB18QfPSF4VvUSjxUUVo9LzT
b9tWRszoM1Y9Yaa+9QM4seXu6wQ7VgAV3uG+gWD+97JS2bfD5dpgqaqGIpBoSLAiq376N++Vcmst
gex8pNMpGr+EboFAYJhAcffkE5buj66bHU/j6AIkJpFL/hx2kLSnlkSWGdWLBZZniQjwahGl/dD7
Q4r3zGsIQeeQTL4XNL+QlhDnsmpjw0Dk7XKlgMpBFzis7sAVuzKBHlooQ0zQnxTcBP+b4hguo7/l
cUPKq4JCaBloLBIC+KpyoMoq1NfyDzcTwXv8rV8wZMevFtKOd0OB5P0KA2fasL1Bb9uP9O/GxPq1
p/Y2UFT6un9S8ale8dheOJ0Od34jjqTWxgVytvr3RyKMIt9JrXrrZlL3UYM1KiDVdrTqX9h1vnDp
i7urhGPKfUKFZyTkUqK6DwOwBiz0BkysqoiS3NDCKor7Ueje6XG5dUcjMmRUNwcJs/JfCFwYEGkn
6DxrbN36xsO4fAdHsoPxpr+L8zA5pqHMJBWQo+vLWc4tSpxEduZOZav/DuZLEhlT5efhXB2myoSx
mGyuOZCM+hTyl4xcvqBMyawDOg61kxHWY0M6ZNLYIxwoyrB1LWHZw0d81MBfYVMdAEsTe/En0g9a
MgFMaaZdXDREK+peD9wOvo3PuS/k3vBKshPdWUg5f8aydpRYjcBv2PK5qrqvIayihmlRY14E1KYe
wZvPP8B8cM+F+RS5wWMy4c/HJ8WNICxt+PzcgHUit3rcj+GKGgDZpj5JeKho5ygo97vna6anBFcx
8HyPuL/WvzwzcCUF20i3SrnW39tXAd7tkiDCiEUIdOGYM4HciLI1KtAyDNQeSo0cuMFLWcMqUiTG
G6LwRGUUyWAWS1IQIoxC/LP47TSHKb7I3kzfrPHjlKLB5tunsNev7sTiHan0MGrCSD8SoE1pGKl5
qPVpTZUHbtaYf3GUKEwLo2RJgySPTUE4Igh6MiZ0N8yvVZzdTlhovOraS/WCSwylA7EoCXNwcnSi
nSpz3tyjItL6ijWIv2H3pB5BY/+Hlnc3sh9IwKUjPgjpwdRQCrKQQkBHDLpR1akOBqDZf67F95RY
sGsinesHT03IIHuNWcXIw6GgrR+++BavuxVswy/rnoWprLI/zwdYIIJFAPvTFQq9DrR9P06fWX11
XEh3S9hLL3wBsny0A1Xup8De6EzBA2GabnCnoKLTrU5imiRLLPvD0YAi3tE23RaDhtDF/nxof2AU
Te6PlTmLRGAbznGjfa09bFGMLRykFg5405oXDXt9G6y1e/Bbxasy9c5374kb8vocS9EpERlfNkUO
ogrohjEd8HacFfCt9Cf8khyPZNjcuu/5vkxvNt5e4LDLdD3jMi7pe8SRx/3AtEB2Sm1uOxstFASs
Z/DIU/+icMvuOgUWldApyDNW6lZu6jOaSpmL8Q5Te5Vb7J1STgmAwNjN4PeKcmZDv+LGT9pMp/Xk
Qbx6u+oiDQYJJWGIZjj/XZwkBnikmtZCDZelVm54TADNtYEQ3mYav7moSAJ19ixpWFo/x0vOGE6b
kI6ofPwJ8DctLkQge9/JuirqVlh2R40pO47wEPvkqdIs94YxyJSuBZhy9ZRKruZEtVtai7kxuF75
Tc4IAtEhkGAlvPlGUDlMe5IsR3Xsv8USPnOGLYuHBxkDF5pkYNXi7QZlb6TgLvw21wsSUHFrdIQA
SgGwnCBXgEk4RRDH5y6XhgJWIyHJzydVL/9fZa7f/PSOgSiuaG5NkC4c3N+swI1AUWhSOjEzyIuR
ERH9Kz/a3J0ZxQRUgt4Mg7ii2UnIhOo/KoaFXaa89asiUZ+2ZGQRX7QcVbTJ+J8q5NXENKTLRDQK
qanwRGobdJNMyqn3GDEJ0Vo64h3F4B0wM1suwVSJmquGf1e5FNi1s4qyzf8/twoxqd5Du5fDpkZ2
9nXP0ou7bo3hZ5dwfuJNFEFukMyaXe2hVbAXHPi0C70xSTuw2fmAfo3ffEiFlstl9+r1PA7OPoXV
S46sDd5malu0PMXwcIGNehG5dWeG5nRkNXvxAynTbk531F4x3eIP+HzpTCnOOXFlmRutK4d7i5bk
ipA9gbIbQPwZrGKYUQ4WYh6NuOuBxLjf+z/WL6XtDJHmbPZPwNwCrYVxW+9JCNvS48qQVLm6ZpdN
TyZvpIc57jJRPHS5RnB8oMI/5fYhHrFECIltK56Se1AUmU5OoY1tzxB3NLSk9mVPz7DVDYkyXF8b
aiN1BUS73Bb6jP+EiJTFIVYLcp0obhcb8os6O9tVSEszdBHczzvlos2IUHAUlGUFQQ3EjX5aFHOe
j5ba6xG5N6APwcRzCoRVDhyzthg+hlND8+TS8lmAk/Y47MIUcAwLT+fvmUKrxvUhgfOEg73XRAmC
ler2tXqpQzNfG9+67Zi32BqFCqeIaxryeimMJAidCrGcP1rOUTz8zorTusVn+tKTdtpfK7K4D+5l
SQvyaOSNYzRMWylxNQhcKG5Pso2E3zdi/du8tvQdEJhkXqtsrr3jWNyldTPxgIPwb3MJMQBfpbZY
CJJUdY2fKlTbSRbYugD6x0+pPQtNSRLddgg8uNOkwHSV+3a4QoRySabYihxKgkUIHCnpuV1d4Uhs
kpxi0lTqDUjYVcWymHhRW+hqETc9Zq8Noo1lOdivwOPLJrpeAB6uOIMqJwMKr7PiQMGg+VTohUIb
v7AVsHhGcx0pifs4u7Ee2gW6aCvga+vD1SCUhZ0H6xMP0jtO2OQ5fOPnFIqT4aWpvpg8h3opdv5P
SsN9liP1tNkcJYNgfw8//MnrNlRohcXcjVhGzyggRhE6dRA3ShVjZg3P/jSrMJT7e59tuIVN2IQ3
UU6kmo9BxqHF96uGt248lOUToHNRATCrfCZDlShvo37ryf85/V+FIpMR5/tKDTIcozFRe9KotXqa
j0BJ8GIMlJkRxKhYF1/sSvat7bjIN+dN4sgp5Ym5vr6BeF7id01qkn9LBes0bYSb9zuC+RWQczhv
SepEA0z0Dl52M81nJCaHC5FEDUTS2ZbbpKGeTpUSZXHbNMzs8u1QrfUA4yqb8xUEVg7kV5VRWwUI
hmKgozLA8c8Rk4wLjwqvVQN22lwZi9RcK1nFpu/+kZgvEJmWNrtYIb4OifL3Dac0gTUE6dbe3aqh
MI2uBIUeu+c+L+rRf4uKeNCYNv5qQRb/qhIhrpDEjZM0skXkfUne3SEPoDcwACvwlv0NrwmHG47I
/SOCxa3BcmOVI9+a0Wp3QUmGoT7bzViKTgGe8xkMHXl3Y1UwY5ygfQCu6OHNIVsDlp/q85qTXtrq
qG4HSxSeUzXwMD6/lABE6DMSLlRzyttRjiBNffOy/58DOUWy1FVmT4FqaRhW+5tko0TLzCFKf9P6
CmMuKCNtegfoLY/IN2GWnIsVSSX4SRTvDYHUqLjpYG4KLRegAnf7bO/U0WhJkmuXNQQDmMRhdEO9
6tTpYgbbBkzb8SwcS3DSDhdB5Mhn1DAGQdwkkrculN1YVadDUNYVybMFcCtwjhzTZl3/L0WMQ203
qO75wrDhr6sYU8XYlIiMk7g4Pw0cUloa5Kw8P1tl7sWGP4J5J5x+4iDgMyjbYxaSac+1qRvsd0aR
WRX2O5CxnLuuaekOfSsE3y2PRAHaGqesAP5R56KqAR+bOz7zDe31FbJiHy0KZWEOZ+hWyYY8EXiK
BfNB6km8Lca5YJLC8GZKa1eX5yWu4SxhlXrxbMa2UjFSa7sSf6d0Qd61Ss+6T9Oeae7OinSDWzlC
2CY62N5dr0buOdtg/XW8hGsRt77GNWGr8nzQUqDoQ3+srbTV2uE2HSYlGJpOdVeCNmVzIRFPEMX0
0fEbLEjldeiS4vSpt/ygv7Le32tneApFyBoexY4BDx1j2LEbPrBJdOd/XBYg6qViyeLfayzfgaUZ
SwI1iAyFE7LOntPdc5VXr2sgaCdIsIjvH02haMJMm736Eh9UnI4FpgX2FIqCCWSIK7ZgyxfgU8Qb
pKfaloif5xAEGMTBiRjOmqukfrvnpedcx3kc1UBBbfxpcSwIz5mBTEMe1oo78zp7UWm68Qi2EzRN
ayxplCiQi2Bw/XwfZf89bHbFAiAjNayMKyOyYFSzd4DwTSgnGvciQi8Y83NcQQNJ/jHIWtK47V1s
836R26tS/L8A9BAhfHHMGSJfdlDAzmkmtrWTFZJSCKIl+F49Ol9ex+xFYhDJOq0oJaXchaM6FHNc
X9DdtcLXAzJT/uKwtpDigYYLZdhOGSY+i3ck7Z6ONApPgsy5MaCnKHwKdNp3hNJobUUDIoz+uHjd
3Cq3wnmeihFBUfOTWwkZxeD1rjZZDb4Mke0PmA5HGSioOinwl7c665Vwb7mRNPQHnUtOc92P2OVM
TAVNyMECZ1zixQq1ihMP5TzKO/4MAO/vLqttl2Z1apflTHXDskhWMlR9GxKq6eETW1Y4YXk/U1Yh
OoumGQsyA1uBIrpy31vKsoHuOcAohIQ3PBAN0WDFlsI9tH2fHIE3R6p5Em1RqwGAty1/bnhXkaAB
5tPYLIKw9uRom8JVzMPrrqsvrvQKe2rgHRiPgeT/95NHgeqylBedMy/JBsAKVwMQPrg/HyoPQwIG
7soYCPDHOq8Kk3Me2cAEvuuCcN478PQkq2bMJm0q4LrXJcaRHK9LIT6B7xj5vMqUAw1g8ukv20D2
R0k/e+lgGC6cvAiUslfp+pTTREBkCTfEtcKLvhjf9hC/T6LNsreyt5P89I5iTsZ1LFL4EATyBXlZ
M4HfCpHcdewJeS4z06vXc+tlij+jOisepCAOOR3MQW9xAevKu9z9/LC37KBsHN9HKh4Z8gqzA8Fh
3Kh4G0CFXmZATGmd0jgcBdMyasbYXdP2W99YJ9quzA+5RwucsKz+aWF7VlwY5jhKseL72EyvcfQR
vEHB035eqfQz8YWfebtcfkq3Un2gmNGomy0g0iDNN77xi8VVXmjDN09gKWMyu8eK0v7riAeHwPt4
4JJlrgobxhXBMMPuuuoILEcH1UhlnO3ON+v36WnI41eqi2r8KvX1N1ZtgFL1Cz4/IlXlRXZ9beMa
sbHY+MZD8mNF0lORnXyeKBUUowbtGgIklPOq2pe7tCnjLNizshOpONpedmdFaQGl7vjZrUYUNBLw
6RFg0tLwfi3in3xfI3rS9LAADvK0ZenwfdycBwTMgBcudeurqQNSpa1pbgjpN12AzXk+ghpWQUKw
lgXAmZceuwqT5ftoI5Mzue2FK/OJ/In7QBg6vvVti05fi6G2igMmtMIksVpBiV1sl/7X+b/0mJXe
KRG7gOGfCoj4NXCTdUw6lsjCCW+iFoCKuwT6kvmZlKpNFROcRmc+tHmhbsURO/+IYHpzgLiUkR4C
Sh87WKZMXHO6rmmtkTMnHpZN2vZ+7XBhc7PnWR8nPF9qULgiyr+h62Y45zO0frcE43gsUZwjLt3f
2dEtklgDLHAMWcxVqshQK//ijVAKdSj/2bZjFvSD5nLzAl9mYnYPSomvhHnxFdip5g3RC1z2UfCy
0qSbfArbnIaEI5qU3wkfp7tIresLDTTQshu3CgM6egG1gUOgUOyZl69eBYwY8K3Mva0qA1RSwMiU
jDVAjIv6bqbT1KvYCE8ICrbVDQG8FnEtZtM3KlEZC2sPAao5gVm06Ao9pmPrpaKHEFFpc8v6HH5f
DR/kJ62apDzIJT+KF9VyJK5ZUZsVqGd2XUNQBL6BCh7a7jRemf1ItR2xj3CbcfwT2UlMAd/tEaGy
m1Ji7Cu3wszY8zZHO5wsPZ/jqtKH3QnwfOXBC0PrZ+fphm2ihxUgWHlVFJvaJZPpTqiG+sGOHYkk
W598wXQV+zP8TZujrRxBt5AYqozpfv/O99foecnG0/6s8XmDJAjootuJk6NuwLxZazJ63f7PN1Vt
yIatoiYGEhsFVTcW55fZFy7F28ahFJ5cn6BkOvk2j0WhaKmiR+bmc3tHrM9uVPBgyfO9TvOTJBz4
LjCD+YkFK9rW/aQpef+KL7+5ei56zo5YLuYo6AcaOe5hlw7VWcZj89+mLmfg8tmcTmo4zzM3ceol
4U5eIos3Wu6sHC+pD+kXMWPDkDPInHHRviCkOpnT4TQj6IaiSuCfLmIsFBOyatPTBA154SmmwlQ7
IPpmuWTIKK0lKEUSkm47H/0Xpr44qg11hSbpJbqxvCfsg1yc5xxcDN+/wzSEfAmkDtRfE7PmHxFb
W8D92pDj7pMA5cQNF7KZqWhP+i8DSZJK2tiEphdspzVXM2K4zZ+1AeNsljVJomX5ms9WZdJGNoFG
5lUeY6CttfDKbJ6XVySUX2piHw57o7SEP/i4WmPPL/3IUqO94mkIf7QUGx4FZwdaeP2CB0n5qflx
K01/zCNcjX7p8QJTJ2OTzQKHFPXdKSO5k+P3frVuS6hPYEtgq5TIbIWKOGtt9HCjWgU4z1glNVcF
G6JavfAnkEal+EE8iQ0YgDdY5y5NMw77goN2QPWUXj6AK6mfSQ7FLzDtBKb7pOcMqCBEzGAjnMp5
SrQUIslX12AGa9u/Vm968z/I5C1icTLgQmIUQ08+JguUbNayu5pX25Paouzesq4+sDS4ev7WtDbY
8Wtjb69Vh6tbkAy4N+k33cLAiXKp7VcDk3KBq4agtieaIxikNbPxCwyR3JeKfe3EsarRIDsAXmJn
GTGGdep2NRxQEWYTd3XdvyeBNh1rurAIEzSz8sA7/sddEIfB9Dm2uqHLZT123CVPjU1x0iTH32Le
3DL9Vbbj3lebeC5ClfuP7m/NlUlptEsYc4QpISkrHCMsPp9I0iSi8gLWa7lHVlEucPTytpiwJrKJ
q4KUSKX3ep0VQQSkGZWBwZBKhd54lCfHvMuww42QQyGbGJbkzisFTGr+ggAYnE59NN0mjgEgZPWB
gvKj805wapPBj+pb9KXotguPALUPWZ4JSqveJ/OI06Gihk4DvQdInodW90xi1oEI5fzq29CXKCcp
WQJl2jRjZpn87NAn0s28Caqx60ytz6fJZtBxz77EkWOQ6jKfEd8lVVFCoTqerS9ajmSbctcoqVQU
jXn0/+65EHUrabaj2+JJhpHpu4IXQO6fgJ3RmSyn5G0VvhlySdrp7GLE4xQiyu//N041pFT37E+I
36CW9kbx/Y7UCB2ZoEv21MQFfD9smZY4AG7IjbfIpdlMRf44/8CDK+LG+ZKcJtiVnUcAPA0Qr3GT
h7+vPCIVdGNEp6TuAqhV1Xq6yr1YaGq2W5gtxZ3DOouCNNSUT3oJcPcFjiCX9g7gLLf1KiOAnXRG
pqwr9Nxdesikr2OZABGcKAOBGtHNFeOX5t277frGOzAL0rCpaxnPpm4dA+G1z0wngaNlJ0wbOQ9H
sLNjGU0RF6ESeRVNoccW910XQ0BV/D0Aoot3iDED6251Sc7zilVk+w4/wVQ869+JlgQLP1sbfjg3
2iV97gvxrl15lJpES7JAe0WGq/TO5OG+V1CMhxCbPzKRdfPVwO0QPvaVRmJP8ZFqvW+gl6EQXjqP
xHEWDQ//fCCl5jugXuZ2S7lyRN1tQ+nvz2Fmte2wfktsZyNWGTF6DfxduLrpLWd8LxaXdwD1IaEI
7ndEFn+43aR1xlltfY/oHXCWeXLP9VPaCgRQE76AJeTRHqPmPfP27/w7kws+8DXVk/8gnFoEBrXw
cBssWOY6z+/N8bxTQNf/H93a3NgQSQ80kEkoMWuqV7glMXU2AjlxUGrXQKn/SG4zChzqjmsGaGrZ
y9t4ycrc6TOvBFgIwtBhB7uMAQPoj6fQN2tip359av9h4xDBkc9300CsR06r4kuYpF2ZeLoBc2Qj
lnMhn7VJ25/9j5EzRW9VldHGFeLpo0l86AZ1t4v3B2gXSO/wTwfxAzHGcS0keRhGtYW9lZW+ie8Q
nl3dhcDq7NbxaSma0aorgiM9k6Nf0x/CCI9o2KoJ0YIMPpUtLTiGQDH9apzUw4EawZViXNPfcEbd
B6pHW0DR8Ar6NTqPkiW5VpYW3TjTOugpsjG2x29VgeNJCB9kGY4K3WERoBRzxBMaMjq+M46sa6vs
lztQXP0fl43ubdrE2LzqXtl8W9QQrIZrYLaQ3e52yJ9/SpRVtz7cK5ovVZmNoKDtIoTRd1xP5pe3
aQJQcpnpuuQNaulo0qiM9RlgFec659le2OOVR3OXhDtLYAZT84sv1Jjymn4UJaYA80xGhcbiENOf
qmYfgPQLB85Nuo3KzFceFWjjg9OOLdJpPD8hNU9t4XwFdt3NgFHAVvN1+5r1KWoy0+5PMR9QE5nF
AzP0tkLopTC4n6jj0p9hjpeYFBW4Do9k+inHbjPJ5JpigvDPW0zZB0liQIXQvNhtaDxX5T8pavMt
PJUvARCX1pgpTYQAcTkSKKCApOiPtv9FY5ueWOdCBqpO0CRgSWazImHDm4RmoLpz3lIxdJZgbC6z
95r1a7/A2XlHVNwt4b5Md6SRy8FK6hQwgedJIJPqyhCnDFIIxXE4rUZJgUOocrKN3LlqeNE1kSFp
8326N9lbSXiOo1I/v566q3zWJeL5MG4q0BVYJMc30rq/Jf5MzjBvkG2kH6Au3EbfTIddJmB6w9bI
1u1NoA0Ys1byfbj4uIxpA1yeG/v9nmGmi8gnxfNZc8uUWRUc8n6gtuB01ZfJSiTmzofacV8mybzi
N24ZO+bMFagZSYD8CHb/nK64h9o3K95THxTkaRG7cWB7wlJxaaMlDwdZI7z38WDN7AJyO7vDxqI6
ed+2rZynhi+/unQprjllHQbns8x32yPUKidZ/t/JiNR+BxKrvnza9rEg6OhnurOi2f5EY8ukhOrw
rQw8Z/UAuZfz7Mt5GJkAJlUONY+p+mOr4hEZX2UeT7AOXBVs91OuMkhlUvZG3yCB68lVMALgKlCU
tLmxxtFeicmxtOUSekJtn/PkwtYPtvJsLUoqqCNpOrjN9l+zdtoa61sWfBob/ecvYnG9qPFV6FBk
7EhFldby9KKHmz+9PUzXuW1wcobMjo+r42fCqZJNKnOP/rwwpxcZQGabpOQyDGhDW4x9ddQCInWf
v3tHkvrdwb70ksrfGvB5hfI7vb0nfkFT27+9IAZV9PmLrj4I/bdjlldIjbQJ5Ff0C0mxdsbzSQxG
Yo17XAQsnwb3Hb66G+6KxnPw946QK4HsrjjF1Rud31EGDAQfvZ4tv6liCcGZMAfHd1AsqZbOaIZQ
NrdfceIuqJEcnOUby0Z7FOQEAWUxKabi7ZjLEC6xp3EoSkYqFtw884iW63tsy+rr/WLzrrrrHl6U
zIZT6uP4UGWeCnfe8KVNbvZ2E+rXf9W6nhL+xvvI8aZ+TksSpjjmOdTaPMBeZQiBlzJmcUS5AYfi
PLSug9uxEGAlMYCsVVxH3+V1oHLAaYfkFNadNeqlJ0wIlNHLa2a3e9sRDFv40npTuwRH5Dy7DhQg
5+g5fZ/z96F5GszchUgzGdRkyvSpTWiNwSoG39F8XrxI/nLwcNKLkp3X1CCsEt4ZpENsKrp84NXJ
IOy38NdVSgq85d6skukjKEw7m5G+r00NnD6U3LzPjvXNkEoV4KjdPA264dge2lbZxkTRq7e1CIbk
wKmBdtLMKjbBGE+4bQuaZ0clmJk7kDQklFQy9Ng7jUb0uPzfIgNuFaVgFZTAQ1LvmJcf6oT+ChqP
oG8rNrH21gs2Qz/xjL6YPPmTqKy0bazBiDM9ez/jK/S4DE3rCdyugvrj7KSjbEt/BIVQZwcUoXPz
PNa/+53Dc9yFmf1S/5BiYsye1QrQ0TB8hi1dZ8TII40qMKHb9tMIUZwUkvrdBIU5GmfCGmyaevMl
xiY0B+0S+cSHmz/IPzUP0hKa8HEtNe5PsPYdFaVKwRJ2KMwOiq+89D+NOHvgLXWJyPuqM5171t/g
7Zb2NoWfAS73Dxs4YHU8CR0wLE5o4QURxkL/n+q6KRYu07d6Q8ePRlWIWQMHaF6Dx8w8OIgYB9Vu
O5KwGlrdZRdiC2mjZe5LCboyCvQt3l0h6M8n/DDriblojHpbTFFvgMLJ0nWqJSvdRYXcqvT12c6Z
JPBK8sT0CA9wLzPBspOBLqcbCiTQrrf6XrdBA7QJH/rNIStALjafe4exXyH1x3PZcXljzqqeKN/X
T4BnbHMJDemcBi6XpFA+Kw59e63agDAC3/kQ9g23shNZCvRwXdIcufrWyOBR2sJXjaFFN11cCr/f
eg2zoArx+yFD2MxdmV1KEy0rIHtvLm/BwI82FABi0E6uF8+Ko/lyYvpy6kquNgbtWcXeAle5ogUx
APWNd5nda3MmdEodBHuijBhspqs0fzzvbNQxFht9PeAHs7nPjzhyd2e7OwbwSo3bjMv6/3IOLNdm
XVMH1PIe2ciN9WeZ6eTITlGlFEPhs40BN8pDcLOxCqLsRRLCO9OCbvyf0N8iB4s12RBDQWpV3nGF
hXwgNmSN4u9ep26bydhhiK1Z0iLsHFt5cjJtEqg7lwlJY5X763hp2vg+KtPFWASam1ga5vAl3Ttj
HAZRRO+YOyeNHX+ShrPUYqn9KiOh7BcCj/HzA08XWuHnXLDPeMe2lqRwOC1GnU//3QCtIO7idYXP
Z4cZSL7mmltIjn/4hifmrPpUOEA5HmKFY/o/VV+hZlFcPzF6fuG1EvJZSZozd6rlCMs+0dZevhjf
ZTlO8ihpNWzmwamcBmUFPPLnLWYO+/opqPL9Ba49jgkAOMcxCq/rBIYu9VrcpJF5aUGgR2J6taEW
ZihBt8qUvX7A3we/I6MxCrgeEKNBaXDd4w1M5mVj+lBGpCm/Sgdbe8Wcs3KPWFOnPn+hDOqSyZWY
i21WBtc6byeLl+0fm5lnSyg+zD8AYDOstUVEyycNb7y+Q4Hyw3D2GbIH8KYnrh+K1mEhhv7MqJBa
n0oN4moifBSmtFauPvFVZh+Pz4zUXMSYm6PaYnaW7Rm6FEhdWvI7h7e3sJxvrCuF6NBzhEA1qpXN
AthJEmpUWhDCJwj97DWCtwXUmB0Hhdj+8cucsRHYNBVUefv74hdKITxpBFNn1HZPj/5w9MpSmLjL
gTMRYeDbHRZoYVTP+O1cALphfdi3APMp47ukSC4PNkx25AGwrYXVR3UpZaqu9xElqX1SpaG0Ii2a
7dK3F5Zj6LHf8TCTRdbLuGI0SJ46wM0YuUD+YbWrx/xM2vSQKq4yHJE6LsX+XETdznF+pJl70noc
e+i99RAU9ROt+PM+HSPM0Js/DEe6wH8G+kzWMyP4sbi82SmfAfzysgg30NZzYB/RLhFoBgm+4fc8
/iGrH2Kpm2Yj6FwiFQFwBH/VRz2jX0+K9LD+w7eWnBEt7XSbaxyLZWBIDmUdYnBhdgJg72X5gDS/
SFYUgunU2EQx6so1iyTKDyvyKEsLxf/D65nn6mf4WtuOq9lNDbFsNHn6q74asM/aMEftj2Pl5SzI
eGo+jEMaq94D7M2cbOXEY3fwn2wjUDimX3fOhkxNw/POQr7vLcajekVr0UhIngiUZyywPmgikbGT
/NmHXv5i9fg0PUaA/6JW0zlE5lraG1Qtz6eBNVI757s156tQyfELkfG6H4JfS8Trhk8fpcQPlrd2
mnhpxhhD9GnTXTJNv7xXX51PSiNnLKT3IU6hLe/0+nMpccb7Ub4isXw6DdYuYZMkV1NVkh4tugy/
XhWffJWeJPK38n4XiFM12ZmnfD9M+xQrXG0hXB7/fRuYRPe0DV8i+UPqyALPLOI93K/B8h1nYWs6
m8Vog+OFPxkiMMtk61OBD86uZR9KHbKYxGNBHEKYPu9WgLP6MivFuVokV0Py/5I+o6p5LrjaBBWp
Tm1B9L9vQ23QY3MgYTLzfHeAbuBZP1fJPy1s51ILZeYDpy7iyOi7fmb4Em2kZq2wlFyo1+U8wdIk
9vdKYnHWnfTpLDKNhlK0xcFN5aGIRVcVgvWzAdbH1YkOPvZGd3f/jQBtKUTgxbX5aGHbnYCtLMCc
4dgzmWmALT2e5jFN+gIZ0G84yOBo9BctBJwXsHZ/BpU6Wdg5wPp4KahC3CEcmGSY1oByHAmN5vZO
VCk0M2OtyP9M1XlNMR4saWjTV6fZi3GPU2pCIFjMh+QIt/ZCza++sGywrQyrLmkyNAwZFOgtxqkp
LPg14ADUnDjUJzCGEdIefXL7x9mp7sMypgfCtafnudmXII98INVnDB3HYJNH8hYJ+/bAfDTXPXfL
RUsTVHf1AcwWT9Xc+LKCHRhR6usYA/lwdPw3sZflngyOlkxHpzA2fCl3OnayUKPwue5MK7YjkVKY
4nhdt9v++6woyb89rW+9xCmVMou2mmoLpt+bwj3aDtXclZVPGWBaDSrje82l8TV1AOVhPSQWtde3
bDlrQ+TF2ZSefTku2eQBZEY3pNiKSpCi6tBF1UOs6yiofnCdR2fExADo1HoUr5xu7oA47BPuia/I
hgmRfbEnTYJcgGYu+OknX+zhm3nvv5m8XFmA9bx8q4PPbiUordMKeOx8XyO7Dz6Ld5jMTQVPLawz
y2CRS61YWtz5fDWLzhpWqjarSVxFkQlkZey6OD06Mv6jEW8m9alWybGcOFM/gbmgFFWOJ4JfGz2a
ta0e2SN/WdAtYa9zbCIM0fiMm3bHO7yPKIsprNkBjfmBbe2Gz5Xc0Fw5g4wDAA1Z95FTj5/aqXXE
yZSgWX7ernE5gEE+GU1OkatVPRgIoSeE+Jmw7+UmgYg/K0nL7PcpCEZPPlZj5XQS595lkw4tiq4w
taZs0OhjVaSfST4lBFyfTH4K7fROn82MAWINtwReQmMnqwrngLRky/eW3Of900mB8I8JvOm8cpRJ
OS9K8RNMWs6TKUpOd+Lug0SWMwoTjZ6bteqhgnGw1j8RD+Wyny6v2Lad7C4UVIvugE0jq66CWPOD
DGe3WxrYjPKlYPTyek6ko6cJyogYUw/VhR1mbxBhK6PoNWVrcdWx1iAnmPsRoxEeuMvDpD5FThay
bxNT4jtZjn1k0bcrxru1y8lJQ99UAuLptMEaOaPCInlx2hvgcfKkwIy+QohiyC2fgMmSMGm1utMj
FIV5mRlUahX7w88wuK1yOedw5ZD2n9+sPVLb4H3izTfx0nGqK40Fe1ye/R3lmwoCW29SzkCT+bH+
NK5IbzmVntD3mgSkLkvF//W19NCLhKgNhRFE2SCLwU50e9rF3F6yVwqDZceEcYkDTf8y5a8IcVTf
AhKOKewYa5NbvwM1CusLqV6d3kJbaV7KEgKzLaCtJo/spJR8yYjWGHyXcsm4GLDDugDJTkdmrCef
SkldlGovWaa1dJJCCnF6VGdLkQ2mDBRQ8FCppBalC/bjfwD7BgBa9HdRvfQ8I4UsZKjoIaptnNHD
fKi3sBPpYgmHV953VPHdruQ3tNExRRQRsUdwdNUSqPnstMJ037nRCZjYIYCK6DfLgxj9QXUaSqkJ
a979THqE4g2iWLRda1nm4bdDrzL5YKCQjOgrvrVE4hqR6ht8dN3VuO0DOysGwG+kwyW6Y7fl+rA5
8IDC55Y10XDOi7TqzZnogsmKftofdzzLgoR1Nv/h7UHVtCCrUkpVTwS4DNzBGag6nsGeN+NpqJ3t
NGw3x5pAI8hi1NEhWMliaEBYi7cFVlc71Aog/I7BXXf4Zv/TMqpU8M1WySoliuqayBV7Ri1lipXt
iTtVDLQXVkvZ+wGyU4MbogP9LZFgi3rIkvKuZRDZQvqMZ/r1Tj+W/KUCjv7oloLMgpQ8gfbOyYKw
IDFTfuZ18pPRtOUiInZAqMw5CgklE9/8XxXTVI9lssp58Mm4m1AaXSG+5oFWZIncdNxIM/zpjzEI
Jadi7MgVlKIakhoY99on3OMFs4L7LYRatLHAgdYoqrSSg5+Qq21D70ZAY3oqdm6RuK4x8CqbtJ8w
br3qxm92EyYrg+Qv+p8KILaD3EACvT7RsQaXGQI3T6EqdPNrBXAeWT+HI1M2AZotFub7mxR+yyE8
W1AfDg3zwXQtnwPd4Fp41Z6U4CTT8ni38GlfvN3om8wU1+UnBffVNU3T9MAvfp+eRRAbrw+pv7P1
VYR+FmpcCNOWcecucOahGXNTijJEl6vFXu4kOYrUoTOzclIaGxv/EU+bot6N6DswEIK1ekZDJBEx
KkBXEQ7J48TMyi2OXVCc5SdKvCZuE32GKeLAzV+j6+Y9bxag2q7GoCPvYL83/VXFivKARXetgE23
oHPSi+qSG0MR13XoD5PstnsutfEo6xvsSa3sFv9kQ696p330XoCxi2zuNNRpGT7Yu2o8q/tE8/MF
3c1YfTFh9SwIseKjQbjQyJqvwtdI3koEYaxRymQ8ZXLSgOlXewuhBt0dHoOw1yuAmD4ZCPl7Lkdf
VPqEOh80y4UicSfpW1jDZcBfA4Tut8rWVNC1JzCT6f6FydQvMNoDwr+bcH+tvVrtGRQJnTD05KBl
WIf7k2fDBppPWLvAlnGZnbE4HcMoMEPL9Bh8TB4un5jvTZVpA4T2l4wrfZ9GDoqJHC1/cAUunu8s
+M0Ka2wX3Kq6wFzqIgnwfqZBQHRtJavB8wf9xaVtW37CoL94EhsPEPCQZsM9dAFGK6g4QmdClf0Y
E6yHEiG/h94bpMdqcznblgij9MPDS3Y7w/SdZIEpsyNPNiYL5d+jbU+BJpA8utDrFHRKiauL40TK
ane9xQF+6060uUzPbSh1c+TsttckM/KK/YJIjKLPwWynvVlBMKDJivLEKbS5+yYlfkYE6YOXMszP
gwtRXcm2MUtxdBi5swBmp08c5YUshuadJoKcZi96li4ep+YrePd15s88d2J6oZAMZdix9YnJ6PcD
Ql52ikW1ORDS8rAuUi/Ue+ROcnqz/xyu6hv+OlJRcTlnAUxR4nI8CoGxmp4NkeIw+DaPFyp1b1tR
okgFE0s+wsx/oouWlre714I2GYqHb8lN2RKl4ue4erTCdh5OfgDU87wMJ0eDyI/fwwW+KhLP0TR3
ZvIfNDUxxZJbD5D/5SalO0hXCnXoAcvwgPUsAHm6qMCAUSsr1YGZbzUCpwpgGgvSFJmAtLSxKn7u
v9oiSYTcTAUtt9aToob4weayupqp2mahg2vbSUM5MHVZXOQNNDPKP9/wIRYDXZAp3UJ0a6EgWmwf
nxvwY/JEPS1adwZORdZ4Qv82SQNk4S6sREEdJ/oLd6n3aPOHiedth6/n8ZbqqOKGoBMVzncxFLz9
iZYWQmzrctt8GIGjFjziRVUTTmUq2q6O20SLFUJ3EOmHCZ68ZxcS3hD7BIh54udi3Mme/jtiE8Nt
jLJdP/JBmUVKKFum2ZT/beQ0R86lCqPzLgDCIsQpyraxLvE2jV+9bLBBCPTxAdBfPhNssmGPKy0D
SznnVI/X5FECvfDD8AchMpCv4iCi2fJg9x4S1QrRELPjuDCBH9HmPVcsIoOWaClEPwVZ2sjFUFAe
mCiaBAJ9tidWcytb416sCb/XlITq2oaVG637/i78RADvEPnQ70kVsxefXcj72AX0rLslRw1Ie6GN
bkCOp9RnNA22R6fjbWyjoMaQk+JZs22Uq2Fxqh2dENYZKvB6Sn26JxnmVjR1uXd0NZWuA0v507Aa
Gw+clBz7Jxp0mhvaMYA6mKWcAhysA9+nueJ7r5r4dVI6ICwMnYXqUH7hRGdl9CK+D7uL61R5En+m
hlviEzi1yVxJ0gQEkpxPMXGLSar+Z21RT+YNghXdz9V1w+3X3040jIsdy1a2169PeJm306be473n
mWh4sBxb5V/AbmgVYTpqiKAwAk2X7sUgUQ9bOlzErvExM/cfnsFAR4k7AVAqRzkJ0yxkVzXX+2mb
hFqih8q2Qe1PvFsnH0sOA8R6ARcYI8LJOG0ZQaNhBNLB/U89xBllqaOow0ToQ+L2d2u1xuqNjsQc
wX97axdNwLNvbLDA/JF9cIzoKiJ4V1cIcqlhQM4VCU/CGc/8QgeV6BNhd5Gz+vLp++UOOjchBRMd
JltHSCUv4jj5q1XBn2YB+Kz1/oWTRv08SGrZGa4J3jHoYAGZBRG5vXFGNvFRL6bSqcTBuio5WjOH
eVzLXATXGxVwrBt5gj3uZjUpScWVc3IaZefqd36bi5DdqoJeU7up8nrsN0iUNtGAgsr3GLSU8c2k
XrjgBVNL9FAlsoqnBsk5VJQ836+CQrpy+B8spORpp61vIBv3wEANLFWfMgK5Nf5alo8aCTEwgyWy
ZiYVyGGMgEqX7EuSL9NMpdGQVlmm+a8Gqlf9CPNB1TEwTf+A5S++KLABT5pBqx1RtzczxjSvCrTd
o+L817D2oY2i5U6RrNXOEPM2Gw2EWp8vWQffygqOMwoYw9tILEgdR4KQ0Wo455lQHzGimmxINsLE
/GkrN52fhi5ZamRpDq7zYzgTMily2IGbA35TCNNhjrNClJpiDMsUGc35JLoGbJz6nZ0ISVpW4d3H
5g/UJxIxXQT8GQa/nBed/npX0iTjGAJ0Mtv4pWdUox/ulptxXpIAnPu7oI3uGX63Ozk43EkcELEF
HS0Ehsl9uZLtS/HwrGho6lLgGSS+wvO5gGdvVIUSvIx2yCzmMse6+Z5Ksw49gN18NBcZ6rg5UMtN
6zECOWGw5EkakoQvy32Vf/+5OJ/NZLApHk+dUB0nO4JRDoVpPoTFWrk/tfU9+G7ShdDHQMZlvaKb
hFDO+3P/A7mMSYsQ4ECT/mMenOB5JzdTj/YlOPxJ59zOYki9IlBqT+Y9IC3b9fImft9k/RKZIMys
RihYvW+ckzN6BssYwOkazclw/n2kZ7G1wIjaUYExl5WI+/n7O708Df3u/LcjrUSHNkJ8O7UmzUcu
+kwbIYvHpYp4VEN1uXEgnEjtA9mf91sPkyFR5A5NenHKyseKDOUSZFCq7uMXLa4vVcD2ZMlxTUoL
bYJIv43ekldH0xpe//pR290Dw9GTqY+wjjnGwRh9EO1irUB8nLtF0Tz0pofExHZ58Hly8wlz8o7b
kG8D7Sxf483JN7ha8rfud8fCehS4o6mtJfm7AGwR9+a4hIoMaDfS+KCyXNj/05CKJIY7aCNBallR
SuzpThY/BnI1um1dmhHN978ZZFhsZXqmC78OWNCBaFFCh6qcaSdGEOsJzi3aMlsqvO1u7Q8x5efx
cegGSwZZU34xDnVCE/CisiN214li/vShlKCp+/cVjxAadGeQvGp9t3wj8NgfLn+bWQh7tEm5PHfO
+ycRVIhpxWx1T0JhCSf+0WWH5w9MaRBAOtsJFgC/aen1RqeGE7chDqmkdT00ZaZRYj2vfZLDGYB/
KydOfAEsbzMPlQSTbQlf7mkGGOS5fZZUq3+M+6W7jxhBK85czGfaDYZxAt/bLWkEzf2f98nlpYJw
WU/5tfrh/nzs8LP2OZRkGzgKxZEHC7XmlrWBn1Y6mQWlvgDgiVJnUYnb7TVO1/Iiv/G0zBZvpCz7
ieWGi3gmTUC08SBXAWODpnLnk2+eesPeHvM5CJ3UFMEEWpCsI5SMKrwYeyvGgyhNuaEPCylYzLrn
DJiMjBm7GC+yNKXYD0I+MFXX13MA/1DvNK/EMME6s+VZFLl9bYX5eCLbJ1wxZfb7GGTZhaerSeoa
v6I2Qoae57qrkrPoy+vquDSZ0zDB+YxMCaIyC1R7tErVvWA7E0kR43KQln8yK9crnV3TAgOcqa+a
OTsi/h3JgDfd+b2kZPGNePd5DRJ/FhYT601r6wTKYn3Hw8gv893orvwZSM7AFea+4CNrRVJv/Wnn
uA9wR1wxQKkNAX3FDcLpyJrhn5+oFAJWA0S6EUq1Reo6Enup+EcSGfcoTjc6BJqO0gyNlsssD5Lg
QKdctISBXSLemJsZlC3xxIRSXa9K28Ld+3AZKYKzdFrm1QANp8xKIjRZJpIMh0BaYTjmaVgJd8Ht
44bxjfzxhupM9MKSRMwouk8lFDzHMnRPio8yVqvT2hCpmWTyN+0KnxqYWCL+yZMDwuNReuBozRbm
9DySsr6Qfkz1h5Iyv5jeclJfDPdGcax8boOSaOA4p0lSpdgKa1tmQ5krz15rDggBkazqDiWBFFjM
nyrKax1Emr71JfSn0nqCkMY9VuESzoy6GcZkGQbYxmva610XTfIQUIuagAGr/RoDubx7B2jIsJ9a
TNmtVYGvID0Uo9ZMEpi88Q47+0Cj6+NsAMqMDfZwtqKHPG/IXgMz8ppRz3zl3Uk6i3wvdSFOyySq
5JIKEN+hflXvqe2YACjseeuVCClw9OBClKQYcix+ceiAmdbOs1d7hFA0oeF9DwZJnBC4HhmffWzU
afV9prc23yvMl1D82iUjqEj3Pyc2eqiOmD7sUAEVzTtFqNxs/vcjdoRdllpqFV3dUfs3sGPWKAE2
tQmUbyjJMxUkux1orLbRy+B5jhCWMVNZ3PbJAlVYCRZ84Jnl3cxDHR+uMVAyjoKueZn8jxB8Udbz
og+KeJ4nbp4c1heAzoUS0bAcu0YL5lgP6BiPTDIkLe1DS1W6LBRhCkjk524Tn5tPvWcWjvsKUn9l
pUn/5HRAV/jqcDDBXwEhWO+NtJA9c45CI5knV6Q+/bdSCyFlenP8Y/KtF+PpsaH4lU1pJhm5aFHt
c/po1QRpfmfGpWDDCm//2+c9JSDVeICKjScvKaFN0kv6l6NuhzEkdP3NSfBuC74IEG60QtwQJ4cr
o8YnWQtdPdQrCF1jPd2yF3EtYUcmv5u4O2Ff1AChdhWNBBOUDEJeW7G3sNEPIgi7HcOvrHrTII0Q
xOyeLDmFJK8n7GHjactevlo/wccjuuG5Ucke7mmahA0IQ73f5+6xVkOdMNTyqawtB/RmWJPyZko4
2TlbA9NsR/LLw7eXvJAY3D2NkWn87C/y3OmVsd9rJNsbHlh+17qvWpXthbnfNHA5MvFcuHY98pLg
9re1tTPTeuNQf8rD/kVd1FbeilDNqZi1dOMtXuwuzBS8m2s15cZggZukSVhQ2Mvd2IVBujLCZI4e
22GGN08O9xVVIRjtmwdjYIT7JEnDmFWTpG27C6kvw8fn5gXvX2L3qo52HJmgp30U3q55DUtDUwDo
Q1yJWKV0NpyyW0eAt9xk4qFHMnEQxL+x9NB6myb+Cr/9f86FCFY4MOiGonDn8ssLa/Rgh5yn8rOh
5CFpmTO0ThOw5D8MpizVvZZxZgo+1yeRV7P/h4cna/9MLuwGlgeae38E+Sm30ghMJQ/3ybhOFrJs
XPKzK2NUS1kzZ1hagxZtHE+jEpKiZWeedTX3zUpFYDr03Ax6S5GtuyU35FYDfTqmadAalsGYy/0x
ivNgLEy+SgqzztYPPfLjSRrkC1kVVr8nfHhlp3d8JXuFuVO6yDOl4SappufqDiAj+v3P/I/Znjbb
qdN2IAs2q1Vr9AfD58YkcLllXqa4bKopZxVN5pbiNWJd3/KGtFCfjhV+6XmSy1XdmHhwd4OsVZ4b
QjDxhRyMAtJCGT8E5+J61ymPEgB8h0NMPw5JgcFmuYhNm90lGqg54GDc5JMdU80jyy7/jtN4tTAk
5VpptaZRf5/BskpV6bWv2qu1nfX0b2ks5odql7mNq4Dc2nXOtDUh8GKA1ugyw0hE7wobT59+Q3Yn
pbnQ0JTUHfozsjfdwlEUUyS/kcy6E9iYv2W/HMoW8Vq+IbHMjwy5PDLxDH6/YyGsd3cRybou3p6B
Q+2xa/Ha6/48Z+3CDI3C9rNaNcfU/onXfL8O9nWDxe60XgdDAEC7w8lFwxBsIbRjAlguuYxIa3hK
79riE2FwSBNIMAPc75lwZ5WZFMzpy0PXA9e+99Cs7h//B8YcZW673QV+eFu46WrKkXmyjfYuoKcQ
rypWrP/1ZMh4xYCe5xpX845DKwDYQFaLhy+8ElmeP0ywBY4zrKPxPDkklycAaqs2tecN5YqR7/2T
3JjVIe4CuL+uQiD1JZ+QYuOMpzeW1YiBhN3i+ac4bBL+cbifqn5KylK5JEWKT3MorCUTm3x60BNX
3DhEI9I6336giQgGAnMhvvAn4OM4PZBcAELDv/u4wHoaBkQT4TYlVUc+KHjy1RM90laVFN/ZHrYN
yq9L05Uc4qovQMDAddDwyLT8yvuxRzBSJUtQGVFZvU6JqMXBTqsgnzK/vtBRuiUQzqiF427wJjFi
Y4ImDKDBC+Oz0saRiF2QIKa2w2XW/Ba6PCAPE5BbHZEwBKqxaSEJExNkwoi2yeXNV+42QVazssTb
Z2Dhxct+OJA1ekkJQHE57F2heVHoNbPXlOpgGRF0W51CBfXf3ai+0DCbLFiT3KJCldX7GM63JrdW
Sf33Q9Ya8/R9jvL2lBf81jemBBTFEjGwI2ATLOJ1rbxshKobFpv/v7D7QUOGsK1279uVhPs3j1u+
ttp4JASxitYarIvyWoG3zu26HYPq0CgK/48Dbv9yu/U61LLY7lb6X9NYzAMsdaqXNvtbrf6hOY4S
E/AoH6+B6+LCZvUD6GLG1C4gb5d4ydP7FQPrbtl+E4k2rANEQpVniKFseen15gubyO84q6776Smk
Gk6WU1Hmyn1QVF3S/gIxzjW8kZt1GLBWTYxB8BSPTRxbs8Vd8D7cB7flHqKHI8nL2mhA/t8s1w65
UhwfcsqXLnjSPVF1rgZpvKOgLErBspIb/mBqHx+h9x3FyricXyGWRRfYmPBvSJdj+kqTsBSpthjn
iY4NgLZYp90gPItfAr+/PB/SC5X+6GJiEugBIw1K58ex9rSVbHSqTu1I8v2siQSCsnWICh7Z1+Gd
TL6zgcWBsGIFT0hy2cs6SmuUf3UcOMiNtXLhuaLa6gVwMZqd0NurKKtPeh3p1jLpQHDViuTa4MSf
U7k63LhHZQnQKlATtCS5Va3pNetFqAF7aqjkbsuebg1VeeXN/0RBYnr5YfnnDgQt6vLqcn6mkOpS
z4CnG5c+Ooi0T6exwfLSS60teXgWfQf8kph1MYhYFCTOLZSDpRX/V1Pgl7QldbAukhVJPx6eyZm2
XDUmleMRZHLPvgCtYPtzjenWkaxgKjUIuBaQANHH4Y9ar5pVd2Zmv7rbh4z+EnLzCOImoJjlfgtc
xER8ymzDlBuFH2KRv26FZQHGqNN3jDIyJF9aX8Hl737FLV2AUVVhJwkQfGS5XMjtch559d96B3xP
IXhd9iFQm0anzPEgsNRC5JPeWDj3Cv407e1x/8Aqfex8yh+GaAycGBsD+KBWF5bMgmVaprCZIOLl
ETOR10ujxbuJ1sYLu34sGUbfE4YsbPEzsPBT39OOo0RWmNkCcj1SMmGkn2C6oPhYb2jTjIBHqE1n
Bc+IwwFG8K2vMjHYGyE4x2aW68BmZGwIDi79KtWNHkeqEY2HMZ+j/c57t/aIUPof15WT2gMcBwzw
4zVk3TmfoNOGdq6KgnVig6jMF5hpkl/QEbE3w8ZM/MBqGeiXecwix4vHcRLX5ZQmqMKxF7fSHmAt
9XaAka5Lrxjd2HuZudVKM9kU9+3n768AlYAv2NvL8wNv6ZG9WftjtCn+9vbt/OjsIYtz9sFFrTzu
uekhEejsAAzeGN/8zZaC911nji7u09+Gnse5qM2Y55ei/+TZ5v5IMyNR1BASxjXAxjeZTLmnnATg
XNIfFcEr5wSOrnuW1WsRIcptM1PiPqVe+BrIReiezQQJEpSh0Acqv+h34RpbJcIuUNmQmsj0osMM
3EzVwrvTwMl953DGc2NynXffX4JUJL9sBK5MabLNq3eBMZIFU5U9KsHKIpLu7R7IKdOnODxFkzcK
trkEk6kWAB206IEzs2O1sNedCIXJQ6IDvd0OA4H5obzsi4myhCAVMb1p85viJ6fgnKfTGL49nZSJ
w1lKId3z6w+Hrs2k2RAVc1UvXTuXWxDiteCPE5pQGVxyczoU+ghGs6YiHb9qqnCUiIW7tVessj4i
q6sa+B5a41a1epDJu3PTJ2zbWB4OVIlLXcFJa0lnKwOWiLBfTgSvxtjedk44DOucaIoaGyjbgfD3
DVGtpRQTT2IYclWVXUmeGL25gjl2DeLV8PybY0ndvpAl6A7I0ER+HLor20+8BnAUM0rdqAxi+94q
TyLsCqCEV3Yp4vPzT/DJVKPYP9f5PM4ylnOMoQZaH90dZgxSo5CAKh0uzPXbALGZJNWG9Nx3pm54
cmIkEhzE59WjxZnUb+ChTRy8GjsrjxHCRZLHQtClpJyu4cDNDeiT2vg43dyuyGitddM8GECErBbz
FLwKMND8NNQmE0nwosfmh1MLkQhqZOUbQvuZUHwYtflQw7jYBu6Q/VQ74IBgVVsQzsL55UHLWaz+
8YaThaD75u56aUHxVC5eXkxadEQoRqRQo3HLP1/iBe6UBTEpAuH23O3Wc0x6SukWkuUw8LzQ58+m
r1I6PapillsyJz0RKRqzS2OhLbeYrmyBLM/CoF5MWQqgfHW/bZKs9z55Xy8eAw5HU9XUB33LixQx
6iIgl10Fp0Sy6IWpaNc3xit7pZY9Xru6PC+zuQvyJ8Q0PKVlqwU4omdXHj/isXk9G1hJ0e+Uc2pw
4cl0Bvas1AmX6lnPxccCAinNOSJZDO94bIW8Uz2W4ty2pTke3h4auywMTZLcMcLufV6OnWoYZhPQ
3ZFw79UcSwMD5C9jn/ovKRBD3fl9I4HdJD4J0K1mYmKOsmwCJf4mzktPv7pDnaR1fUZYmDYnpAw3
BRu/1KHQWepJk0iCL/vuAr6nyu1T0ab3iN06l4QQ4TXd9zjReEsLNd6E04L85tLIuLPctzhEhoCI
Yz6eWvGj2nm4gx7BQ/uQPER+2PbcDT6+bqbrjc2kJsVZ6KEJ28TN+2/1ImBJ/FDKHqT1UvjhcdZN
CUq3pLw6omrHU7FoCTNEcTuEZrYTGLy/sCsZvFilfVpc45fvyVHjhQhzsnwJEbmV5fQ4javwOL2K
zpAIpAyriFKQ1vqKAQsdHaMzD0Lcp8hN0qG3IE5SwxQ3u+dDdOA3GrdCC0LLo1Gu+YCWdIfTTEGD
WpX1s/mJ9s5SI+TQFbwInt/C/gyJ2BS62fhkq5qIPwHMgYiJ3HgFBodZccqsuToYjODi5RyNaDiO
l16jKQx8WAKv4fP2lStaFKYhVex6gk6LFLFLW1FGV+bz2coAJh3ixilrxZCpnyFE7CLDXZXBemog
FNKnJKPxYCVvDvehF9Cmu/ga6kNlcQ15fC7Ao8DYiWgxUCVEtJ6ec60Ijml4j60QqeQAepJSu2/n
StOh24ZwD0BrPTpkOeXuWsb+hI8J28EVTl+PQw/IzKmAT+SOV3EbqyPS2p76f+RtroHCFZU4dpMh
relUoYx9tNAtSPHemgtJhYHeZ9pfaNNIBOAN1mo5DXPfSw/do7BUSwCn8zz0GOdsEMGMR1rEQq4e
+JOm3gPrqHlnzaAAKVQ9iK7mEnsDclTTw69R9eHjtgWTg5J2IhCyipb3Qhg4dJmOIoIjNTzDEV4T
U+/sD5MjYkMi/GLhZCaRABOnPnHJsQvDe3QIhcCbOdsozvptFhKylzWrD+Bb/oORpKn0FfWvpdsU
BeAGUr9iImODANFar4HMGi3bIqQZKi8cJNpc1TjiGMGAjM+RUvRyqVrlobK8xI6/piZr9/EAeKrc
XPv3HZrD08NbxYC1syY8xLuwxIQ+EYeiU2PC1ykSdeGr8QewgJKXwtEUBCjq0PEaSCrTAq9RiqMs
Dfld8bXbISFyR03ZGIH3A3pbbErAJ1cW0f0NewWd8mx726eoyeLrNapQMrsb0cb2rQdmi6SnWMoM
moXPZpRu3/kbDb6IiJ/8QXtUX0sJ4Dw5I1HkNDsHlSRob0Y46BwvPzhAu9EzFPA5aOTDOTK2/Zqo
zAHU+7BSqvwgFWmR5xqLMEKeUPWMgQeht82aheO7RmnNwkYghfPxDEMvS7uyyaw2OKejSpEj6vG6
eTucESSoCmBotZevuRZqjUA8+pvfaTS8yCbpwG2Z9V+8YYuC9szhbEzk3IkrbAz8LZDLjr+rAwK9
POMYLg8OEguetc6v2T1X3cQyku1jySLH0S4BXrMN/cIBaksAqpGldymY+mOXNg8SAY04g02xoSzG
5A6bIB4yufcdAhMowxzjdY4o8LMxpXjr16BcOS1aUujyh8cmNnH+coyASrOJA7EerjuQOZTCNAYP
sj52bM9KQR0vsCnHqMcy9q8cwN2/EEREpiQ85ha7azzIpoWMZI/woNaKOu+7BB05iuWQ7NDW4z8m
kyAcWgaksVCrmkhajrIWCCWHXZTIPiB+SzCRe7XjmBRV/AN/iW7QCKCCrpDKCGGFD5xKsukCJcYx
f+T2B76YnisfjaBF9zP+k9GnE4LZkzXxBmCjntyCofD1sA+qBjrAmmez8nY+WQlOarjXr2F8J1oe
F5qr1yINhJopQUL2iDFWnnok3sGbg87Hh+++u2UyOvYiiPRYKBKHDNa0IcFC0nlRZAq0+fvsWsmT
bKcSXIpEEBLPLoSyEitbSnik9ucdFgJwpEIlZOXToMDSmaXWWqkbsNXLaS3xfFEyCL4L1GEa4qX4
jQUSC2I/FnJFELoGSUNvf8pZ9wVplXBWFXVtSje1WWrgYI6WdGlZmpHeFoRBJYokguAFKagxD0A0
HVrNufBj2MHD0xwNfMHw4RJn0rCvM+X9+QnfFRASNvjIP7VO3hxAvpKH6KFBVaRkUMOavarooW7z
3mvutJWoT6U12F02Psz1mAjJpk2cO1Ctxl4XqzF2aVejNfBqJosR/e8ViAXYnatBgqMkKnH5AvCa
VyCu4But1rRRwAlMZx//e38X264rq6fEIyQt6VWVc0VeIGYKV5he9JTaDJQdaVGbl73uMANCpbRK
TPTXNMuRERSbRNYAIqrAh0T94CRagiJDN/t+dYwBD9t7k/8OhvEMrP6He+nZU4XS8yUdHuq733gQ
fyZiiGWUSkYRFo5QXqD7Acl/W8Jdl33V8NUTL2yOH9qxh9c2qcb9Z/ZPpJkLKcQIeT15adzwh06E
BPJOjEL/IwHuqsjlPe13dmkScWik/+qWkezT/gxCdwA67wir4AVvhexFXkG9OwO/nJhmz3/JVTHq
1flgUPGXU3YYf+RHBaqAes/u09l0/NURcTIEAfv7xtpZsBX05MDGryz9rCljPB6C/yWEkNsytgB5
EWW6h5aSp4DAXdI8qUW9XBX24sGRo8ACxiPWmyW84UNn6MVnXDy1vDBVY33HVyUHvay6VGCv/ipQ
v63k9FjX+nwAO/JRyahlGwK09kiArarO9XR3SZuCiL5RkWySvgiE5YCNRTwrG/YKKAnVfSoc6NYK
CWpH599V7VJIlQf89ey9d4Q6h3JhW3zpRytIGZ31UA4Wa90YgO9rUYQyMO5z3ebV4a3S52CcsggN
fKpVuB2Lwc7r3UGU+CEfaCCuGyCaPiSfrmgII0b/QlKBNZ1uIWpIU+9MYvjArSuoauP1UFNWUSsp
Cahv0+5EoV3QwCeH2hqeH7bW+w3BFFcikSEa/cH74d2jB5x11A0qVulYQngLcLjnMRfgseBFInNZ
etP3rci5KCUvPVnj79IOC07o9nbOsvfH8MGH3rUIElMX4s6YakGFNKYM62Wam/7mLWCGB/qpoXvB
llLNBq1j3vOVQ9v0WAcpDEzKJdhDk5uYtsUVT6vQrL/XDnnWwyJKqBwVqM7lxqI4kd/xi4XYRnap
YWUIkMycl1TvVot0z9qCgWDzP9Y4dZyAYdMfeQIvFuRhobJmhMz5g/JuqeRH/H5mqu+9AoioEgXd
5eSGGFppuIxWTeE2lQ+c0ZwF/iWz/rQuz6KOITJ5ym0t29WTxJPJCxoZWO+Y4fVmzTg42YMCsYEY
6GazBO+ivZUw502TRRocdyqgPaBfOd+6do2xZMJNyS5rBHj7uNSFk04ol1cP9OtW7LnUIV15+50W
MS3Q65CgE4eI9VXnBvk6bCTjxYPjuJHcyBgXIXkjKiWr+gN8zXDVWuMsTthP1i2OCR4LJqLFvOuv
fP+SWYvorXGryRmAdkesT1X8ovXxp3MkPuwPpVyuPJQu1b7otcWEViBqa5aTOxPdwwqysNLp6K7O
af1eV90PYW7jVbgRg6f0vDSELIPDLzefNsBNv6GHYwjL9gYGkQT5zsRuaTKxGQz6EVlbFcaZfHRw
rFpyFuVHWgLjk2GIGrx/l1qhG2+XJWi8VUoDavphIeT7A67ebLr4ELzYcC+l+ooI3pJXpyCVIdbB
7Pp04JP8oY/SkZiR4OC1nKEskQglgx5B3oTj3HrKEtOQ6BRLvsIkzoilmp/H6KWFFihdOd0/BPaU
s8jy3sFYKwfysvHr9lAxiPmo0kgbvXf9CQqGutPIBR9wK1JbDvh4PkVk1Q0CfpMMh3YGqPw0AYi7
sN7tJXqX6pMfyEBPhe4WsPsprvqFbDewnCSDOvLXMW1udwjvM+Yx3cpZZjVcuRvil/b4jg7frVlv
syKXMoMKGLG1Tf4Ixz40JgciGISmnG3DGQKXqOVHyaiRcouZWwewQer5lMlJe6ELbaawovcElNJv
GksPSDRyMhmi8Pd68OKKKvH+qEFP0q6dx4a+fBRIBM0AmMv+r6d9tG0DSgEWbynIv0KXA+7uXtLV
gPFtpk19dpyVlHooBHXosTqQ+xWRdOph+mG9JAbmhgJa7L/kgZNqTNhlJ4/JdI79NIBMVTK/PVZ7
aaylj+HN5SmA7bnJUk0raHBbS47YVtXuGBNV6EyfNvXuxVoHAhy91IH7hNts/G73J81dvhaj8Q6I
+mbjQLh4ND/iRj/gbuRXqqTuSm9Ss++gqBG2JZeQc3zTbFW7NV2WdRW5WOEMwWFwfdtvPOwhJrg3
nyMH1h7aCpOhFVHt0J0OwjRn+6S0yyy/8T4seIyBXW5zs5wxLJugwGukZi/DmPdcOHpNSDzeSDrZ
8FHVAUr8xPYcMt6ci1aAjpAxePnF551IDztTtkFMRSmssJfii4UWz991SMjQH6Ih637Jd5nkCoTV
4eg6gdcplcrb5RU+w1/Ht2a4M6MI+3aHhDforiTA2MAk3oAHaQoSccOzq5W8040QqmJ4WoXxmHjo
/CWguVrhi4PDTgS3fKOZmRz5LaR5PEuhJtZ5zGw/zGI1tafbCWUFFeVnjdFcs2GdfZ5YXGEMvHEb
OBdipWMZncaWs26UGMYdQIVV0Nxe7z/2+ybXbfIGyEo4hVYVCGiOAy+qo3PLmstuJitLfTNE/WDl
4bxmUSVslmwe4YtWl35bhDWFXqP9rpgWhLphpNDvZ8eIAwwL0sjRE/DJ7IPRcybhFAQzV8DkXlRK
2VxYdmTDcqwHSRpzwn1yVsvJ7FqMJIZ2hk+iSTyllYKUVYeZlYpiNQrscwYX4anqLzKJmoKxbm8z
g2RMsw4GUFX+2Nx8LyNxTstWbYxDEWpkemikPKVLh+UG266/5qH7kMYbRE7H65aajOHA0Qpm+4lu
pxMiukOQLWAIv07prqjNPLnlU78V/5JkA9/q/XeKIZEWc/8+xTJv02xYj/9/A7Jx4hBbCzngsUu5
A1EzUuDvcqkJ2AUiU2XRrRQ7mhS9L+XHB3pUiv0walfk6FI47UgdKeCxTIpNPVjxynidiYf7pve9
ZFH02bgG38vn7I2XfcZzu+qtG6NZSj6aJ1ytv1o3FR+nNHJ7SqAd+QWQf40ZnDpE39cAR0GehV5B
JW6xWNpdzhVcqYoYGO1ja2sB0MnjW2WnvUcgL+egYlqdWoUtKLx615zM65rZSVhd53Dy+UG9//tv
ZtMWCMdo6m/Qtea5fqTGT6LOX1KWlrzRQ2z0VVU8A1o/Xh04vB2rc7faazOcUmiQfpclY5Scm1TY
iPwUQQn8bbIe+JIpFhNT/Di7QCPzLriL/sew5qcj+NUuIEcjQPHl/cD9rPytbSecKz4YFkYeKG37
0LwMp5fQ7tSzQnv1sYzN0GVRId11NiET/ai5VOXw/Q/8wg96EiQDQrctNym+8hp4xoadH4va989k
i00d1nbiDPJfhOrYxIg8iRq9/R7yW6/VBCqpmlsqLTtBDvYv/AP8qt9mEoZEt/S3DxnEY+DrS0du
zELNVLbsa3PEgVeAEUQXVv5oUzbWNWxO0hHsyIj16qmENsxs1/qPbDvrKXOV5g5uA1GhVGFcgQ/V
5pxVujnE0ppmDsRoiepPrLZ7QmYLAy5bk3tTQXm+n28ImId9KG5DC7BJ+lRfl2pLxeU2Ak6ik38W
1byREVlG0TXybtfFyC9YkCXXLC+lNVqmaTuco4hAdsVhPoYrWIbseU2inx0OfpSUYfHQc6sDJ25B
YyAX5OcJ2yOhi8RrVIylfcWfV047SRWrlyqEblwnySDu7cRfRIv++/rT2O3oUEkBUO/4qY695qxq
5XY/owx5N0uuE03jv3xX96+P+ykQToJwUyQxADfJXwGFSjmwAR1pnY5jB2CZsrscg499UxHI8ysP
Biv0I9Q4aG/QvWaudsZo3rFERpIO0kyIjGLZqGa6dLzMPALllK6HIgdClAi4ayfcpJLdkuc7Yg33
t996BUspsRYtP4fwVz8I3Fl7jMslO0/II9OnvcPbkeSaOEtxmmqAsE4VNFeR/UYlY05gQ5WizRdH
0v0TQP2vjN2A+OTKkyKxp99cqMraG5FQMCjUfW5UsH9o643vKBDEp9w0t8hatKpeaQPGCB9mQwym
3b5CNPESknB+7ohvny3VnqTdE+emAK3wVdODRKEkF6KIlRIt31+nVW9ram4/puB0ouVuvlnIrKCr
nbRdnAwMe+AXbLVLygTuv3ruR0aCjLsaNjKUZ5Sn6u4BY6VF0kNS88AdGDF4qE3EdlhcbQRpm8an
4LjLIFRUfSCPVz7uxxLy/Uli6KowXLSzvW/WZR7erDiMDFcRTCANbTz6ZxzFIZ5oMxljSlqPK3IN
N6X6ySDyC5mCWe5naQgJDMr8u6/1wgsU2JV2D85z5wbdkcjZE/2EZ6nvJ/Crgn9dY2rx8/j954Ks
Ry70Dav7GenOXzNtxdYBxGACADkLzJxIPe0kcp19BCSB8RVD2/gAIVf1eOxHSAyFKogKoTkp4kTY
5nEiDsT/scOx9w95Byx33/ICMDlL7u+E6LnZkjMQ/CtIoEwB4nTBMZniJNDDRJ0tlGmS5j6/8v4N
KNiQY6XmYe3UjPB4sQR+kN0w8CM0VvfLW4sUEzTh3w3m0odrMw0LEnWkFvhJFnYOlNaI2btVkp0+
rILJ6PG3XqMRH6sN4rrG1nOI00PNrpHPXdUDR7wgU0KAovykvb/1coGfjKreVIvm+J3V6eAwODfa
oYaWjkzVh29Siv39AVy4ZZNr06wANrHwsOTY1I+FoSr2Pxd9sblWhegSWqa8T+XSHQFR3nkn67SD
5QU1pe9OUwZ7WbRnl78IEue9Da9OAoPmp4ekHmHj2pFo2BisaHiXqGol0vtQXB2FGZDE69p9Y5uK
g3CZNHLnum0kWtLDoBEwywIIuC0g2X8hA9mYAxVwmB5Ss8GvOzgva/z2gvMIpAYUVZbSjX5n4UYI
vYrF4lmQ3tvxo5lvMMOG1AXiCD2xxr+WGVrndJignbJzC+aHpyl0LDX9yrV11tMViWIigdqpysKs
dkRpIyy4nwXVc6AXt8+F9aI3o9kn9Re5PvWne3mngYxB0ZL7Tj/mx4sgtP/677MYSXAu4VP8tFGF
pIIwXXXr7L8y+rlyCH+zPlXASl3+O4ps/naaNcsxtV4sFlxEerMMzdyYc86KSG3671+UvOl9/oZ6
M9uR3yS5rNjhHFiHoHN3dTfY39j5cUEpUAGb0Tot/NOzpYafB296hEbtyTPDjFUWEbk21dcWmHaS
31ohbHJF4GGsjbGO0CH7VuklGXFABH19lkE3ENay3PWrbje53JjFW7ztMXo5kj2fIxnd/dSl7Ocp
E+XK6YKfeb+IMqvCZm19IQxtkLTChwmddeW3N+QenSe531nMf9kP2bUmCIhKTNtR4w7sums2XxlU
bIq3nofqZ7mZD1SEZETeF3F1ic0UCOvjSMUNw5x2VpG+XiLj1eISnwDx726WzV/67Rj0KLu+7XDS
msMSX545sV7rSo1oGpPuSANl3g2ZAKi9aEt1swTLXnAUSB+xBs6uAIUDrReCNCZb1e+YamWJSis9
Sdag2+mROfx1qJU0uZMxDQZx7gQypqeSzVaReOgZsLiUApN9JZU9rKY0wE0Fn65jr31uJ8URXwyq
2SL5DKHpUamnH2m3X7QYfJf3+NjuzFC6KIV0VqCQvv8n92RuXpOEFkbq1/lgvIq6wgj6LRf/KIN9
TushG0Ynr13jRf8EMEu4cbGu9T0yEE4vUzxzpODPickb1/OlhvBeR4Tl+GXv8xxrTy1hqu9J63n3
FSEZi5+jQTbMQzGJvJ536lEjsYpMgKSzZWCn4x6ER0q9D71BqLhO1BKe6WQ7+92YksAo/rVd7L2G
RCy+3fuXkfr0ylPB5oeBvBo6kZa9XjxZ1oVCDdAkc0sd7N+sNHWk5Fhvsq5L7PAF1rUuuh8+W0AE
gOfhrmokh8adq3C1+pyH0wh8fRjSNUqccan8qL8sLgC/pb65DIvWvfWaKrP+rAtNbcJQkL922zVU
WQcw9D5GZxqc1KTLWOKmjwqMTu59UB10lOOQ3PRLvylH6kEQD26/QzjgaKPEacYZ07SwP41bfvvA
oxrT823p/Lcko8Sb6YiQAdfZ1azSy2TmtqH5ER3uLnC+HMWeeNhssCKk7uCRBs6azAemVbOQrBIB
kRwJNMx1+xjJ8b/EmGyCklism39p8lKJ9MfAdtwSSGm7ISaYullOYghbxmQXhZuS2TDcZ/buoPbN
dAHow8ii71sRQk9RBL+3YnBxs6H+0BsH9yOyiPUI8nnzLmEi0tvQcPahVygFq3j77ed5rHiluduq
vYYrv8joXQMPQXmtOUl90/b38/Z0UYkGt82s/goUOs1uC5ZLdy5ix563yBBUlKJGjbNPaF2HjsOW
YxN5cSNmTuXfK7M53Vxu0nSGIYEGI8bN2L3SUBJUpwPsLM2MgIc01Whq32BOAGTYzjxHNgB93IOg
UT2OewPqArxfsWii6hKh/eYqf9FxoGY/tVxwawFc3DDj4g6Q4cWkz7WC8hhzZN2zaxtQJJqV09sX
Vcf6cLUDv3m29KU2juG3RSrVcMZcToxMQgZPLgB47R6jDBE7rqOXMfI6D/BLr8h8eUx2dZe+xBAz
HYBGV6MgC+EBKZw+RQ4/UMhIYWE8D8dswsR7efPLVjsr8+pmRiiiFN5d8GPHs7v5F3QK938vKMIF
9GQw7c68mPQRWIaPOIMjvv2zgiAnkbsnUCBEC5j/QdDIvx0NLjKyqnioCZckrKVra5JUYMSPkGlP
HcitLP0AvBTjh1OiDpBXqwGIh57WDAqwRuVjtf/n2RIHw41OkoviVCQnUtrIsHzEJ+kcGSUGD8s5
EjB7PL4Qa3913ZR5ys0XG62QJNQycSxuGMX2hsdaV5NAQ4z++XYy7cw61NsC3LlkdaNrPCRYVmua
XYwkUkEl0dwEXu3xBA+6IaGKF+bVkm/e+fyw81qcfRds8D0/gcvhmqGm6fHD3jel79QM8VntMV15
H7xBp9jQnNF4YyevW0LqZAlMj9lv002z/OtwujjlcFAGlvwVBCKaMzbsG7rfe1E8sgUDIJPqhMHn
0F8H07+gNOtf0Npw+zyoGy032ZhZG3f3boGKRNyVtPgm+P5gRYuxzEEhmxnwcQlJWFX8Rax+EDSt
fUFD5EPytqWcKyq+oRpeXZS8MNDLt6mY6l4/29RTPmIGvZcfrzYXHmrZ0B2cFndUusXx6ba3QORF
rmlTfZ+d0eqrlo9ufQLOUa4TVueKl7DFXsA88ElDK1ps3VyGmC4VOEvW+tOracLNibZecuARgdfy
M1U+kOKQ4ayON9FhqMwV0svJ7qDfWoV628j1II1QeG64GNH9Z1gDwYTvK+IhcgudOKP2JV4DAgPe
Wy3a6L2nvLbwnnywqPskjjmrfltu3PdDVWQUEO4mXssEX55lxSwqYRD3+EesTqmkadiWRlZe42O0
Ci4I23nhnC8JVHhhUC5fZ2/oIq8JNFAPrq7+2MrBNhsfXgaE2xZFzV08xqApexlJSmc8E2peaVtb
tmLq9o5zxgdUHs1DLfK7TiFge97FPw9SYzKFk/hMCC/aDJhZ6QVAecZv/8D059hN9ugwQIrI89rG
8OOLJArGuKLtEaR/khM0u7QQxZ/qvPR1U1LoTx2LVQZrdM+s81wgX5iTmCwiZ6nLz1NcTKbRpbc0
IHOWKnuGFVAyuF0LhAWy4HM8jCI5Z8vBzk19M3wqxdQJmBoMf9PoAinyYjV/3V5rhOe+BLxd/VDb
C5259wVyaTb218J7Hjd8I+8UlDeuSNTpS9k/P1Z/x2dEst/ARbvxBWx0gxUTLeLficgi8IvQ/n+n
5MiCH6jqJcTqjLYfTMb2/EocABxPCNlEl0Np38EvJhFg5oIRG8aXQ3HIUdAifXEykae+XJ3fm/lg
rYXn5pVO2kphPJ7Gk2qbU9Sf/5ygnjZNSZgzRY+7jiaKW9iWVCqU+nj8ylCG27ChZyT/9H4sDqbp
sDXzz3rYQE/2fxj5pv8Bkv81Sn4GfGhii9+ZqFTXS9qXwYqubV7tQIyR0k/Wfn1xc5CzKJgjzzs5
xF3Cx+oO/FFFVemUZrUxkkBPFpGnRIrGx0EpENPwbD8gLA77rQ4lNp+47GuwKCKLjicbiCWD0VKF
GnKJyPgbDXG0nd9a9IxhpkNsSpidprMcyr7Wqi4l753VGeBsPRBrMClE/BjWJY3f0iWVboj66Bbh
uK+EjdfFcj6Qsefxdmte5xi7CdEQUHPpg40nAue8sjLWXq7zBzuY/LG8EQzGHzzJaNgqhWFMWDXz
xRNsKgsItOhqdg1GTtf8j2qOk7z8cShAfszzVZwrZKasNXbNp76LsLZFHwmdQeo3efz3mwkztxJo
NPXZQ28M5wmRBW7TWvz62sTieyOJlSOkgg9Y56lWDTBt//9Dkq16VIdK9c9GZl8x9Wt+jmpbmDco
a80jbyBapfSBG+vz+uqlDo1FYntDGyvS7K/RRc90o9avSUjmLyOoYeyjLjBWnH/aPrOeio4pm1Kv
cFLlqSYuXtSW3OZFEoK17orLwV3DqHbnHCGTbx9l9ayB9iwsIyW71zYPTuAxqjhF8F3y3J9NsTsT
MsrhqMhWevuP61ZT8SYl5WcKqiPwZh1vCZMZtzWsFbF+ZglB7YyzY6Mht30nW635nihwW4MT2W3h
T8i21yFlt0VzSQqG7tiKqJO6y28Wb6p07qF/ly8H7rtEVq3NX78fIQBQVNkhDyLgBo+8T1O/9Rb/
8wAKvSsJSwZELSFH5S4a5OPLxCbmNCvLg+EcETXYC4+DhHil1JJ5hO7fmO5LU+hSkSNCvZdmXfyO
4QsA/vaxg57TOy7kQ5lebv/YQjAucxLDdSwxAjT3YEH7cBx8s4ZLKoUh4tRgUzBNES/lwc7qixvC
lLzrBhAcdm8R3AHnIQd2Lh+fN2g11dpP1dg6G053P/AtWV4n5/JsVwRoGTYTQTkSimvAyXhAjy6y
eZYjDQxI/JrdaIorFb5Gn71F5lH30GWDjGwFN2OqgMe6UMtFeAe08RsfF8UhYA77xkEF4IaxB2wR
rCF69b1+w1x5flwr8NoMnhwE1Vz3NNYrwcF2OUSuEM2JONRqXJ0BKYjZ7dtDSMKKfr5PahCKAz+S
ExhkJmZLovQWXDgqzklzqvCfsPrEBhcALtdL1dh3AYS5fkxAC/8+ejDZZfEvEUnu1vA0LyLAuBPN
VvRlWtPa7E5FTdsEjN37gGK5o/PZ09AFP+InN3PWUA/SAazUFCmhRzr7hubdUy/85fx2Ks66aTVV
8fL3Nbx+/+kKlFXnG0Z/YeSZeduMy+hCkEQVq9hivo4+X51XZSWXDDl+p/LnZsf+ScJfhSd5ONXZ
c19Ub38Ol5mvxnwo6e5d++zFbp9JIGiSGJ230iRwqd6kYSddHTaqi83z/gIs9M23I8PCYO37KNW3
6eVSqhAIIfF4/dsw36FeS9mTACAzRgCIOW7HgmiUyqFQPof9biJQvWfLGLSxT/BQVpPa4xbfO1kq
lZWwgOUKCVSEi4Z7F0I03nq0eMKznH4gP2NZ4PBJayMovQg3pp6uFaYwqG62ONhjchHq9xqTyA/Q
139yOA6dogcSNx6GbjCLKcNGeWo17bd23DlZ8nG/wwd8VNRXTNdGy9nKmfCWevelW8HRW8bNCGCc
oPquf1Qp1Oe7+jxoPkIUjxjYoIoIY9PRCAlPFA7WsMNUv2mhvU0cubGhCIlq2X1SYWT9A9MUCmcC
GvxBLcf+YMMFNUdy/M+RnzZ7u7ClBCO1a5OPdB5IRqdtq7QmPyTH65OgFZtIjywMwFYYKDBqfpz6
scumuXun64At92VlQV4IzvMmDM6tAIlPi2vF5bYadWzYxpFUwmWVU5Ar9oceeUjhQj2BfE4dPUix
a3V8H2ovtNZ1lD8j/6FnTHJ/Y2GugNO8kCY50DbzuPzmp5jASG87O7C+e6BAEVM0zuinY6U3PpH3
pbX76T9UuySa6tdAyjuA1hLIt7ggIxVoMMJn9+EP3f4BemlV+DwKjpa9oEN6MIESrvWXeAF1l5Fc
xJ3hm+ymoKUgmGEFCp6cOQ1sN4BbrizfPhVGp66qCu85Qyb5331LnFCkm9LVKihwGHqEQu0W4BVJ
D7k2x1uqix7aZkdWbEAkkjgS7gogt+9WzE/gRjNz0DvSTm0LVBZoaQvboiqRIr4hp1FeiyCzl5kn
lyNG/J5xDz79zoAQpxkUI46tpDsbHExmqhyz+/Nq1xmzH7lzKjty/FBKDEOgaDvz1Az6iwhGUrje
fkU6ZQ9NwBCBwIsNu5EGadt+5DeiojVy+XPfsyX+lufnCBhPr7kJkD9/wW5VtvNY/V/rllGNBdwv
MZNBZuacxW3wXQqHkvQ+Lo6RpX+xZDnJzuVYerYLaB0QuryeIsYKLHUshWn6pMJYTx63GiLM4oqA
gldHVEIa88fl3DV/4TER13BMlOo7Sge93jZ2hT5RmG9uUV43jOZD74fSviDxYvAR8RCojYZUTSbw
uZ2SIrjcN016D+iOqi3IqdPEe7+Xd3JimzKe4O/6HsifFri2wMZeONpu1E4Sc/kAAVRMGlQ+9Ssu
VvpiKUPm4K9C4y6dcj7QOc73EdqSzqhlALYjzVUvQV8hVSD/OFcXWPdtxDF0kJhDcAlzY6htGIPU
0PZazqHbAv79uNcAQy9eMYIoIRkZzUNJfTyhl69CnNreTc0zmWjWXzQyCAcOcupRGJNdmTmlXYa5
tydArSxUtPCTfx8OlfEIX+Fhh47Hp3Pyz0ZMwH9PEYs5c2c/Dapeeu47CDkK8zLrjHs0M77ild1x
EIz7EouoatfdhQeyVl9aLZyDL0SHqdamgEzEVfPJIEJnL02k3XAvq5zGeOcS0ge2iiA2L28qSmGC
/M1npkfXslUEKIzs1OnBZaYJppJx1tOjdV8OCrX0Pws7BGAWMjzKoU+O908tyxi3NwXEiaGTzIyh
9R9XZePJze1Rj9AIXZctiEKY6FfXHMc/y1GOwR6DUvHm48tNfNsBGDnIEVnb3LHi1HT6bLygVOtt
tAqt7aopMyVscuSRI4uj7jIZjsti5y7qT9hTmj0xAtiav02ElMS2gg7p6WQNu2xAcCO341sDCB9/
UkSPGZuMZg6cDOcvTBAgrEE2nXMURrmhcFEwIhR4MLDC3RWaPMvEaQUw/NM43Rz49mygfK1Hv8F7
KUSSgd5cZKwGDeTcEw5RCU8sV6Ttqpr6QdVrx7Il+EhgkuBa3Wyx/XY170264PFqBM0mRc/eP72v
0oV9vpTtcRzV6bGIcTt36Qh05z9kAnyMLIzWYGXUTG28Wk3W6+Ll2NH4FrJovRanyFqUns3iExkY
ryszlSMd8U7RHNd8mI1bIepPUtukphBHYw9bd1ifneR7V8uuhLYR2d01KM1Rg0QiUhxPPhze/lnp
T4Uh2b0O00XFX304RjB7IahfGeXEtvI1w1JbuISaEs1UXSZz//N/Db66TUm+CDc9Wg6WxibPuLAA
J//pE4Ep3iUDdHH4cSZvbWXkMLy+TqWGe2VMPHkwhjavSda+FE6p1q+B4VgXeJgYMg94L+i1UOwk
k5ESY53M2ZMdTwdXfa6b7AldtxquV8pvZ7k7I3Jinuf8jZX6YDf2TKJdaotiy+sHUNOyol8K+ekv
hhugTLLtOE3zs7SqdAVDJjl/wv0xLqJtx7VMeIimM+yAzGzewR/Np/1WcIT3WY7Ddw2wIaQq2fMs
DfMS3qeJrN4TBYfn1q/Mzs3G8lP7O/lwuqVFeagv42oSU/K4H55HPr5XNMxepPxFJG2q/2rOxW7m
BzV6OU1jBOFH6hR/HAKuEjqc1Jc8LY4yKBOquF9GZjYAxNnM6oUZZE6inRrNt2rCGlkVKHA85j7m
ie/6ozkaWhV31jtJ3Vd+hihaDdac6f62A3z8JKCkF0dW6tTI/a6oWlASH/jY/y15ZygGTRx67hn3
pbPO42KpYcYeBqUuDaa+M6kXN0D6K8kTuqvJmduZPhjWQkPtlwW5CqGLbR5N3/8CoTx/KV2CpCgM
M2UQHG5I8HbbhMblHxMUEJUPOsRlv5wFvxDI8wRKBF6jMbGXdVv3BweivlmL5oVnqrUQze3JRenF
f7nfAocB1Rzhoe8kEfHh236MYXNVjQ7XXy4V+jPgUiJGu7Gcs6rpVXXuTEFlVM+AWJoI+j++1NOS
ZnL++S+k9aGXkl5zbV9KpqvaynwQq+beDeEKGTGPWwqSJhUp5LDNuWnkSkCe3896XonbdUCn9fCb
63zRJvD58PVGf4fIf6OCHt6aaZtg1AVIkjtSRwb0jky/9gvBrXjaCLc5Lx0VXMVVJyT3ZAfCSnYz
Mq5qTUTyYOfNb3yfcpOE6tsMCvfmr9/1mTaJJVRp3UDMTpJObx6ReT3Qzo5/cTSkgTpkrIuWAxXJ
JlFv/ifIdEuUSbfbORPNU2BAoZn6aJWUmVxTYm8LwdNyU87ATquFzAH+tmpOYayiccdh2Aaqg/b5
3a2Z6HS5vsYcTGUAjcadchCyhUGxfGNVnlo0uVwNwb7nmmXLmu1ubnnknU3XdIMImvgDx6pjS5Ji
/apcQ+STFXWMmTOA5bas8oAVO20mnqj7CsJASrTeHsDhjWWLyzxTCMb9AOQvKtfPduUbRAbn1yon
J9cQSctpmB1wO3vSld1NaPFd+ixekFDRJQuKquzZvzZW3EIjzwPVPvpOn3de/+1ZjmZFj3BPVDw3
6napTlxbD2vrBx0LPWWHgWOUqiVuXxfhDSmrByrR0EXOuDdf7HwcW/xrBxox8wy0z2zEYfZWaPgK
bftdLrjIv0K5K/wPLL8Vvl6dJFsgpSIsE2TBZDmOFZU4Tfj4jm46oPWhWZW3wdfQanyETJZESZKW
qJZVaLbIlpV0izo2G70vETotmpBQprzG970dqekAwVadVv+vm+yRbisUyYWLjV7MDR0d+heQ8Dnq
VhJYN6Z7qPWqslTAe++fqGTqGDTxZb8qMzY4RU1g/S6BWys8tZVzYfjiIfsitlggh7GGSpojJT2X
aYTqrBnXwtS1AqIIw+VQYlVmLwNSj/LmipoTk64sPnRi0VFQYdyVMKGGgY4iBTd/Ij+MxzPi4vs+
lGmPr02mf0VWxF4VCzLWpoyDyU5Gko3y7Ck+MyO1Df/omVyuDwAHTkqEhnWXmPMf+8h0wO8G67P6
wdYwTFJWE+I68/9W1EH+j51YnnIQPTCRE7AFdBjPbn80uvl1xonk6K3aYKysjYHRPJh5y8PhZyyV
IYSDr2eVm6FBIK4nkK1NeHVABl9CPR4cTHAPyrTfmmX03WYfLNAJrMVCfjS6Tb8qYLyn7NCFOxJe
kMcNR+sQ0RtXhtSVpMz3QbQfst1oDeny7kSTruFfCYQUwBISYho4KbcwfEN0kAagGtEJljpS5f/F
MRfkcN7HvRqrIl1fYCcFyxhUg58EPYfiHD2JYdrTyWskTnadJJQ5SsNknZqyju7Jhu01/EzjAgO6
YTH23KfaTfYJRYssLy3XBsoI11RG7AWTnGDKScPpCOHKzp8DKjxNGahpEzut+6pXY+QFnHv7zMIb
C/teuE/UQavD0MZt7PgL8KnjSSH6kznuRoeA/MHX8lTCEP1QtWRnTOcC/jdL37IO1rXefS7JI1C6
ab8YFRon1/KAC+rh40YL0Tu6jcQcf6VreuHDVgP2S6Gt7c1pWj/E3X19i38Pl53wOZj+UllaB3Dn
hPr3prgXa/7l4sGwZXvVFuR99vEOZhvNgznaTn/q19raUSKD0YuK0Sx7KJGdW7Dx8bfIqvty+dMO
2CbRTFgKr3H8QzzOZdcJlknkkuDiBzBcy6LQ08f3NdPbC8K9ucG1ju4ULYos1eAPIbTYXw3Bh0bD
H1d3eotBQzxr04Ktkw87DZyIPlchK0IK5iYo0Dm95q+W9N29tptFitp/0FFSAq6rN/f9oS6Gifze
8Yxipia+XvDeToNM+msnWnxtNAMxlJKHHlbL8v9607TAswJ5FK+lvkwb5qdYv17R81iG7c9mcYgP
l1hJPE5bu7v+ChAtdlEPkZ86QAfH2et1+n5STSVgUfjBtt/EHA5ckctLxZEDM7PYzJAnWi0NDCas
4IYp4rwpXsvEirQjFMxQjRUm7jXALMCOqtSR8tpeDmwO4ZJ67r5QDolshulLueQgfc0YpoV79RY7
r60XfhEEYTnh7H69lUtMFxyvIYxsEt83/oQbSQlcTMJtcJCe+z8AFu0Y1rQHQsIO5YbV/IkEFHnP
jv2E7nJhacXhWFcSxCwyb0Wi0L5Zeb1uo7fbWM6PLnalDLzKMFaA+Puw+imui/x9+HpejVUhhXeA
J+cylHcjTrLEgWNcZ4HO/n8Ni+AesNIWxL8itdVB6zZGDvQ3lRwjFlPXSjSvODYRQjHwasaqgqkX
68o+nvRHcH27URr0x1PvQCzxC4TlOaUlLn02uWPIJXtc0YMxRfvisOyS05Z8bRGSYqqeL4fBRU/P
cChIPGzHtqzxULoqqgMXhQsUY3w2Mwr9ckBbT36iboYqEVsVGje+Xq7b6CgZ788sNgVawkdsGx84
+p9E+uoMo9yl6Aey4T8WVfiw5uf2/Oy4XurJLSpzsHUNeP4Ji9abq6PtBbXYBMCYt1ue4bIvB8nC
rD63snB/wQJIAemHBecsBvXRjmRYzyIkA65qGvkiJwk9ImZ8bycaE+FQ9djwFOjsICsTyJp3Fs+C
qXa52hoBcJ1XTNj9OehJBvRqDVbhLK26nFq7T9VHeS+QXhxtrCiIW8Gk7JO9JmgEo2ecUeCVW3ts
vfIN9UEcubiLDtN4lDzt/tClKAUEm8Z9vX5pMG3Sjwtpne2mAoIXmeKzQ+mv2mwRJcXoh3tpe5Nj
85puZVe6DfzlbbJREZcdEsg605OPLNlUWAAVzRK/Xl+ctxWaFG4ouQmRspepw/5aVNKVuZIV+6oB
4HnkHacSaeDigCD5S23nBJ5tv8pUMQ4C8OapJAAoVq17V+q/vsU87Jw7msVHYvOhys2Wjs7AyJb1
wSLE/3IcP62KlwGwo5fy49KaxksUAQVlx2wL3FM/I8z0EoeU8bybtNy54BqlyJWSScaep+hW3cf/
QzgzPFEDlP/fiLd/nriYTyU7IqVwu9NJ2P6JYEgRhs88pWgR+GsTghCSvFpv0SklidqJAc8QN1Ov
EM/zGD8ZKSCW3nph37J+kHhnkKpTjOVKo7qyed8YYRfNq8thVItgx9KZXdCzS1pD8+C+uKkb9Qev
UqNiIGWbfefHhZ2c8SJiu6hxB6VXINKnB+57c2mVXkpzFzMadIdJZBicDJcSoSfgimfpC6C7OJ+0
V2BZroIgk9Ofi3KJrJ+HJ5Cv9F1ZkVbT9JT5kH6DeS50HzRoeq1F6AAHcyfQmYxcD8tGeMFR2cxB
nIlpdB+vQrqftfBznRaWW3tfPMQdryWVyHKD9nYZrwQ82JF6l1IzmpL+aPu72c1JTgv6lxR3uhiv
G5K6dzCajwrl72eQcVNL55pts3ykV8PZJsZLdciA13Jhp9117Sti2XhMfAE9k66DfAv4i9W8pl3Y
NkTT5ZEEnFuVjQSC0tDBvF6r+y/FTx/iY8cP8t94EB9sDd3ICjcVuvqvZg38HmCPxAHT2wCv0qpB
sujFqPppIXy89sAQ7F6Ju7yAnbNrtam1AuP+8QFhHxLeeP4Eyl+Ul1HgukkBCXDkbj3eklRI1tdd
uLW7qY5Gcn2xypquYwsFTfYsN6xEy7AtlD01yoEw6dla/oKBDcBnUYipKBegJWyZ7facLULI1hJ+
7NdUWJ0XZaxReTqfmvKBNKtLoV7NndeJLJfynWsyxCoODetts1OZ32VRW7gqm7+hcxUN1er6qLP8
RAcG6AL3BLD7Hh1TqbnjphPFKTxlgiUT0hvyFUvp20wp1om/Z2lowGT6unVdegQ+PIc4kVOSPhHI
n4A7ZiHt8hi7ABDoXkL2QjkN2dhU6ZoeRx/Ars6An2Qosh9NDePgPmPos+626AIjbRD8IPnCoyKC
jV9OlHzTMJN7JRgRFfgCHssaEZyDcCS88iuMuRjpIRNLehxuvaMsJ3bqdS8mKnoGvPqdVMqMkT1S
pHI591EiZ5QdlncCfBelaDasQAHZOVcAczWxGc4Ya1TT23TYTP13bc3+gNDGtzmstTkuv9ozgXRr
RreS3ePupXexpp2DMrRp6nO9d9bCGGQMIM3JPHfMyYL8er+4yOC7EJZkwj1Ga3ErHSvjjCTi6lh8
hswftSX799q00uxFkZ/vcg3diE2FGihQSCvEsrYs2EUttXxl+EP/yO2pBWuRhgvht+bZfVSNkekp
H+XIgQUL43cYmJvU8KCR/jgjQrdVDKQoeDD6zBctD9iPll7cz1d/VhcnssfkzdcKvnKSydanWO7O
HAijncRrSzwjGPmYDkQ5EBdTXKFRG9ZljculkOxEus9V/E98mkiOwaVdxNbJCtK+Kul9JnvSa6vM
2Eb642K5YW/+UJVHr7NTnRMJdqnh8vqGR61EeKQHvDkIYaZ+zn0WBwY3zcveuh5aNKJL1deNO44X
yMSH19SgvNtm7eY41By/lK+l1EKmy4zfeQgoWAnZPFjzotpagZPGxATRU/ePThse2GWB3oi2g8jT
B2mi8to+69HhyGqEFY/3J3dzEK3fG4lWY2FdhryOTzZKuYW1GNs/0RGs0rGl8o082L3U7PV1ksyr
zNJK++CAkpcbmZZ+Wm0VsEk1XkYTSY5CEkYRx74yTjHeZvf43GS6ejb62oK3ZIMLaWtIQOBvcDFg
+O2HSBtWSvlxA8uj/ayXj7E/joTI6lZz/Yy1jKwVhJqjy7yoPACNMWh1WaESyRgHxNAZRVSE5irx
gwE6s5EP4m+vaXD7tHGs7biNS6Y6WWu8rR0hUKDoF0KkjWM6Cj8WMBO8xF5zhqp3vM3LK4In04No
VStJO6ztuG7y05wLR+SoItEGYAOxu42PsPkAQ38bdjbI+M+zG3nmDHN6ztI6PH2Ekv9PKH/1EXvv
zq+MEc4Sc27dl+kdZ71QYF3HkSBsRfy1cgEJtfN3if8i6LWD5gVjGik9Rd8Pz2ksEGVqcuiazh4x
QoF2GppjojNHwaDllQSM8xO8w8WWI8xdDXcQQfMzSuv4hVfCi/nmIPfT/QpWBx27yf1q1QI9CKlP
OfNpNYxkqn+dN5H4IwYDeuMkOhOwOwyaMJXdGhcUym+22eZlYNMYkcPHKiVD8IzCPLVpOR3dOYcH
m4fO7tcDaWMOuW0XTVcjZ5y4qL/qifGJHnGS0fkrbtHYfCkLAhr9RkzzIk01bMFT1rFguE/XYEnL
9Zs6QyPCMo0vHCL4s4JPop4x9Hd4gM8WkdOR2YcDm0X2ERZIXbC5cB/ucSCey1PVY/AwtImRXx4g
3QE7qHkwVGJKVcJajmLaq+MI8DCS0z/Av3S/EKzgta4eEqYgacNfu2kxJZNzm6Aakoh4kQYE0S6O
dMWLAX/IcPXE/1cyNNZq9rjkdI5NFOlrnq9rC72zHL/kManWlYvBkZO4VyMcB9K84carBrUOTUf1
eAEY9yNjiFTpFzvcgGE5p12pn79DrMc1CGtndwPzamPk0VJppNdyJ6VjyHUEDeUUgaWNWflgaNCU
KwrJUh0DENbxYCYm45qCNA2Egz0HONS7n0euNWWW4qxQ6uzNifx2BQ4GYJfe0m+6GJQIDVRIFUg/
bTgDluLS3saCUNbQ4XdStmOgsCotOEizRayzFepZonZi1E1dKQUiYCDf5jZ/tDqVna1o+3khBiSa
ShEosubQtqDq1oksnzR7v4oEpjNTTgiy2pglThZ/Efl+tdkjRYDJAL1Ay8kKXfGIwaNfqPXIQAih
euSOsizvSO1HDyyHZYQRUECDwMEOvJ9XnfCWW4PmWwAgawDQyrPGQEWSKgTPVbbKpFQm1falJDPJ
iWAg5eHjx7N1aHl+FQIGQVPZcqGMGLsCEVqPujOzoaJFehRj9/CDoe7xsISrrhIcpBFoN3HOhijY
5Y8mDdpUd3cs/i4W/oQA71mNvQ2mW1EQs7m8gdj2vLqPZliO+pI2RvSS0EC6OoX4sjAuz14VdwkV
GNF7UNv5gtBdrQdWWpWhboEdTGvGGhndhzDg6yLD3ebwWo3HJrVhqcQFQ2wwJRaYrrBtrd9OGRnW
bSkcl783oOwnjYwv0IZNIJf5DVOr+a1Tt1TGdJpZpDH8mvNNVhZLTylU/I9+8bE4fw6I9f/5o4zB
L295zV+2w0oJcAsxfT/Uh/waMm8z2fX+/OkGs9BCwIS/x85fZD9S/ZudcDLTpbdmoCxPIIU6mOYT
LaXyS4qEgWL4qR8vYHs3d5cWM8JquFVKAvywJ/ci5bBIow4khD1oR9K7nZzNpCm3K1vpcGPKquZF
71CZMQmoSB5C6pwXdVzUq37n+JG3m6c6JDxDX+fq1I58pzJn3SD3syK1uTYX/fIG0B16PONxgqOH
cMAFUDLK5wt6Vj4rncb6pI7BvZbawJvcLZtdT6+dqIlIMVHOAnhs+GmlPhrixWV37HN7Y+qBjqyO
iJH1hOErEOR3VBdr2Uh/2ggTv8i9hEcTqs+G09bDGv9rUUjYm9KwpWRCaTVJCOuT6Tbv1xooMwa2
pSnuMCQFsZ9SKxgKMQ9zmJtpWN6nU3eIU0PMLLyXJn/yblOhoq6BbqsPgPUblYH00EJL4FTy6jB+
+qD9lr0SV9y4fPQ8oylgLjOF61RBpPNmzq583CcFlk7yCbFWxG2i+1Wc3BGIX2SsLF2pXgJG24pP
oJkvgT5QHkK0WsI9v8k7yRA/qZp8Yd1/nP6fG2Acz4dCjDm1w3efAyselvtW8ZV99sQ5Vd4dC+Oh
9zvdGcbS38YnvXernAgKzGwQJQx1yUA/nkysBfN+EkPYUX0phwWNlqrL6qTM5n2ATkEVrqCB5CWh
6J7ka+T1NIjGXjBqFaqhuCOwcbpYtYoMTO08foiESAMok8sJUU8sVJZAaSt2ThN3qyMfCEwvpnZQ
wVh0eVLtGe7VLV7HnmnKpZP5f8BNlFdf50syANoVP2n31j9gfoKiN8//xZFcw9SkxtDDxniJdVBD
N7U33Jazpz2tv/+Kcp1RVQ/YGCs85aqHIyrfhNwrQSpo3JjILEtXiTns7b70VAobQYiVNRebN6X/
g4p7ML41YyOeXStCHvTo8N/BptfLxwJJUz2dALYrS6pSyJCZbYYhrgSA2dOcWVzjyf3x11erCg7C
n0nF+XDVXAi7MaCXecGMU7/75DBKyg+Oj8FclfHcB6XJLPz/meLeHy6XZPVEG+B7DilG0+zUChvg
d3a3uuNW14ruAN+mUNHb10VxCzVZaA79CaVM9ZBLgSPMUiene26RdE7aUGEYD+g0mqaTcLvr/72J
W9YKh0rcnLtk1uyLc131VO0cSwtNtz8ONh4gT8cUcGHF9nSJtt4f6Fe1l8f3XVkwIM2WhjhxuzLO
Misy13pmVEDZlu3r7pVBAFxgyL+0zFFjlVECYcB0nkr+rxzv45vDsXKQgfaAAepEMseiHovHEy7C
MItIVftOPsn2ENeRXGOqZLoFMdFhyajf7zIAOIR1sct5xn/Ue26bFmXvxJ181M2BQrFgzxKWHbE5
d40tM6FvbwU7I/ld6R1xzEroVhFnkl+rQQOfkcaPAlJMc/Af6wEiv+OvVOnYK1bJfkuRMtezwpqM
hYYOqdbNJCuII7RruvBw0KRoMoEMA3HY3WIcDTTxifVCpn3vooN7fxI+TT1bj5mHlArMbEVpQ19J
FlHHObKx31KP7eJkN/lcrSBF6JbWKEDz/Xn+1sYLDiZz3Z4ZrP6pvziq+CaiItyI+hALkDLpAMft
y/RjIJj0WHiLt50DsAKGs324hnm3oFXD0kvoBEB4QiLoLP0K889wrUhYM9tBQTDWuGDUF5e099LO
Wck6Bdn2p4w58kphoGTr94sbwqkzBkT1qb2GyLS/a+6ZI5JCdEaECPKfBFK/yxqS6ETIQ7f6Zdn2
PJzLca8EBGCJfKvzkvbfT09i5EaDiSOS1u1Cz5arY+GMZCMWauvnCfH9NIUpLoBdtKQfdq9ASJUE
9T1A1HVfqWrVTRWOybcfVfTKbd51OIo+5NSbvB0Ys0s5iVnbzqIgPCiWHWRGv8OW5dcKSwSWJ6Tr
cFDJWcFb1rpMj3F3uswqVU2lkXbIWA89On9AD9sJp32JLqn4i3jRtyCQUEp7o5BtlidJc1GZ5p8T
jJk9ncFgj4n3FhTsdbccM+le4FK1c7GEng/e4XwT2N41OHp6FA7PQ1Do0RwoNczBDXlIcIf6kn9C
vF7AmOCHQ6/+AufT+y5OZok5cibXDqsK1J1juQffmDhv3ylc/vNZyt4dVhZpQyo0Bj3b3g/HhXkg
MaOsfi6+CRtxseeRrzJfh9fq4+6qnCEO3UtTGtZt3t2zjOLktAKCywZyKlv/l8G3fJAt8DHVwXCB
MOU59CBIW8GTwiBzBcbfMJSq+qFMUvnKMam9iFTdjmal6ckdPBkpWlBWeTJ0dbcP3VpLOJNor7Xd
FUx5wQR83+EMXP/NEqznqXKqWqBG2K1bT7VhWAm8X0Yey1coWzIXVoJw4jqYd/Oqm1x3BBWFKUP6
PlvAC7PQoTZ94L+RouGutnvpnVjP2JQQJeZ8NHDYEeA0JONLrr0HB9W2izkgZ5O+uGvpDH3ipKdu
lf3GF2Gkb1WlxyPu8VKPAXGoVj58ExyosoemJuPpH0CKlw1QYveZqlQajO5hWtWLZZqDWNlckHSs
9rrZGCV0Oy9SXmiKEz2QGxBG5jHqPbBi5wiPwLpMnsJj5tEQhVMjlnr84VBSumEFdIKYvf1m/haG
miykFF+cyiZBSnm9mihd5mpGXgWpueYBibxV9ZGpOzCQrgUgD0VC/MtVc3f+nhAPczoasuRxgiVR
P5vhQn1vBcY6nlDiZZ2qJBfK7B76rVgRr0hCVkfU0Xhef9QUOCu+DI5wP3XLkV9cVahm8NO10N/F
VPQFZxjFXHbwjtybRGD5SU8b9JMv/VhoUYqakaTHHJNdmq0LU+naCn+xudN4TqUL1WIw9VEE3dwS
olEy1DYRR4n9pCdUmUJlS/w9BPbqjs15aCunV7pTPppTVW7Ux6oEsexsbewgNF7GQ0UC5JdFAh+1
BTLXjjdEhw9Byp5Rz5fS8gQMipm3Xf4QLA+x9z4GiF+7w811g113b3V39gOVd4X64a99V/LOdko9
fIpe6188MfztPaaQenecta73BjynRm6EhnH9fFbfkvwP8D1RY2J3BKpS4eCg/zp5rxkX/Z/mU4eH
lVmeLN4InMB5Z/4lGWUfB2/w3yssKQmOjC64GMi4g7uavVMGHonFqU8hsg6dVeT3x1uNrlhyyhoL
oievrTgaa/M3xqQMeVI/pEFsE1752kolFTOqDdYiChnO9wPPmMoIpQcGLdHeB5XqTt6aCNnqI976
+p95dseo0SyIMAWzQqIiN7GaF40nIb27zJ4vKLYGZnQG2JLmOQN/IgQJcP8kWJaQNqfgtLuyjC/2
IK0LLLhN6ItkOJywIdAr2geVmDwqXlHlHqwhGacnKXNwQ66JD1Nr6LI/XjbbPXSR0KaQXpxoOV3p
y2W9IQ9LieVEkhu5vePjXYMAy3lRQQ4zQS4skr5E+olWB6JWVMuTAd9TzQmuks4Q5Ajf5JCIa312
wENeT/hcIDQmXPJFqE/pBzBFYp9grw/+gJa442ywhUzapJpWFpH0iahkeIrt99zHMq5YANMSMpuA
xhd/ImgV+dFt8g7bJ4FCPFpm127Sl3iSic74jAN4z6i3QF3qn22+gfukl3erPuLnL45qyCHyL9EI
oA0yc6q5qzDglv7I6IfNiqLek0lZkXu/QwAJWu+a3wFNO68t9F3CHB2KU7Z2TA+kgg4p2/lewPcp
Bv+fibTVj3y4I8sG9gaTsDhp0kIoD/u52lm+fZFbSlb+ctaIyMSLeeZ8Om2my5Zp2AIyDGejRm8G
f7vvUNBAKrEBUDtBE0/xcAl1N3IuegoeexB/4fgeW2COs/BtkhdT0l/n2s9yXnQs+taOOYlNS0Zo
J0Ek5q1Prtazefq8+oOufjLjH4PXvHj7rZ7iv0yzNx6PYZtNX6aVDnY4UR7qihF44iTs88GbMH5g
sV5eUwGBaQszZJ2s4+ugtMvqjLF5UxYtrXm4GiC7fMW+AQZT9VLA7IBKl+VZakbGsmwQsI5fchnP
VAWbMep2QmJWiobRZgUIgHy0Nfz+R3gEGMtDEl8xyo1wMPGo3/oks3mPwF9ce9eioRvIlj1TVJ4d
ZWj5Xi4vTYjqA035BJLiWRYvevmGkV65eNY1EaHkaNecrmNCeEk4REMydN6Rr8YN/8ykkdF+QHbA
9lm42emmUd9pIhDjHW2UcVvvL1hPG55hmt44g4yrvQZYLiLBToJJmjPOiDSKav/DCNS4FEoyUuUY
wcRMJp80oBDoOsBqD6BkCa1rbdO/gUk0hF/oEKRKkUUsmCuRqbBVD+/IsBI9eMQ2repMq9YJ20Lt
2GXeojuHdweBNtF08hQ5QFk/02rmslJ5l+AsGoWYJdhKP6k3L4DTbHwTPFcL25Rwgd7qPxnxOntY
scGFHtjUNZY9nRmGLPVgoWXloiwyw6le4aY+WajNyS5ZawM62DRQsHwr8tc3RR90OlHjjrpQoaM+
4MJiuvbAGgjNiRmYB5h26ixvTq+7VfImfFgJ04MFur+u34gUav47s1rhGAewOv6OdLGzOsYct+3w
2bptgcWhMQ53rg8tpas19zGtP5UrfG1iolE+BZDqe6BGVO55B24/iNMyiIFFpPSNFu0GX9H5xLue
HoKdzUgVfkqSGaSbJSVbKqT6TAzomNlfDNCQlUS3+zqHzeLHfY67NxOIbTr6WiQDHJyOi/wNPcja
ysdJLfajSSSnJAsYFRzmnwzIy2omcPVVCWzEXLreKONn+/dsr+KgzZh00iQwpYdaKkIr0coBI6bA
7fuP4AqNGQaTbsFp92BhXfcEZx1TCJZnRZFTbpuHEULn9PbzDFGj2DJs734JfqVSdFJhbzRIXD/t
+urBSxpSFzcRn0EoFAhSXWzad0PnbXOclY1FPqddY4+8aGCtAhxX3a/BycgpFtMjFmIcGvziN7y/
nkkEJHrjXx8iTBVkC4CxTCnHctEkAPOROsEdAbVUSUvbScDdp2OUpKILJ0uAXeo+yQUQforsn1Ii
vRZUo/K6QmlzFWEHDb8H6CNLz1yQUR/sqtcjd+wyLvPHBKg7E1sMwIeaUcVtNtMH+mI2T4ToDt6b
5RI/DPuRiI72RS5C8zyukq8y49UxYa14katX0AW30kGVkSTPpkTXoXNYxI5MiX8NbUjvmyTwTNZF
zOSI8nQJPQgNDxjmuVPaTNVsVI/AYD9uG9KFopildxfCx7GjZpuoDACrw05QxL2QUU+A13h1io9j
Bu8G2n8SLFsVkZocg9ZaizSi1Iu4J6iVHkkeq5z0hpHDRtf09HOJSWD7tMzRsu1X2UNbYwynma0s
zUkF9Kg8YP9Zz8pATJxas0t7R+oauPhvS3g9B5LR3usdbLRKO962yJXAmRT5mHW/KIdPthDcP+1C
o5qPyv3l/lDB2tuYqWWoOcUoLBmwF+zBfbIaOy7CaFi+XDx4nb7ln0epPLCKGDYAiDIfNscenPBr
O56+7owlSoKnjpsjZOZzcnc/ePhWs5t+Y4AUGZ00U4DdhED8HCdb10TOgnhlrYNPYX51e0tlgSiC
Fx50gUpZ5whW+iy3GXputXhXlrnhwmKGSEFcYhsZySpgXE3we2Lvh+x4tH+KT8sEiG5e1XhOQXoY
wenQjGh/2c2zr2Zg/O2sRFq0yDDlW0VJek5+DphMhBZRiU/s+TFsCOeuX7SPg10d18xPj/m6nL2G
ja39rO1DQPFKc2kVoR7PjXNEq9E3Hz7OWchRKkKRTdzZS2+zLhKCItOrf/JSh1BtS5repSgVlHcq
qOsTkRfIY29hn2ciu+JqyM0QOhRXdN9FnGoiKHDcuyFggxNTWHIMAapuo0gsQx25m9OtEkfu2nec
m++d1WGVX8GZkR6eiCVa/Y1JM13+cQJDddS2VtsrptqIuicQVlwX0Lcz4BH1dP739PttjMqr6R3Q
utvlYSf8mVhCIVFOHn4Bw6ijtcGcjkgQhAmwRJLlgzOF30ExB5wg5a6D5oQgyQLHEEiwiY7Ky+sV
bK8ow7OwJqtJvIw9QiFJdjI1+iNAWys22t5OmeTtjrPdwFTWEWrVfH3YcsU1XGBc1JzllpX7rhkL
lFy5DVGZWS83wlAEz3gmo5PEsf0sXMio9bCr9vUbSoChVaw4L5WjwcDkDwuyIZGeZi8MASEk4f1H
GLM+VziydLtzAX4kIcnwHrw3QEPNou1IV/Bp0tZBD7KtKRlzlIVndbZeYx0goOi1l3lwGh+B/zNa
+DddcOgmT0Abm0xVQpCxFmjinAKF2hecQVH6WqwLUIn5j+q1nAH6r2WW8fi9EDcDc8OCL5izqaoj
mD8uheqwbMlsieEBHjM04nXspkVWLwt8HMtCM0/TAIZoV7bgXm2cSox+S2fKJW2bAlJSwDlsUMsh
mp3Gtbx9aR8lkflRnDNqhIBmcno5RMlABZdO3+Ptc0zau3N1uSMydJex0h/g7Fe/nVl0KTfhJnY4
RD+nAKnxwIqIrHu3mVra/5JHx5munKNFC0nm0mql3mDszx/GANi3H6Nm3MStPZVFtl9ngbYcN8Pi
KcdZD//k5/CdkQ3Ie1Ong9z39dtISR2QxQwh3eFyxExnlEKovh44FnovqmIAhbaUdecvMQFXjmjg
vOgPnr/zX0h2cwpp47DBrLOhunLYW4uCsFFIOSCW0tnvX+C94Xn9dd5z5Di/WLsF0tAmcDo2uiKi
EZLFUIVanQEdyoABN8cd7Ru6Ibh9CMbcgNwCBvJTt5HhvZDMcJCelUdPy8ZySp4tAUI+tKHs7UIE
5NZPHKxj8W+cACTDOiJlD/ayy6nj/hiuFt8x8yS9Rg/H8AMZVoE4MEuXDgE+POq45GTFdtX5c/Rr
0x8cJrrHdYMitnZma1SOEbpaBunL+rnqgHJ7N3Z6/6rceQEuU0/b4YUpz92oyhWTdVr/i07JrbDd
j6XBaG2+LkvZTQ3JnRYXiOx94Ftqo+CVsiuBt8Fidrb9Cf0lbKSNYyVoeQOzBsCqkINvO4BFWkr9
xP839ITDWtAPc4t2u+RK6NlQBREYpLBN70udp+Ww+T2RsPUpP+H0bRKoQwHfZ1vSQ9ApVxbjC5/a
pkTn2jbIHZb7j9Dmljtys5JmuGGvqcuSllChlhwocvxgwiwgPDSfX0XHEcC9pGBrfOi8efoqCO5z
1raYAC/xcVN6ifMzDSEY1YecRzRhoGx9GhYPZKNqMe151D8Z4mrhcwQwFCrIvwBq+ak77TO1cP/M
zAhIYtZWNtbMMDRowFTh2vjvmX9uzqId/7OSw8zoBrqVNlqjSV+jsj/hiTQX84AB4BoAHAUIGjh5
ZC9ditR1MPJ7OB3ys7u1NxV+UroLw58qIEEmBvNwFEYyY8xd+uhGaddJuRjS0hiBwprg0BjpmaqH
Lcd7OVISno1POuZSGF6wS7P19h8iGseknx1IQdvaFlWCfLVffq+5Jf8D3VVv7T4YKCHg8pvu4HSi
ipezalMyZyiTqybWQpHxjlR28V/0Hri3wWWoHL6EH83GOqygZ01pPpgFFqvz6AKAReG01lt2JDo3
i1nvFJkerpsZA5hbRNVpRJ5/oCyuj+GCz7YwEMzBqH66Cjg/Ib/Td+WiGojpBr5UlZKyFeTL0FVG
jqlHa1kATOvQtV7tV9Mrc1KyP1ZXLyERzsxfkmIPTl9Tf9n4EGQUTyvs/O60xns5FuV1ogmuv4yK
goTQh1z/iyk03Lt90iW5YvfzCm21GXEpCglBljyDbP/jyxUwvPTFG2mAndxtb1itarjTaLl8jNcp
tpA/W/DKIXGGDC1sBeaKsi9xr/WW77xLLKGnLJPruGk9p9iMyZUS5clBR2sRNcEvNWkoVzlFmdwc
DJTaRFRCmCY5ktRj00G40Hf5GxsYMR+OQwZ0WHTwllNr6adBj8wjakWV8IeiK13N8GDXgKfSU3Sz
1+dn31DocWSjZ6Da0nZrEr/C6fYx7E/E9aV3r3QT1nTBWsg+Hing3UYl2X4xxq79hnF931nKOzKY
TcS8NFyb0aUNJPO5Y3Lpm2Ry7cHa1ockMzoRGEVZb0h93R7BQyjokuhnEH465Y+MyaNylXO0SsFb
0pK3hkYJv6nFFt2c8++I0HkEMCCAg8LiV4jxIi72GvHtWlMYm2MslntdF3iK6ZgFVJgRzZQGTRQW
aXZz5JnYyFfOHxwa2TJ+WkDAviHNrWdFudLO02GMAwFf11Ptzb/fxgR6ZahnnaVx86WFm804vmPO
dt4rdOzg9ZoBXkYFUbeLWviS0xbBV89/+mbtQSfyB55el1wiSejmKiGrb2KiG+k5YoK9Y8BHn8N8
SNiyWwZIG9MQJGVZi0jIraZcikJb5bk/ZLPPlq1X3vkALNsmkjD/44NrtHze/87pkM70e77gi1kJ
Sb7dmLBx8Va2Ri+Jx+L+DATAuFJ5uI9FkWZTeU5IfDwp93z4lidSSlbHlzo2jFQ9QBtodD9VhU4d
o3J97k6OTpMSBzKOzORRXT5eP1dHiYxtELmR/pQ4UZtSJVNAR5PN4UkyEsciKRlDFH+eTqojsrNQ
KcJ18rx8MdPIhvj4ic3dh/9/W/AaIoeRnLWqY+nhVvETLhKXSP2YJCH94OddkQsjN+7qgh7cS9q2
untW+OEG+z8CgnDwcg7R2HBXO8vExlsXX7Z2ukOjrFAbj19ZBumSqqgMrF6r9Z49Bw0bjCjXoLuU
5G6YCFreIm9lQPeR/1WySnPmabi9RTRyC6ep22LLhweCd5oOhauiaHOhnK5wBE1lbA9HN8XD5I3c
l3u0/7Z5G6XKdlKj+oKmbbmu3VCnEqjdgOTKv0K/cpq1iTU/55ok364yW5VXj1TLqlGGF1j5HYid
+4ZMOeTPxhUwT/xbrvOKmpzGfM05YNexO/cj5u7raSfuRc+uQhCY/hTGIsWrwq3kSnzhoTmUHN5N
5IyNCMpUtYkA/HsokxFLiyQj3XIqEpsVDN1HArMFiaKAgAGMLg+pNxG3luTzOC+VGt1wjFAO2pJS
yliSyJhduorFd5mgVYN8yc58uooKWbX1BJEAH1aAkDpkp9BfWreX9hyoVjmsZFLBwMqlrsJgUkRX
8cpiSm/LdW+3f4MatubQwKFzm87kc4upr/PHme5A3q8mbGc+exxHZ5uzqGsL4U772NIg/jte3kOt
9cusp5wl9Wze6MFGjWGQDkJv5TC/Kg/KjcQNXNGscmw1R/H4+7WhLiP9RC8UzVMhD7glBTJRIGWA
uHIM8XSECN9uEcFcZV6DfjyQ5Y29vI9Bkb4cP4k/WlseADmJZGag0gr5x9x5Ci6c1ko2I3UuPALQ
dso9+faQnfYRd1nuVHNNGTO+i9wTMekrlf/psrPYTP/BsjB5q7zpqtUR7h4/WcZ1bG19VzqGbkQU
RBQ3UscKxi9bel8a76c97tS4SxnYE/OOA1Cdi5QcKA4jTcqwwD74tFm9ypTOytZlkqV/Ty1PieQ6
SXDjo0m5htLVeG7dcIcDSUNSD+jcBp7V8FW12L8GfsuKlTc/WW46GODqj3FXQvKlrXPlhbtzRj1Z
ScXjYE9DOXpmo3nlHRfPfBw5hkpme9kmfT3UmdTo+pYJOp1Ewc2cvexn8ivRveuQ3Xq+beHDP0Jk
giI/HU0Ucgd934/0IJc1nPR5Y9aUL/oxWe0MNRDMbrrZScde7x3cuyJVnW+yEtb6IoYBK+gZpUus
a9LEaZgpW80iNznjHntSDD8LPqd3NJepf+aO0FiMJ88e+eY5T+y/likuN/4YKPHo2EstqZAADZHI
+X7N9IyaQ1hj54HOP5sNMlNb9I5fzm3lH3sYRpxGqTOZK/t65/kH5PPXU+JVWtHU/2ooD2U3XicD
uoYGp1FuBC78dC5V2+OXKY1hYbAawVyknCP70L1LjxTvjCGO2zVK75zKrslPF1UjuP32zWlKJI3H
sjPmR2I9kFDysYlwss31De3m6ioDSm5sKDqN1wXAkKfW9SW6GKsB26Dg3O6zXCGNeP2QYxeRNpwl
yM7BYZKGeQy7wLwVWWIufnXC/R7hgFykisffSbsF12aMUlycNbDO2V7wdszRN5M7aiyOvofMsWH0
NojjPKYt3+y0jJUjBtg5BuFzUkpoM8VwqivoLYlS4IOzD+z5OMyeOcAEk1BrYe/qhLOgHpZ1bohz
6BHIbAUNUIRJD05UehRncYlHQwnItgTMBMoYwtkiyL/RiA53B0YMXcPjOWwXCWqXYkq/S1KAljX5
A2AWAcw8Mli39IX+KbvHyJg70CHTAmAocTURzgRkAr6Kwv7c08AUe5RvJmncIHtqFUauBbtK3h2h
GF+Fk4v9BFCJSSJWbHd2jrS/TD/eHqp84u2shQoSn71z/CNieA8IbCxndwcTjgi9UB5jXB8HlTdF
BAWX1axp33wnjORn+Awpdg6my6whOCsGgnkGfD4fENTRneEE7vLDc9txrPsMuMBoDBKkFnVK/WLB
G7rB4hEIoet/g3XL786w4lq20tHUjITtalw9ra4vrPVU9iio/jwK5pNG/b7DZgYYMlUQqVpTK3Pq
5mHZQduGz2SoM0ZcVT5BpZhdl+OQjaSjHfXbUZX7AjHVod2/+0z9R2uo/RSPS+fvG57SZLPvoaW0
emxwKBE1g8FrT3LQkVBVzZHw0flL5qJJD2ytfL49G9Z5GSnQnsUcVvpzxZnOjacwq/yIAAeDH3Yw
Azp5ZiOqQDINPqokYYnw6GKjPn8rDrSlgZJYNIbl7grk93ylwSMjzMVIdN463ye5/mHWPQneVoNO
lEzbJfLk7teidiH9lq+kdwmCDEYc1FVWrzF18AdHLjAillO1bwRC+q28+ADBxauAHGfkx8JeBFdj
XyeLVOZv4YJ6x0xAE9Dxj3HnBlvBBzZuTfJI6vvlJu9BMQTRa2Y4KFjVn8Ijq7Y4iMXVVMvMI1Bg
kw1785hQwYMSKPlAXQQwNH6L/lvnxyPa6PBF8bnr7faMyTTw3j2I0h5/UwaeavUnPPnl4wm428XL
us8GeYD1f7Oe2+b+avqnRCzYFRUv0qVO5PUVKUqxXehhzUHl7+vpIupsQh3HeXlWL77c45fttB9x
tR/Eax2ktKY9KQp+XPOfgJBpiOMkViSF9l+DtocE09GqGVWCoAtWuIv3gYT/RRMYd0NJ79jbLBJw
NImkXRRK4F17Dm+kNYZCAAkF8rctIzz3D6APCFRYjY1+2M0iCrS+PSTnMJEs+DXvUG4fN2BMv5iG
6GmTZB3YahBORulSSOBAvmqflgJjxYRndfwcPARtoKjhUiv2WjVCJ7N02x+7g06KRZh/ATul43dk
vnghAqvgRy7v7og2U2MyeltdYAGd6UcegP4tnv9z8Jyau2n6HAUBz/hcdD533cvYjMAPtPasmnEL
r47AwrIsilPimsEH7qRvG78XgEfwY5DTuFVTVXfjsPj4hNAOVZHub8Y00L61jU77w2S7fp5xQPA/
WK3WhcTYHWz8SquxowacqvwrlPxSh2/4RruQNzqZJP7RJgnAjo5vry3aqUvKuQaAr3FMFEUo5vDq
c3WagL4qN6K+zc1NSIrV0wzvsMgu8vl2DpHourd44eD+TSVs1iWvZFUck23E5kq6/pWP8wetJK33
YIW45gPiYvDP0X8un6A1rkKJ23Pvz1Md8pvD+LkAQ6S/wxg3Utvb4piL4kJnwQloGbaI3MTf8gy8
dqZ8qOheB39ybCAGhptnmxGci8YFpf3cU7Fbmkpxqkqoz43KAWbPELGwX99qjmSHvgZATH5TLPrz
x8qjkAytEqeNJ0oJD9wEs7/tTJhoxrcnkT+mGKxWgl9CZLEDEwrTs6mzamfxgSCMtkb0YNAa5F6p
QxK0KeVxUY9+4yewCzDYGm8hruCpfpoOcTD4ZBYDOPAAlkfZTDoZJv1g+ZDZdFIB18uVV4PNdiIQ
IUKrF8bHGvbbR9Z0Dl5rfsXH63rPntxADfFM/646TfnGx5xsf7OaIoU6LYplvTYzjtIRo4H8Y46w
qoY+5GnAmcGdrZMsrZZVbwUnOkFq6qnsn2ECe9Ke4k4zzZ74gmeZioH6vzoPchhjYEtUfFtQ3sb8
Za5eKAVCpzKhIlehFgOqcXDPmQeN8LYYPCynZFikg+/qmN+kR+nS7sXSw2Wks+KePFu795pjonT8
RjaK+BbbNIj/ciIaScJTdXjAeyCNieoes70sO8OfB4f5abRgQZXv+tiDZqYDfAjCdspJelKVjY8V
dhFziGMNRaCAdryLUzJ+M4gbn0v3y7R+vimkuYoaByPfOXII+Z069cTF7cgS3vSBwPxwNmbA/I7D
8+HwU/FzpPV4Po5e+WPRcze+/8bPi2kAB3u97CIaF6x4OfijmpctvvedBoOLaSw75Nx3WKGYXQmK
aplqBx/e/GB36yPK/VTPGmIP87s+kPeCh1TeWQ4Bhzq9xi2RD31v2cEa+jwPDc+ymkZzsvJazVPh
jmrlTm9ovm1VQY9dXNNZkawnyVbLXwnRDG74c8+WN2S5qBJCFCQ57cmQUBPkNLRLs7HJV1hmIPaQ
zH0/S3XOtm2asxgev0AJ7297boKT8r2d5LfOvc8iIdhjrX36lHhhT1hbj7McXPgvnFwhdIODJnD5
yuPNgu4qyCaczZ5OMUO3sWkILvjJrpsch5O/OIlkqH1arDCO9jUkVyI8sbDDFZsb1Bi97dEAnV11
YQM8bqgBtHtBxk3UZ+lwHTLjJyNUT/8mzHuCP8HNrm4/hH4z1odjRAd6Gbkmm/+EXse3YwhLzs9u
bYle1tbjLpejS2q+02Z83yqucjb4f1rVehv0/gVLkQEQksOBVgt915SnYJY+I2Mukqt0O6gXO4yQ
jPDtgYCqISe2W2V13mqh4UdNFvPZ2LqfygiXuZ5nEUB9ZWJ6Dx1oe4Z9BbdpgWmnU/7tteoaSw/0
OA8nUhLWXQixBTBMUwqNDp12tsaPC/CD8SVaSKsoQ+n5RYhYz0yGUTj9D49/J//kzx6ZYHR/QNfb
3Q4/kbhmcWLw34pC+WOVoS7RoI0KHGkGPiJHE6zFqFOboo5z6yQI+STYjlVC3fDZOdoG4WtGkZzX
MO6qaJH3mqWALCcnWUPukgw4HdM+IQ+35mCW5yoqkNm+05S/Dl7dmz+dV6WYtrLY0WODzIxql82+
LvxvFcFYQs7X/OQa2f5nCFV7xESw9yW9+P4s4DMS9Pnu/k3/JvOTUMfcevWnZNstbEiVyL7IKs+H
SxnCdw0Qxl5xa+PNaO3bGefIEvs1NcgiaycV+D3fGne4RrmdLnypPwFfNrfqNiVHH5Tj4tEzCpJO
qjadA3fj9vi4Je/dybows3An1fbwjU5tTdBJylRoTLo6go77FCFk/q0CoWz4y3jZuJq+1gpQLxUk
nHf/6Ko8q/CDc3ln0n680aMGiVjBdDeQBKN5qhLmyU7v9rDqUcX/l4rjfMML+wio1BUux91SC/l4
IwfK6YW8UkBfgCSN6uKs7vR1U5TSqoxW7vVJX+xTMiPYGkVoHtCgaRXWAUCjMjvy/QvN6daF6HOt
XICw1ekJzoiVfxQHvA2VT80dR4jBi7/ng8h+UqsdpJj+9uk+c8w52IyaJ+R9uH23X2QimiOxgT1x
pPN/M2oFQNOONlGSbCZeCSwbzvKndShvPCRU9V8y5B+CJEB+rTbWN+wVGTdNMRnPQcN2SjTJpuD2
70MsHaSN8xw33mk1AtOPT7W/q7183wEtgtc8ySpNGjXu2ae/LKPaOny8p25hgxTrQmfb7Wo1ZDJ+
D+YWxeeVmopSFsDK2YQqOdRHwf/Ea7viJ56gUWziAAytGCIw9Z6dGFgdgTCQ0LlwGaph1ckc3F9P
Oq00oJ2pGoWbJzggNROG3Hb9m0ruh42aubpL8SF4cbhOLvKz5J8vYOhj0OADMJevxSPm0KhAXWf2
vzxr4gy8TKv7SyGSU8hSPT1HNKAR8TRopm5CszwQB01TwkPsoxMeFhRONyY9Xvcw4B2EyAkcvbOw
8pF+A/IhFqiZ039f0qpvqCGEI0Khae1HLPTtlrEzJV+FTBGxMdfXVbARBK0VK2lfh3JUuNTm8MY4
OhcbRZGkhLG3sAtqd1YP3KuFyKYNaQf3mB0EJykV4lq4VlKAp321zv71QGTp8/lBeoD0jUTtBxV0
n0QLHnKnMr9NctFdXCRjt6QrKA9+7vnQeALlfjoonbSl3+tj6TdalWZWs+IzHLecVQ9f2Wq1cz84
wg79/UimAzHeVfACYH5p8JlNVZdBL2uoZdkG5kYpr2J1Fc/HVx9WzAMwodHYn+mymwEErWWvPKOw
7ROAoeFS5ntvQvXO891KNwtWZYlTifRowh+iXAlQ+ZB0NN9htKEs+/Im9m8yGfn8bVoeoYCX8O9E
esgDPCfWlYtXFeqXJBj8L6Zfsp/zoigQKUc1/ZHF/Mrog2rNFcWduyef7hKOvgQUVEKRaetvRIcO
OTGjncdx6Ne1CFkddsyvoi5XIDWjRzDN29cQNemqpXrxZ8q+ncbGXRuiuITJGTbJcjppFGvYEfXU
ic2i4Jel+IOQAPMzhud2k4uMgbXt/g6uR7MBYD0+3gzONuVTVlJDXtl0OWmA8a+b/Hm1ZsEHywqy
zIvYxYlnGl6Ft3zodEbdHmBxWfH4mUlPUBdvwXG27u8iwlzdYKBzm27jGj06fPjSldAehhYVBg66
m4vUQJmgCIlo0wylV2/mSuZtg6Jsn3I2FZiP6cO8N70nncAjN814ErzbyIqgvVrZOeHnc8m+p3tA
7wi/ieixtO9J6kGSW9RkUdpfI/WABH9z7WZB26fLDSQapH1o3pUSI0GQAxXHqZOZTZcuuZyRoKKs
6Cb9yyaRtcQ8HBodGRPViaBbaTQ+MNvZsHwgVuZhClmlBk2UX1s+aSMhIakdwH63pQ/YG9Hbl9sK
3L7Oa0liSw2zq9dHf/ast4w4k0/X4qHlt+zExaTX8eC3sey+2K9TAacIRYPxyml3EQPFwUcQCYOA
vmdpZaGEQDxd2Lc5wJGFKF/paBPnleIoeSLiPoMmQkqUywY6nUgGZLrU2YcB5P+SLHCnOivBrdYJ
bn7pkY0PGf9mQl6I7R4XQn7PVIZQ5+QUDpSujwfPtWfA8BlXiCwEloEVlZSBLTlBHqCyMefXXzI9
2i2xTNgXoLKgKw0PFT0lQ64cdzszSuwR//WYKw7L8stFK6wEn53/B87DFjgZRMVwzHgsYMfHQyiy
sYYqKuNJdEuTy+iOpT9m8ds0IM5c4pg4XJKKMPlk2NNUtrEeZ7SahA4di/8DVbKvJB2HBWotdGx7
2RXKPI12L6yKaJRNycp4WqdKQMMR9Kc2ynjVHyf6zlUVYBZX93SOP8IATA6Mwy3KEcWS5Qs/ah/a
kSoHe5wyFFoaw/TFfhSdVTfQjOKwS4Vkgc/nuFqF7VGGOmeN2pmtSTyxqPWy6UvjMkLJP0cJ5akZ
ibuo3nvJjqlqwJmXX8PdRlz0RQVvLN9UwEaOcoT9qkuqKgnocZUZAFmOL0RpwUf/AaXFGwrR3/aG
Z+eTpYjCTAUM/s6OCDyUBzXjULCKdbyWOFKYbgSCgNWq823ZdGGrRgaYOw5czomzq7danHGImvm/
WrJ9ElerVpNO4Wqx39cqg0FnrRq9SQwJsVz7ywICiIV0SIFmNJlZwvGHdHKeQUogPbDCtBej3c3V
I67LneE6gQ2Vx5O0wN3cZUBP+7hAOuVHNK6VX60AYXzjJ78PZpDkOLHglYDPcKAK6yxgWARiEjS3
JmopBJbGVIbQGLNWV9CAJ945aaO3eWUIH/VClvtveirx7cAuvREdJ3HT1HU47QKddKIUwam/UnrC
qWLK0hc75W8lZzrBtzQ20rsPqAFtdQMcjOWXhEPvBC8xaGdbjz3lkejStGFiyg7bosJvRqt+hl6P
Kv429/v+PsomwPZ7jij0Gbd3XSQLKsvpCCQcWNLhr1Cp0divRZGM2xCnC8HvywM93iCXkqd49Kja
kcFuRsE7PEiTeIwF1UZQnON5nnG1D6u99F7rUYPnkScNO54dUTVq08lWmvJPzSBWanvTUNJ/w/MR
LGO5f8XAEFVT/AYPpNwVJsDRwIMzGNLPgykp4IgDKmWLWD3bt/jVW1ThmtzQToDG0azjb72j0gQk
w89aLfes29OcU9vR6ZRGvkx8aplzCcRc49/JPDBiquvo58v3/oy7c6zmDis4AnQjhCeDeRoXMCtx
XMo/gyIiWW1x5FVUNPy/qMkFLrEsVJjBlcpXdNg0erRURDpiWBL5hvo3bE+j4GIND3SAVorr3tmq
wyY+/0th0jjm9LKuNYul/DCCp0qcYP2iFr09HiO1X1nh+lgk09mo5xc4M1RZ4ZZ6KO+EqmHPWboP
gR6cIHADaBsc9LIMaJXDS1G3poUhB2BwMPEIech535zzu2y1ANDge5YIgnHbDu7UAdN0xDkORhpJ
w88M4LQLB52Ras2w9f8=
`protect end_protected
