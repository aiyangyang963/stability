-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lyPjXFW58Tf4Dmq+NqPXqxV5vQW7Owzg8m87Tl84xpljri+1dvmM0U5M0B00MqDCez5JM08Ir0X/
19bO6IdxKuZiA8jAdAn/bk6jvc7zAa+YttUfYAwjg/xDntsWZjdFAWYSKtPvlTwt/7cSS8JkrKVk
xuJkyUHJeDWyTEb2RqgLgmHCnaB0BK+WlUqvoGnyPDO7JVaERqdxizM21r6wmLbZp7U9SsW3Wt0o
lXkVKjU+GCFB0wKJ89MZuNalnf7YBndgBkkRdMvhyhDfqnmnu01Kxerc294BgQpGMDCrdrhKejZb
RVp2BxXBhbuW8Og/MTzQWtXT1ZljaNzQU1tVsw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
yrNSow/Sxn3M7JoDQ+aQeo2/vg9u2KgCBzpjLaglBjk6rbS/tIEFsbFLvqcrmnxRspQk3xEkNnhS
RZpfmaLxyxvTJRe9DSBxHQt22wDqaT2wsz8r15DSEkFvwJ3FkZ88Yp5gmA2FLi/StsQqUnVKyfmZ
HTF2SDeqw69YLFUiqxrTKBsP3dlYYXn+Ica6+j2Vnup7Id4AUgIYeJWuTTc5dJipXDdRUxK1yfk2
9sopYytcGClTDHtSJrDswMrAysa7ywzgpLsFnLz8zbDq5KT1K2CTXW3nQfBZqfxznttqeKUgPdLH
7g+KkBaLi5VUXGl4V73Pb8vTePfposPSQmue1IWduMDWBn2p+d2+dZ64hHEJaQZx83aRFE8rS+gE
83c+ILyFfMYeEniKTN2JZiNLFerQEHwQ8gb1MDgOIsrwJdHwSwigYV+YcxQGQ28xGKP6Xlbh9tLe
qoYK5aoHX4LH6Eq88SdwBaj8uJXYDK5gAhO1OVAWvHPni7ZPrtuos/j6uqMvIsdrSqJ4/HuWgIAU
bk0jEKA+doLXiFtNNxSCnzgA+PilK53icZnLYfItgeSdmYytaD4t5T6G7kBat7B5WRioGqmjmYvf
EXx/qyfePopLiztPyfHXcZhnj3JBpyc1Uv/QryaVAwO6YWu/N5kk5qbh7VjkVLJYTzxQe/33pmZB
jyqGPRBJh5wbmoqPx0S8eQGJUh0/MaLveO0BvnLWnzs3BsUOiiW+LKz+i2g0FHkDiUCF/xe3ITzl
U006l83d1Kqq8gQd1YhlKphk+H1b3ZIfxb1iDsG+Mj0YdMRbEJJj+9DizyfHS3tmFZINtD/7j1LX
bHuapD3xcNJ5GQG/Bdi71bsEQGo0iXz9cuYIAEjVgc/uawqDQr725RPjjAbuE4awJ1sRUWh23rhz
Gj4hNE8O6zL6HYIj94Hjr0I3wFtboxVvjH+mvC3G3iXn7mPiNKOogOJPRePdY8JelAHx+U91YFXI
p0Q7IhIdTsR5xMROmFV8zyCKf6UW1QU9iBF0UnIW0ZvA8o3qejnT3YgzdCNpAtJPkRtw8P8n8kfR
m8lqYLP4grctR7LTtkh8ma5lBNzBlM00p3Lg8p0ufWgnx93duZZ27VEsUwuDHyQJrtUuyn+2TImG
cShFJN7Wfg+z1cTQsGqNHWXzFI6l2Y2yKYbWqnho9ELBrXwShCiSyqgOy/DEXTsnf00uTo0w3vF8
mYVBCg9zDawAp6ZrmlPOz8TYd88/6m2jd00H6F3fKyrSPcsW/0mhjjm+aSC+Fickhzz2gjVmH2X2
xRYZj2Jk7zRTCbXvRBcil6QFFgg6WyPiHaW2MjfRNZbPsASMcY+MZx0lNWQx3E24gvb/7IbssQTJ
5JkqLKT/9JjrI01yu220SfM1QBsQlS7R1JfaHG3DoXNt0nvV8LuVLEw9tpkfFyzP8VRAHNZVknfC
a6AJie48u1rwtEsP7gYde63WzxQ5K/T6Usdtpu/mdGlt/LUlJ19EsxaFlAeun8zAeA5dk6NY+XII
piQspwx3gEfP34+g9ri++ILNiREN+kQwSGRqhTp8mT1nKKmqsQeDmT81dFeC8hIYdrWvOTNnQl8q
jkwsA4xpUFETngQrI72qeehGWNyGaTxRNxsBtLSMd+VdW2FXij0YzwoCNTGX23GUTm50A8IwWKjk
Bsf9dUjWkOmCfhLfoflBBP9jjfVG1dIlh2GUZAG6bTJtzHF56MzxeIQc4AeM3jD4Uzo8zCdJzHFz
AGMnKX8LW2PTckaULaILJmbV7lajtekBCcVlXItG1fVsPoyi61fCuqCKywPRFrazlERUlgXrBRLA
l4UgRS1ZJHyRpSpPFT2HGIsqRgrYIjacjJ0lvyye+2OtsjAIA4T6gqFMqceDsweJg6GwUWAgTD9T
IKokmJgshwuT2qSyNV0nFHNrLt+huEgnjEWDkEvSBwrjMhXs0oCjr3B2nUGBF7dYoGbqLS8ywqR9
Ye8cEHmOP7/xElXgryvaVLjGtMc4lJhGeHrH0uM9Wa4Ilcgum3E8WOYJsHEqpn6CvpLDBF/YYTjZ
Il+AFSdR6ugeA3UwEoio5r5Z9KuBNmbJjX9zTOoA+eGeio4sY8eeIwBiukpDuVEwGP9khrwj0XHf
Kp5Lm7/9SY+biUK5mRyfqayV1LVkeeRCCagVSOJUvkzebbjfWwPXL5m+ruZmEvDFegISGMqmOxJJ
Xlzcmb9f4DYsr7Ii8AD+sP5auRap8JgO+HJ+V/UKkESvpQ6/nU4epCMhAVp5fRluzQR8L/W3Qh09
lXal39gE2JlngPAJoTc83J8O3HUtZWjkMEmaIiKnQiSEYHvSIsS9WMOrIxzMNKun22wVKEz6HLER
p/Ul0XVFYXN1ulv0AYcPhmOq25mtY13joiFpKLOfawE9ZFwhvsq9B+vhf4HVFmLvKbc0l4OFTWSV
fXl3OQzGhsAe5JI0BCIYCUXUWnyO9ggVef1U3mVqOk7yjIwGp9PPIZY3J6qlFwGhnDypc01V9rz9
wcSfLI/QoRYxJm6vySHEKL9n9gD9jHh9EL4aXoox7aO02oW+hby9oUlwsqHNEJEKIct1MrIGfneS
x5OXi7i/DeT+1EZLUPRlFhJ1IAKSGousPlsDRr1Ii8H2eOSLr12yq6TCFD5x32hRQ9ItwSOdyhO+
iCqhOd70VJzo8nIxHqcEnrchYepsGZEQsonvIToZ7d8oAhXzc8X+4ErW2Dib+s5AggLkQihd/FP/
poaAchgDQ9imgKPrs8JFPIW7ju0+0T4H2t0kG9sfRF3jAnHOQCKG7Zh9HIJSfjTbak2MRJ6LDAeJ
Gt1H41VE3keWorwJeEUOH4pnh7CIxGE/VpWK2DHdsMFwUTYYBbzT9uQG4xmQ9D8gGW2MbOmHxLug
RypkAyk9mPg4/Ulvb07KG4a2r0zJZGxeUh4V7oSW3pR4p8JITEy3Tm7iAZ/RGNZIlSkDBYc9bqTy
NpF7sQusT6ZUHkRcLYc2O0gWRvvk+DMtgnmWhO0au/nK+qOOvZqdhdf1JHMgKTGvkd1AhiVP43H9
GZ5MeSqBYqwiZswvHgdGwA34twJAcKUOhfEIdMIjefIQH6/ufnq7/z7SHhM9pWADowh4zWSaSasg
TQzPfvlE+eu2jmwvKQG5+2BGzn6n3Iq4sZLoImwTGhOO37EIYwyJWXlV9dz7+d1MCsWd7tV2fz8o
9aJjqgIL1oenVdepl2Zo09aRZ7MxkPAx/2jfx0qWJxD8yrgFYP6zZ/PH2OSg2bVdOYelWpcYQUR0
LnWXTVL4eG1WHR/93d3VXQsLa7oRTIVUKPqHu+xmoBtdp6CG71OgJSOCpaNqEz7ECk0WosakEkcD
dfiKHWORAEsmc2imxyQtgvEn3wtKp/MhCnzZvoqf8kyQM7quSbw+vI+mFmdt3G8IJjvJsCT4FI+X
yWnjhLrx6OXyfisoo7za0jOzgB1RMk2RFz4okjKDWIWtJemAXyw/lFXxFABEwR995cKgJUFSVlwV
DKJWPDqQiD1O4y1omA/TmRn2J+8J00S66a8E/+jwJA9NLSvXq9NcWRWXANg1nHqqpLLvwERoXo1X
ERQEiyFI82dMNONLeOiGq0jN9vfS+chEhge3mDb5Oo6nhMvjELGATFpNlM9qlRx7MKuFqw8bhBtv
9xcVWjBWN5uF4Zrlp1VgVZAWBV8Aws5IOmkRsK3Oy6e642LZJjAwDiwa0G7b0VOto3nuEF/Ney67
uSQRhY3ZndkBH4Zsr6k3I574UN3h9dRymiGISsh5dIlZN1N9NSK06CfMtWO/1BBM39X3dtwQf6yn
qgQsgSI3nJ89ojTE7ZBar/XP4xvAh8mKmik1jHaKiCoZDPGYHcKnV8QcPL64VI4FNOh65/UbrRvp
bZ29CNYOToZNvTy1ilJ7gLFT8KhMkaqj2DxMCo0GtV4Ew8qPMB64wtr3PRMlZiHUAsTMroUgo90B
Cscd+uxTco5DBOoKEHSrwzhjRXqPP1zDVHSLLwvEBa3GLB8yWoS9UdfDPL9aMqwBy5rQYV2lfqJ4
/rnw4GT2810WNWydJ/jR5X8XYVCFbV/hum7RbjGVsIsJYX18tBiZLu5X7R3Sl7BInAnVh08VZtxe
wJeY3+dzxA7OdnaxxVV1qWBJBEiUe8yj0uzOB6AYOlVuUWacnZnxLrYl+29pr4kOcgZispBYFlpK
6wa354y2mpvZ78yJDRZ9Xw73wun2kjUdIyvrQvQG8eNVLDMkOn8Sp8kPTzXw9XS2jUEtqcCqNX/B
djRF01+SmjVC+V72iZeuw1FA6h2Ma6SaSfo4/yCmUzFOWpI4TJGoZX2ERlssi7slKbhzqmQXc+yP
2kTdEp2Otq0ikyoENHSNP+68eMnJCBS+GiXwh3yx8BulfhFyLrLpEdghKftOXY0cuacIwZurmVLN
OpqbX6oNfkQFkm3i/RBbYwzXodWwrEKtFWkxJEQRlp9h7v40PbnQ10RjU9aw0Jg9Q+xF8QCXGZtW
kV0BdBdaAguw6xqCa3WbYp6R4CPLdnP0ogagXG1X48Ax/SxMR5uNgRUnip/jSddG9Zn25NiiI99A
rGKzgKfuBKxo1AUdUMpncURMaaSXt2rBUlZSOFDO1cPQ/yFQp4COdQFOyQrEAXOkdbwOqBblJk/N
4HPlbTmXRXR9V9Nbb/UFhg2L9Lf2XponGWwSsmRlyT6a0yD4DRrM9aQ72WDTOiXN2X7N+zd734gd
TgHYjOUPxVIQfI/VBZMdNT9zWbV/SQ7uocjHy9c2X6G4JIzldzyALCsaywKvfKQnBFrf30E1z5dR
6xCbPcvnACcfcuVbpPnrK05+OmQYOFAYuvwBaI+Zk/haHjoyKB79374w4qsnPDvnUMhwXX10cw8O
knHoHzA5LJ+qPaB8eMC4ng4zL8xgXkQlvmgbBVPsQfUKG/PAg5MmUs2eP0yWWYM5vrItNeGdC4YM
JHdcE9kEEhkyM1JDKhIyKaPfrR0Ocvkn2Qtiua2EIWcSCOF+AWCwy7rUnx/pZ8iEmCfkTXfNZNgW
NUVWldyjGtT1JPBgIcxJvWuwpPXx5wzqsMqI3UqkE3PPdYAhggGBBrCn2RpnXelHbNNlHCL8dcbr
zlasrh6T7V7z3goJUSIqgiiVLApgtk4KTpG9BLaf/q1Gva4eAOd3fVe/b7b4s0Tf/wZZOaZuZfpB
kz7OOsDasv6rcquDT8FZ0TjDzvuFjcmlL4NMbY8n2oSZIaZnwpjBD2zHCLk0FibpQeeSv7gmPBF/
TZkEvUvMLX+LSddbZE9o1p4j3yXOZOUrHmRhDpntkqdP1WPRfGyRkZ7nW9f5hQ8d7bk6EVGT0rYQ
fVcXiQXaolbI354N/wh0IPg5VQ/urQKdpjstpbL0zLpAFCqy1WYuTPgCGrPS7RT2UQWfrZk8EItK
ZuTXo8ythDxkfZ1v7KP1lLtntQF9MsoOfdiuPRX1WtI76RWC19UyfU8jkMqvUsIdf+ksBk5YPX8n
Pfv79eY49mL1IFLO3ft5oOinIFvO0Z9skHA2udXlliht+S97PSVDdfpV/onYgOgTFX6+Wk29Y4KQ
Qox4DcI/d/Pu+GH5oYDKx6SJqnFi2qh+h33Xy8UkVSm5b40kE0JP1m366C1YeRJcHnzRI9vMiHyS
+Km0IfgzMdWYNhb24f/d/T7e18xEV/YXj8lFYek7apoVsIeFX1qvczp7i6VMCAPah1OvqCtg/G6n
GOmT0koovKvNc9H9bqogc15iO6O4lneaAwHJj/ZXV9x4UkwFh/LVLZ4HbullF+SZXpkHRnS5bmN1
WBX/UCOagynEKw7RfNlIo+cnBWa+uH8EJSaOn+5FZV+S9ieF4HiD5iCKsA8WcjUOLfKRFgFkLU6S
kWn8D1uLf1dgIE3Zh/moLW16FYrReKMP9S4RGlKOurvcsqw3JeQlGNlfasDhOgZAw2sNnwLGzoKc
WaAdyizYYD9RQqsLtU9zL3YdVKxfR2PNQ7n1CPZW9Rhm0wpcSZd7vrsRUEAtl5sF7L5DMQw9YgRf
CkTf+p9+q0mbGCxHQXOcFhiJUHYUXDCfkuPFE40dx6in2s2dPtpu0QKD6HZmo6M6lLwfd5MaRCE+
Q0YTW3VBtelplhvOb1gCpghzumn/Y3KhsMtJ3HhfK3QBPj5wk/fGBCQV0jJ8nV2t8BILvZOs3F0p
5gurCeMKxripBzz7tJzcOIjN46/cIGFaiSI2eIsxf1q/gUBkvCG+czPUck42wcQq0ofPqxV/mfhh
q9S/XkG1WvfGKVhNDo6dsd+aV9tz0T/P5zCrCCGTKANnyTk4coA+LI7081Cv4os6amGuTY+R7hxr
kSvsYmf7W6sSC2UaGyebd+VllRN3n0g8eo4UjXs4KaVnS4leqoLuR0aRJoo5HJ09clZoV0d8i202
Cf1tKXi1jpL0pQvxO54VwbD85BouYc/BMRO89LLigADjX7gdzbHI967ykZfMIWE8MNAt/gYJfFfd
0PRW8FreV/Q+1i1G9q3cBdHE/y4DRtkW+5hxhegQj8vmwr0/2lN/zKhsc9jJCCwP+z2T4FauXzGf
MJsPH8Xq5hwCQ7FbgBk2YG1qKE+qDFUBtS6YKe2lDya5EOExjV7nBgU8cXlx9KJpcA8UWt48Cfiq
ti1Sy/a1CEe/zsrx9ALPcatstMsJ1a24fcPl+HgcXkzTRAB/7F1HWSj3VYDWspUrc6YZKU43c0ES
1sbDgJlgX07PjInCdIWTI5Uk7bxbu+u9K2itEVfS7/qwPUdarp6b1JM+zb3SbSEDG6Vg4yFuyf6t
hhRY8wJ8tezoGmgKHL/Z3kCQW6Q/Wp9giz8QDFgzMO6pN1zPjWe/2kshA0ic8aJQSxbTBtNjUinn
8sE08gt7zccujKmWArIf6VuuENd3+qYEqTWSX8wABGT9AHO7EN/lbGaoxjNG21FJ8xF83cafPrf9
4sBru//IJq3o+WgXx5rDcK38W36cKbk09Dn/uYGAUYYp2nwVH1rDcEZL92+YK3G5y6xu6lgy5yuj
bSjv1jIWXzn5qVqox/pMJndF7Rkkcman4tZZour0lSyQ97fzO9fMXB6xqk6+JA463x0QPr4+XXrA
7HMvFrYkYEIgt5xHwoPUIh0JBGWeyBM1yapBpUkXpc3/iJ8ar9eGsRWOvaaRYehfLMe0owHsWWre
9HgIBlvYRLNiE7GeB4fvOHdKf1tadzkTwqoN+EWRq8TwGEwEzyP39fKTFr/Gi4LgCs3OyC3iQUzu
G29YRQvH5O6AWV6zLRifsHg9V96awfggZBV8yR3Zz61zM2e7J1nxiJMwdjVbrVf64FuMbqrKw+ar
gPBkXj3Q1yWLChinAtyJkQrvtKr9jSvG0+XpsBbAt20uQ4ytu0tGDbtvJ5Iv8jfN05jf2JDznbP9
o7bp7jMrv8pKVVAX5bYN5wgTSNvLZpl0IumOB5kFaa4XJ+xdxigW1LfHtOVNnmS7X8V62TKncHci
bAY71v/oLaB0EFoFLXlBToBi5ublMkIiRqgMt7NQGUCkl93H7uP0xS/TxvYnE9hTekLRA8ITgkOr
wh1viyQ+Dq2+Hwwge7IE30ojS2VsQXRKXwuq8lgsum6I3vGwP8x96XoqYWh4/hoDsrFeqM3o4TuI
bY8s6XpZHotAXfRymo+rMgNRDiBAMFAEavVLVNtKLpt8qWGEo9EzaQTg7rwoHgVoWA2aVaFtll9n
qfLN7aGg34+XQnoe8isRs/7vsi1a+qiSrt2obX1bCupHjmHYaYq63RddRMqYVXx9pos6ysFmZGoF
FWIFgGC7aFRNFLRNUZyNVrR1Y8Uln+3vF+ZEv0GvqfadSKQ8CX/6SM1eKhyImzqUx9wG6W0yyl8w
e5u29n9WB9ZZIUM68/wGswfWdn47yqdxRJ5BvVHK1XNuExZU0oc6fDT+VZ8AsOYCZbd0+uX/dObL
SUPbtw1qER0+E6hKGG0wQNYKixjWjuXHOKzvxb24tZM8NxE5/y6lSBZSPwC2aJAqon5TtBEx9uFV
6IYvIfMzWT0ZbNhDYW6KGrzaU7rP0veUs1Vz//MUv8NEiDVS6OevV/FT3MpdZsQk2ypKv6BedTBp
WxsfLuTGUUXcUS8x0viHWTy3ks+F/DDcgxpyw0b1vVJGTe6KmLGubb6ROMyHNXk45piyjLQTYu0a
LCZJ/751e9PXh42Kn5d3k/eBHM1Bu3N/NQJ/gM8gKQ5MyjPwjO3zlsZCztIw0YwxuslvWy5MJqBK
/Ob1Ql091SgINI8nQ8WPqt7kiec6QScrFeezZHJM+Ih01IUVWBxXfRbT+6qnSkgU6Q3kTv3CB5ns
zqYdyQQGiObs6nL5IQrqPYCZWMqVLwlUcyWB3PNwbc6FUuDYSwNJ0inoGU2/g4+RS+4ehkrrmRad
xa6eogYY/I972kqeaDSX4i14KUjltUjl6jDSaGw04HfQkPW+dSukLymEm75+9WEmkV3mFIeae8OW
+POByEEYMWOHJU/mMXiqTU5R86Ih+0uA+nquRvoiV+xJCy3jKwuVhmqDe6bfmeGJAKXW6kEeoQS6
MA93CpquQxqfLZyXZiK4T28nbeH9L7wyQrD6SD4NJjWTy5fL5JL+NwWkIbgB7t/Ytvi7djm3cr+O
OK7QuaEh/o/Tgl1zgmYChlsHGz0yOKarU5Gx5WnhASPMd+0y9QtDM0ZMz1xXBJJOBHgQudIIoFsw
YB44wBCaLo95nZp61Q+tselkUrNOZPRTX36jq/gVUtb2SSFelpFrP5Y/irpApT1ilYnmHKx9sRmB
bxby9RY4zTCAsbCJ7Itcvc+F+DIaoVRgxdCjSuL4dWQCyE1IGslEOBpPD2bw5vvpGSOiLNfw+dw5
bhtSNu5/u1ZWKFYLnZctoYHHuZlHE9Tg2Xqlri4Tv5gKWrxUYilJe7NtGOuGs2BahTO0Q26lemAM
V7paREuQnokexmZgjjianS4m8o1gcObrn9Ze3ibW4ahLVSylLAuASnq0fB5fX/xldOPyY8oJrVir
nlPned/cYqSVafS1ZBKM4z+HzW4GTBdNYmieM02P/e2EjGB8irM+RqEF5DzOMXX4cW6JAF4ww2Zi
/ebnrQLZs6/ho9akjr7ibjLHG76kZk/AJA1XK0a8g/8wloxuPgS+5SoU99p8WfL2qk8pg8trlyYG
KFLA99xt1dZpbctAC7j/WRUKy/vv3DkiyTRMKznnFWjadPQBvj5ooVbLTcqInvOwlTLKJjDxrs4e
hg1N0Jp0URkZVd4Olgr7r7uxWahpAhht+CrSKkVMkIqNSMYdLSENfEjcwEfLCvdp+7xi8wGFcLVS
8YM/qBdO5yUG4hIho9hbyee4dppaZRZA91qxoVTZKYgRrzqyKiNE38OXG2noxRP6nq8J/NSyaoKU
XvDmApjOZoOjxiWPlqWrq0vaVvy0lbjWykWHQuFkGdmrFjcJYTXnLLtFAyk3reFij1glsQTyfy5y
A6jvifZNIMLebQamHHUK/jDefTK7YxY/hYsHejV+eOm8wnAyrl9yBTp4sI6+GC/xIHuwVUuf/JV8
KTHHGp6S5r1YSMACm0Itlx5UOb2DKR9emCZKSHtKZeCXxA2zDNMUqD3iit56d0cOBmKi1h6h/JPL
uPq/KOwh/DInmANK40vinp4OxcKe9N8A732VIrJ+FtVGZAWmmZ/wT8g3/6+KQAocdAdbT59e1kOr
p5q4zfJbT3YmVYofzGP1LV/Sxd/m0AvS3g4c7f4+1XMflDIUoUKfMS3TVbJ1IzvcgAcRedo70y/s
mkRO25/tY6mXU5ym7Eoh/+XgrPmFxi7eM125W2BA3fErfgINxSh3rpZUv2okc3ySFfoZu1nTpKcn
s3fdv0dqWRVcQmWc4qbQ4DVYiTmngzWarZWBORAg6E/sXtTxivNc8BWYE39PHgOS/j7/QbhHLthH
1STD48l1Jl96+EysoJw77WKIT0K+So10QVNWIvEfh/B/sxitHep1pKe/mgCL+48WV4+iBBhJY1aQ
QPfDVyuqbZ2HYbdWCKBnBcPObeWpsBSDsVReMeocUoZWHXNDrh4CQY0UMbDrr8oyOjceBinIB4+I
2ZyKvPd+J4zXyGNuM5jtln3rRuaEDBNNdgqinVg2ymBj0NmzMiKtIN6btpKwHoiYlAMBeXF4geDe
9C7P9MKSobPAvT8SHGZsNRieBmjlLGk2lmgSueRIPrA5t4+NBc1yUjvBhyQ2ANJUxLQ9l/9YXyGs
U/pJdhdbD9k4LpxcYa7CASDCIeF2ss89Y3kxfhUgMj3bj7Wv8Grg26DEeidwXniFvu8tLscHjFx5
I1wepHWo4K9UNDy9vg9mxaw368F0E3vMXh2ycawi0bQ89Ma0SPjyACiUMzuWIdjVDvhqe5EsZN1K
QW++pYu7dgBKqSyV4N+MAO8JR8dDzQnZvmzbKp9+bPaJoK2qhvTb5ow0TThD3IIprOyPhS+Pn51W
Lya4LkzSAgwUc3RmAT0lkLibQjG+tlaRRT5cK69TBgt8Uz7FIgs9n19LYLo4J+uYgbrNOQb0Acyd
gXtyCrERvx3qynVlyT1XhNj78PaXGyDuBZouEARfW6m/ogWQ3FGXZjihrfHAmkHrwsGWz6kOOhJF
B97zws2mw6hCXCg9uZIRsZUqbBQgwwLSO0SYALijrg5dRHwoEEKeY6yAbqnHAIuq5E6i1hcixEfz
GIDEc75LUJ7SHnE6zQjGEMv6y7ppKGUgPu6I9X47qkrRK3OnC8W3PZA++39tAdvmoVXJM9Dpx6eU
GccyCbGbGwJnCE0t2Tar8snYIqboPp1md3XI1MNb45QH4KCjCpvulCBvfpQwazawU48/cR5oLRhq
CDcqi06eGejBPuN9n+ms/u1PsGqvUM9AixqFR9bsIpt9+FVfNizdd+BcORO0ZwlA89bR5gZDjjii
uwWLqm3NAXJ/lw77MI9NF208V5hS0LfGy+do5pixqzMIkd1Pfwf70GMvV0HN0neOsoSj+coSTeOS
B8/cMezZYQTO4ZKms3/q2Uxb3ehMo3LWj6SI7yS8KLk9CTlhCMbsyJdpTUnYD4wG21eXfrv5Wqib
4wpwM76Kred1MNRdW18TNc0+vTXdIoIA7dI8caN1VAuN5SDOQmvT3PsahanD8q5JEGgQ5qC8Aftw
wW1vZY/hwlX7tRnCV6WAxzt3A2pXDzzgmjN0RvzMD9PhTl+rsCLZ/Qd0Qa7Cy4OomTsr5xqFeQiz
Bccu19PUmiJWuvZeN28uzLoRDDjE3TapxGY8zolDwT+Cngksz1Xum/Yts9q5PTuvPayrQYEF6dAM
bByTc/NGQ1Mzmg8v83jJlOXhU3vRNXNKVflE3O+VTLgn7ojL9OMg5JcAfXRPHIGrJwjUYIHr9GDl
eYFAW729WGgVIZlqUTMqFPwwFuHi/V2vZRdFJnNm5CAuoO4BTXhAGP94EWQRJcnUoSWrXXO+4esh
AJGGyyCyJQ/wmOF99MQ2wlOZGx2BWZD9TRIsjkgr+j5YBDCTazT+PtF287ylMixMdrRIw+LDh+mg
r11pPP55MHJGpIY6UQ7y1o00ymAjWgy6xCTqJX0fvuM0gL9MiRYvcmZ6/uXKS3IcG+lvEf0szaMJ
EKNjbsP10mFw+VDPK8J7tFaGmGyC7hgfvMABO9olrTglAS14YMU51zi8iDpMPy/755XxXzlaY2vb
5kblMEfCmcSXArjMbKne0AfSwEY4L8KI2KOSL7b4ywqiBIOiix+wYWxQk37s1KDclCwvqmwiWiy9
U9M3y0nbi/begdQFntudQeK52pPOxV4cHMIUWu3surqP+x88wRNuwrOaoOLnHPZIcPNuhswefqlu
IkGosC+lzXwjHb8wtC+fcsGYv56NJdmaFzwboVqp+9ERBv4N4w4il9YCpMY2RndG9ZAQyF4llHMs
wQvp5szYuepzgI/n5UAAQveb+mJDpZOcr1y6jjs8O4v+w/6hSoZ++9ch1WeqeHV7Y5JJ51X+2Brw
AcH4JUL7b2WiQXRUZKPfufeoG1BEMqNd0MtM5qLRbeStzqrqTDo8WcqTUc2JqZ7OI2XJCpDhvyx6
6rhXfRbcgaHbAKFdzkxPCPgiYVvyt+FZu66isMp2wkMo1n/CX2U09N3UjEcAl4EmNJTHw2vULheN
ZcFrYnI4gO8hh+qQxFdfTzTQoxjd0cWxUMFztV5QZQ4mHDPOcyIbuOrT3b4WPKyx5GjcXXq2BBe7
oh9P7Terc8Kn8zLQI9jxNgTorKe1AcKlGx+AGxlvJEpuXyy20PEhXYpog89KhK9fFNnmEPta+cCp
54YgtO4dqwBpfaGroo3D6azmBDlAxew756JhksGHavr+2XqdXQmC9oqA1GgbEROsuiJHT/IGWgHT
4haIzRUHeGxvbOinQQgORyo228qGLj0X9lGwMGgJt0frK/4Cu015NEJDBxfwouBYP4QYHlSdHC5F
gQk50xgOz44EzT0qpxfejY0kkl1O+32PXX9C4G4bAJYcF/aw/VJLy1y8t/Ath7UxANbzGnjRyURj
XcbBj065pDfR8oB7AfT3cfohMYSsIuucXpRYXjaVfeRQRg9CMi4gatYqDS/LYobeb8rQ+/CLqVPs
W4c0qYBwpMNWE4MNRDsigiEtRRN2p5q5lnkPxyIyFlrk6gXQqWHGFd3hYayJ9593xAZMDXY97lNZ
p4Y4LIXN2UqrlnkfMDp1rKO1dE5ku813n9r4hkQ6qYefyOGojWy6vNMCgc8dbPpXcmPGivjnLgXZ
PvPyxd2WHImKPo3W5KLziLmniY8M00UyAPPifHS4wQ4NrC0G8sU114jcl5mMyTOvjaKTqstoIJQ0
a1sPJ3mJzfdIIEUQ7Rz+KciYVFa9snVcOVNLSEvqPpPzaHoB0D4+mFhUmG8zMA7lOkcCvtTuNHrR
gw/DZvVhXMZ9X0fSlnrJ9yPOm1SB4Ktz86S7a0xec1BY+29NMJagFCchVxGf1uhywl40+ufejMJn
toIG0SoNQxTa9ehqjJta/m8idoIifDG1h+4jrvakyZuEQHWJ7HuKimWvMQFEjy1IepkYvYOsD45A
DMx2yMISOgPXts0XXITkJCa5MVtjhkD37RQ9CLjGomFo4570OVFIxex6u42AjMSRcjzyNsPXFhNm
iV2FwxrYO5iN1R8BMqw401UYFRn01+52UV1w2ODG26Pz3YebAdJIRFDwKL89ROZDs4AIe4euyvmK
ZtVyAlPqmAsrrdkqARstJUI8xcNQwQv50L7O6dgW/yQ82qcAhR6i6P9lBS8AMDg1IXRB6PgK+LE1
LDKwvr8HI1+GaRv1pOiAQolSSeg1K1gqP7c8ZYLsGnWDRWeNoSpcrX+DJ5AksScLXyBLQAfznBxU
/Vi8UJMPHQUOM4CR+GEzdOcTVmafgHoU2W0pswM3nDqS4GmuU5V2EH8gh1GnCzbAIJgR7RnSqk18
jKboIviBH6LguM99s/ufCTNVYeO1wthX/wstEOQ/30XYsu5zyYkaTXtoufpDrqQ6JU9wtQlYkenY
78aTVgibURzwiRlhxZ6THqDXIZi3Ndvy3DxEaBi9q6uMrYmZHkhIoGgVFHZ2QGiHp4xrlB3iKL19
RFgFqF3/GJKPyOHHt5180FD7vFK4nxPbjM5uS0MHAACgv4qFE95ge55BV/28MvEF7CyjmEjByNqX
TsnJYqqGBBf67og8vQzwvlTgG5Y+YKEQrR4VTEpiP0b3uScUvbREHm4O6RKDuASzgQCPs/4=
`protect end_protected
