-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HmccyoAiXm57DsKM0GNzKl1cKFqcTHPBW6+JNt8PhWfsiYP9USPcWeYwlB5t6B8vhxfeXRhoMz7S
/VPXvBOq2D7rkUh0+lqkdaZX+ftohueqIvzLkK2sT+1j+VrOtyg/kcioMuJWtI6t+b2Fem66kQSL
abzn/I0Przf3hJQ56o34Un7mMEGPhH8dY/vEzhvWRMXTlf3MJBl+SLQU+8M+U7TZY0eNbvF/zH6c
5Ku3DQjZFC31wPUicEhSMQUSnY3esBXneG7RC6Hjv1YHV24H24svbGVg3FTBSff1BM4vNCKQ++5c
E3AsuS70KfPCpALMQkF/27PAjzkRFqpUaqYaIw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124976)
`protect data_block
DAEK16Tr467OtpRKyJ+KvO6TfV+0wIyXSscV8miY9ZKjF7GDTxRbQdfkYfdynWLer7De5YZlluhq
OdAZxIaqDHBjWNEy87JfNtjo363+3LuCIgGHtX+wLwm/4IXDEDl7f19IH9gjM/azTqgBR6fnk8/G
yUEuKgDD6twNqEBfCJCm2QrVDdoD5CD3pZBcxAo4WheCA8zxbu5TqHySU7nY0M7/MDBwbkQQQgC+
Zp8Mf23D4to9Z+ugB84UmLK67iwIZ+ei4CbcGBrRxsqxBc+0vpMLH2235Rzw3DxJdijKQyDjzsDU
WAE1zczmXjvcTZV8yzytYdvxnGy9k7uzoo4PibVIL0tUkOoIDvXsHZrw4AoBD+TMchQ9EnPPyrnk
TAXgPkkyaGTbDBYK0JOPwwG0br5wel1i0hONJ65Dv2icPa9Y112p2Qm2E3qS9O88w8/nGziPTc/P
XYu+z47NmvcSjUNm4FjW3145xRNa/KvRJXsq4awZI6e1xvBxNkMvRWna2rqNRq9qnViVznt519R6
5xEoBX4ehOzZAOblj30veoZXOAy/PUSNeX30E+vHvETwzHu02YhyRWfyb8a4R2mSlLoZhpZ3MKvm
QY9RlJp7qmF4vOg5ymfH+lw1xi+H7fC1ASLDCQXyu1tYr34CI5q+F1tylSoDV51H/XK3DkjLDqlL
uU4hfUBJsIm4vRZ/CLi/BQB3z/Ml0/sBWiNBAryPNLLcBbgKeGa8WwSYZzW92P9M91iR6QIf/kqY
c9FDLFiR8RGSu3lfzK4JbhnL0qn/4mPZw6x/nAp328JwMa2Ne0mePW4m4pd6xuvMraqez0V5Jc6b
MvC5mj37JglzADqfMJ4gsceI+XB/ymZbRuRyjDU7LjEjVHpgXeMElunAy3juPyiEmLCEl/D7w5Lt
BkEYNw8Uu/8DyorlF1UllcIsAAvpMSnGa290wnAWJEljJiwiZkcPGLLU4tRcmA0n9CoUStQyI22h
21IXwY3yBjCHMoK4f37gUFGI0HUuO7oLlcMYx6kkhGcL1oTLklTWtUP0FJVyG1Qdei0U3RfpIcvO
kZMhE9VZNelTkd79wpIP9AvyBkCVXS5J96ODFyYd8snTr8aRG92K9NqmfdFk+JaTYPBMhXinSgE7
r5U6Guw9+yCp6RIwHoD+KwvcuQ9NlwQmfCHR4k/rLR5I3lvX9Edqr4nk2bvnPpRhe4yix5E7QPEn
V8QC2rb6Z95yp0ATYS6i/kVnnkVetVmHXC2qYc7rXR07Ktd9gFiIm6YlMF2L3zUrwU5Uc5qyZ1lS
PQ3o/q6ekGqfnCtV7wDc3ACYBpnujZlHSJD3tEv/n0j2iNOTM/QMyuthaDXGhANoSdVuWI6aEGOA
T5nLQm43eexAhY5pY8TILqjmujxx0ij1Xoy+RROcYAplV7Iu/HRCKPuYySi7Zn0e2Vkt5KquZYfZ
4Cg33Uu+kHBA4wg3L4Oa/U0Wof+772JneIwceUpjHpgmbxgUyJ/Moqt9PmLcbFghQ4mlVRTpOtRw
Qeqge9VOTwo2qK8q0/ghskAv4lqyE5V8xecLW2UUREJs30HueCnT3QEx5WbzEnlJgkrCYIMW7jRH
3HTFvOneP7culKHLTOPBnEimMDYvKFXIXd9xkEExNrJ8tlzLcHwqmY5tS+byoZccM4nD/Y7zj7OH
BH3BM1C84q4sjNxzl2y3iDRQ7Uedn1yeDrQRpmQTrEk4kTlGBcCKjp+0qwIucJH7tIkGg1cEKFuB
ufU3q8B2Hx9wQdlQ5p8+ByilK3ikmGq9D2XwrRtRrpDTKiGA1bqsK2wMWvit73PX6HTKTNoO5Nuz
GSkM5QakXhHxIFp0dRwfSYOCfdxo+S1wlZ+Zctk8mfv0+xH+YGdmIwyGKRNoub8Sw1grxpAb0Ton
3MKitkglHhkIcDF2nP2NlgHT7rAQU+EgHECwhTSDFJkexC6uuPfBSi528RvWqhd/wrkonE1ZiU+o
JX1w1B6+WqiOMH6O2fSVe9rs+JuLz6Y4YBBNwfIfft6f4HGGI2JIGavIKjHkLhHxeEhr+BGTKflI
o73Su0LH+8ICDoWMAEwsSypU0NXqXKHP41/xWygVAvxjphOGnB6uDqS5LevhFRbbQknKEHOLuF+b
AZhF0bUetrGQaYbtTSyHgmM3SG6+EGuO6UabVq5oJuKrikqz7bFKJDvryqOoxHBPBAVcU9lgBe2C
+c4SIKTfbwGdHfyFj6oUDAYAlKYlUW4sgJUofILhnQILQLZE2HkAWa3TiEIXbsu7Ho/9UqZ88f4L
s7PJ8sYzesBcSyJxc7vexEOk8WtnOqIBxRwJ4A0oEhY4iZW2WOUA91Sw4bB0QAFTWR6d7CEoOmom
DP1TJJ29IE5y1eLkb8xm+vYtT/+TZWDR095Xb1e+CWeV5PLjbAoOiskqYYNb3quU3KdKVrMxcvZE
zTkQgS/hgAs24ay+CEw11UCS+2/CRff52jYNHHP+UwZMvRSGpoIbMDr1eB0OyckNCB//H4gjvhy9
E0epeqsmHWU/H1iiONL1FyaFZLN4VNNOvQgbS3vyAcQg5HNj1U4GPWu3GQf5FXvjVOdzNBSqrlW/
JuC2NYedJAITpOWcDslhx5PBcIR1MlonY1yE+z8geDDt1tM9Q3ui2CViD7Mpq6zkZSsk8cMgkIrC
L5KSzeZJhX+1x/ZT76jwJt54SeuiYcIfW7spzFuLyQwtXDCFyReGQVHx5MghQM1JHNOGI/f1Mbpy
Yd6xvsRXj2KNgUKNn8A/xi0/Iae7jNqfhSR0z3AHXh1EKR0l8YMZt+BBJuPkyGDDGOkKM/y6T73h
2oFceFzsgQRJXPU2jeX7aShOBq2AYXDjV9mriuCpztFViwDEBICbaJUTC7K1HcRW47qHpI37IMUP
4m6AQlx5xUYR2GZ5l3vDBSHG43ppFPwbMy7+4WxTtdH079Dfa1VMXikA69kuys/Q0LDpunJ7Z22o
5KTIaWM5jGqaZVUr5KEftfP0veq76HD6y3oNVwLrO5qxrIVovo1CbqZ/DNpSbneQF8vS9ixBzi7Q
trBA6selQb7OBHXF8sWOuy7IVU9hhBb/H3aSPSrtHdtBrdhLCQbRM9VoZNc7opmaWaTsiE8C7eCU
FsxchwnL4VVU1A8r5pYvN3JBdy3bizqPLl/JuIw7j/v2aS5/aME5ogQFaaP4Sv+TvmSVlkGPi+75
sGr5AZZUBHn4jY3UU3Xr6Iz2imoDPGqwPe1H7jcw80z+bZkcZ9DjKQ7JzgxJIheyRpgasfE9FrGb
BkA5ahC0p23isdmrMQ4z1HnORo0ENr+SJMtspmVojFSIv5sy3jPmlAeMZic3tpwHrORTiqBok6xb
vXjv+PRqf9PvZRV5yjzHkuutIrV2laogV/eGYS6epz+VaDQ/zmfrWP7QhDCsUeOXeEEk1JmuYsGI
Vo4C4V8nnVRR2rchOfFWjMIojtMXHCYnLc9+8QRU6/T/X9bU1aH93EvWycIEJG56QekAW+gMonJE
KfGISV+ugSLON46pD8qmVC3aU0JixV/9veXjKMuQ0R/F0OJHDC2macD5nm2or4kMYuxpLzAlPOQd
bQYTEGxRDXg8JiP46OnfWmFN9MfBem9WeITDdRoHJVjZ6wBeBAdBFTuv7reh61PW7vrYRjl9YJy3
UvFt/+WEubal9oN8sPtJBCIGk7jcEThyrkkBFYduKAblM2gQ1dzXIHAYT1ddE8v+Zsg7jjd/qWLN
/iN+g859dkOK8xKOeqY7Idv+4Ucax4PHEXA9vnC68vPnyGHHLdBCwJhaKp8UCnOy8SH3Sj19RZ4v
Jc+8E9VaZbZZ2gdPbok6SK8YmW9SFcd5DRS6/0ZcAgsmnXf6T2fBseVergK9z9d1te00kMvqxyie
klv1BLeGdBnLXqlKWPmZAG03uJXR0VGY5+wPpSySGn62IcfDezPiaBz++Z983dW0qZlrD4CTZQvB
gYEITCr36R7cDOTk0UtTbdc35ASnagcNIy5aZ8Y8v8PI4melsS1JdPDvECG6BfOi1NSWxraE3fqL
eWyNPYFrO+FepusKKkPnSw1moESNv4qaNjljyFgbr80siye8ghvwc4+6Kbe75Yw2X0smRFg5FAeY
6RHfbinlVrtBVqYPd6OEoe1pth+jQW+THwSeHEZYP7589mD/n/UPaa2ch6eaARyZCQCe9GQEqjaa
s8PjSxGmwBbSRuiIIoO8VRPbAC/jHQkOLDctlcOCzwcSydHfGk+rHwFlGYybRr6BVqTa1bX+h0/O
T5R2F5QVsVu3cHc42C3C9H2SRn+EkYFqamevvWOIkn+zC/kFOuXC6uDrd9CUXXqhuRSBDiD+FNNY
okM56GSMluGc0+/eVNVqKpfLSWul9NcWAk/HGeFil8/c08jw236qJhGdoPXJbsxxJVsIBeSQRkFx
VKwiIUMFPnR/JIWdpfB7xZ+pzy24FmP9zqG75Wf0UpmeNBqPVcLIlq246RkQb0b5XI+5gtI3os2k
4SakBdl0DFkW/n61ft6zl9WaHVOnYohO4g0LusXhHUR2jwo573BQXOX+Ti/O6zGsKrqhlJrxsj8e
IHx7evV/o5ZxbWgSGL4sNMc6oIF16oj2pDecyLwl/N5RxFDph4AZVmEDMMjLsb5HLAcy09Echl/0
1YMp0jmNh2SW4n+WDV6uKahjYJrqub4YLJ85clVbYckmYgDwoo42sb9aGMdgvQtBe0rFTj+Vq4pG
LAvD6X6GQFMQfQ7qvx4iDln3e/RQNgf5CTZYcml2pXxP9jsJfdisSWjx0e4v1G9h9q9JjF0EnssM
wXJKYTlZaFPsBuh6jEMhIKEncRprUSYByquIJvPTwijC6dXNnDqYjf06qQhJpzP/4MB6mYugpnTh
L3B3Ybhcq+SmbpKvf7yBag5zJXvVqMCjAlK+K4t1XYVTxVMblOpor9ekpfJlqqi0a+XtAI+Vtvgf
KgUdcYG1lToK4MUofBsTKudBKV7/ZDyIxG+Y+Gc89P5PQiyfVpYOAWJBC5nz8LXGVeUVNFybTYdi
pR2leLYva4sFaxBpxbLKrY49G81jgsMWpSAqNY6EEI7zwI03BNUGQMP8CK8OFS63eqE3823tcJt9
jFCfJbJOUGFuPFgmFgLDmLyjyd2BAnLL3j1B2Vvbgu+meBht2bXMmOiOV9PgqWHygJzN215pJLnf
xAb8MPA3veUjmgnncmIVpQ9IPWMpC0MkR5aW9k1zUMINEi/6OEwB0nKRrCWfgvwwEDq8lKqcU9Fq
gQQOH+6G95kGmk0xQUGZ6pmiL7hiDRtsqlc/kundJMIko+1oFr59ApAf1i9ClDOk0aZQwwAR9kt9
LSlqlUzb0ZOxLvsYmNlbSslMIk8TFmhML4F+c5GtUYnRbOreZkMup7/ovnV7Dq/CW12jNuhKT2qC
Bb4cOA9Te+D99bFN5wKDGf5myqi+Q3H+SXwMNZn2ZwrCYnya9YcgZeTnpK9RaOX3NucihM6ESUWS
ufGwWxf0d83fAjTbWgDpM9K85vWyjjl+myZ6JjlH9DwN/uB3vhXGJRHJIn4pHmd8UF2YBNHYE2sI
dr/L5jTWcuJbJyW9AlVA2VEg56ko8sF52lLlwnf7nmc44d3ueUbuRNqnUWMcdo8aysZBgYEFlIbL
JXHFcwSkX3hk0/YodSzdGDlY8UIOcPcXKdJ0U9vNCkA6euhc85gD4f1L6SXuSe3GtqEEBLBBeon2
ZMpW3uXILdrfMyqX+QaYRyz7ZEdZ7dQKkosuR+JfOhuPyj/801emfxJH/9tp3D8pDi8p8YlGDDA1
YcD3tQY/M7jjKOpX6Fj+UxusyInl4EHXUQToAb8WS2ZORpT8BplSTLk2Mp0hc0YlwfZV2wa5cdQk
t0eYBVcYJoEoDWAp79U1vBGnM1s0hN7uXCOIpiaxfTXDW8wARGsr724c7sLBc/o6v7Btq5GYRNsc
8n83FlONdOVVAmyrQKoNzQmxXXZEzsOVGi24XP8BV7h1kySeC7wtx83gCv0ClheBoArOuJhLic+v
yijlmZ/alpt2TjHaRs8lI8lQx+UH9eBll5X2lR9tsUrWy777HQLb/m3a3D5q0d1nERqW/7S98dGu
VN207yBlR/m3pQzcKhBh2jy/TSgjOAAAisjvuvtluwQ5TCZdMeBn2m0A8sbAVrFh1d2T57Tpetlz
WwXhQX+/mX/irJhNdTIABS4nYNlgfb9PBd+oGJyhDZxNhw/OKB5t4M6s7mF0acVO5GeFCYpNafuC
sFUpJjslN5tvOWrLLIm/HIAQLCmjQGgJi3N6bjEMazhoCf5V8MLm1ibDKL6A6mDS8OTuOPydtGjw
3LWYiFdbjSYQAQLn8qsBo21UU3yeBMjiqlrc8oEaX3GOO3jViCx8PqE06Wpbum80VNSMMeiyMJaS
rGl/2LJlw8N2f9ObXzDEMzhh4WNQavUX6sjO24tnoNiNwalJPlG2tWEtnH0+U6om3JyT8C+IytKw
Sq7jD54JfuPTYFy0MGacRXCQkilnTqwLicbxv8J4rVVPSxJyue6hNnDuLHCNE8rsPIoOPiLZZ1ES
heYvDMiKEydxwXI4qj3t1WHOuOWmM/eOfGyfY6qfDyG+72HWGwsVSOCjwJXXl6FC5HzB5AtdBLQf
6SjtaxhHq0B1x4u/ITvd836q8mdxBv30A+zVB5vNElwnS2OgF9iLhPM4BzAwVlq0NTrR5me3wToO
rzdBld3A5F7Z2ULgVKSJ1fEF+aqi+LjkeURxc7S0jtqN96oditmYQLit9XTcJYLpDlZaK4HjH32i
3HqaRvZU96rMKQGhAET+i/wD/biel5cRwMac7P9Pk0pGAbnDgHfUQW6r/BKKdXXzks9/NJuoSBl/
iJvmV2wbR+X7S1gRnrwO+3Pq0JhtjGknad4Tler6PX02cwt/wCmYTCYRqV9httCQh2Glp5N6Jdz+
J266xCSidEjfgbTKpVD2ikGL5vC7/yI0d6Uz8cIBUrIBFh/xr+mi6CBTdsVT7Nh3VWj9oBb4N85p
0ekPk0C7FrnOLun51BPUH5JDA+TYEDF2vTB7Oty6fQFzotpG1gO1FPIJr54Wf5JW5n2o8+iEGmlg
AEhpP1rc9Idy3b0IDK+i7pG5NCd78Y6H2tyeJH1gmPCFZS22p5W0DfOetnQ+ECL+VZkrKs8sSreY
/OqqU/D5lBWwdEyiQaqFds9+KWmn06VEsBq3EDEGsDprPMT7s1Tw/mES28mdkCs2SvgTeXHVTlSr
vfyrvLF4KyZICGjrbHFwwst44/4SQDOxwc9jBT/6VSslw/Bq7P7ke+loJFJ+dCSe97NootIsKoEf
DU/YQnhedqWMrlpsV+LHTESUUEie7lfdCcxTocTgj3Mt5zk/QIjzGE6eAR4Eqf2l0qF/tQikThoz
ftzIN08ZghMwzQ0PCCTaK8Y7o3OYTikE0L+gRJHpRNdGjRjM3V2MATzCCcGSl1ghV3T9ajvvdO58
cVUEiytK6h8h3kn4ieBYmeozL5y7DspvgoL0tWMnFHtfqKqiRadLuODo4OxjG6xv1rclkDdU8xQa
zeRLRFHZyzIh0RIpQGNwYfclvLHlbVmOraQaowlrktN6i0BfdlKTnZQcdSxrnFd+AGAFDAVxPGdq
8xpdoUrqG+g9yVzpI/3xNL4aYhN+otDScczuYB6XpgnwNSbFp5vqFiGkLbGKuYrfCugC3drwlHJH
oBf7X0BjGSTQ9H3PARCQg5WpmbH/31F8DQy7CsELo5ZfDE9/tIhZU4oikH8Vvab1r8Ji2UR0ryFM
MVlA6lRM8TQi42OB1KtJam5V1Ru1iq6ZSvZyeM1fFUGR4xoCOqthRHqMx3/1fJV9aFynSN/uEgeu
I5nQ5+qdT/Is8rNUbuONOSkYCbsewVj9oEbXHlQy/M8qAIE/fQwhxQRCuyvG2/amdtiHjAGWlKrJ
ddu0XvtkSuBYNMwGcaFTEAzBhGj9V/6zTBy5BnE1ICLBxfPHMZgk8HXDjf4ftTHOJaCX6Ipm7nm8
trrvSayH6iLkwpejnMhgvbNoX3oBVmx5e4gGUNs9t2YoSGAjIFqYoaWYFjg+smuLCM3ZJiqbA0ph
DdV8XVbuqeiVwTSXM6SEWA/Inndu/HJzN4cqwkhGkvJNkJgUznU7dZDw3bKkevkBFo9NXa/AVLYo
5Zk99H1VesK5dnlE8/9Eju04h7Gt9AdapxY4sSmkDoVivW8IdykgL/b5JgaeWA6vd0w+Xk3I+1e8
fv3E5OQfta73VKhMHPLTgNeekMoI4FoOh5rWJHxrlyVBsxtulqycIlc2ebjuSQyHxGylq5fZqLqK
MsQScw/XwOyhNrFN/30PRtgF9tkwADpDt/vZc0byTSNW66E30KNuNUq70XvS7RJrUIyqckwqBCNu
4+B6ttFrbeiYvcjboB+WZxPMk6LdfM/r8jb27zUb7ihpdKnCC3vFY7m4LXktTfUm76M87b4dma3o
N0pIV672b3AxnG+70lpPFJKkfGSjyaJol3ajC3wo+tbFcn/6C4B5vr0TkABUpYkx7nPw2pjVEXbV
IsUmqXUchiCtxIyuYDoR9vpu9ykVcWghID57nVd3tPmcV5fPbKK2uSNU08YKZotd55nMSL3gXp4e
/xaCvj2RB9d8k4b3wZX0BeUfhaZWhlbL3mJhxuNsWujbNOz71AOpgD94JvDOA4A7sjoLtJG7BUEf
ILMxWfnUlIAyY7FgxGMx5R9rF9/8xuiJUgTTbmEL+eq5asy78/TttxgtgFZSKnYP8rYsdUoq+59J
/NSIOTWQaac4RHfw5JaFZ/QS+Qwx1ol4nx3bSEgUa5RqdQKrOwAt/eJnDXa7X1w1NT7UM1tRa15l
c+qsG6sGZ2eP+cmLdN4fR+OupPrpZFxqr6WibMdYonhvPQdLnr+c/X4ESM8dT3e3GeRoPwJq1f+t
bvwe6lCH+5ZCy8Z22WNvHBtP2F6JiO0X9aTLnS5NuTXHCPH3JEKC6yNR5yt+tRKRuwrICrCxGGQi
goDoW2RnV7UU4ssxxev281aPd2g3ZcA+DqF5sD6B4WLYomfH9lV3qXO0lePsb/oi/SOgvHjYiATq
Y87XJt5i6O0vU/qelZhvPmJVlabwjWCTW3DZcFS2wiTM3pEN8ADiH9YwIZJlfCc+ws2tCK6phuBY
D7rjQxKd+FJ6Xt5VcpV4KmIoL0+l+WUgImf12YEM2pi2OesIJn1ef432k4RltUR7JIzg8yLMYiuC
WHFuyedancXgTxkxEShuf08yeV6zAYbEsbvl0ljBAVzvUkWWqWbK038GBQYqc0DTF8WK3St0OZmG
6f7nTDp7DbBpxZcU69GpRQdcNkTES5yeqyze9STYadHIixUSsvLU/RC0rfsBy6dtqyfNRzWzJ3GB
KmROI0KTPPvnasIS+IgQ8FgquJ87Z6mtBSALvWL1Z1ZigjHtQQ4SmkTjsvhq54dRbF2BeYRhmBsQ
WPUUl6kc9oE7nG2l8trIi3gjLGaF4a+zlPMg6uS5v7XLYq42rVftoW/fV+LjA6qBUkRqftueK82u
rg0sLXCvJFirwzbXCopTLqTX1+4DtWNXwSAUx4o/jNQa9pQjtpT2ht8bNHkugxC4sk1RD4PsJ76C
j9E0Fx+C/xfMTGWe53ryHZFV43mkWOBQmKxTjo7pDtJABg9sQritrq4UKgZnQPqbeksYnavEL8Mu
uI+YU5ZqKyYHBIW0MweaLWxFw67Pa4LO65Ebt9FlWlYdoed/p7sV56musKG9cra4vrOtVl4aGYXE
JmH5ox6idVyaAwyiNA8/4sovrbM4Owg4GVa1zODpADvf0N3h5eT8ETlS/YepsfvCOY+V0xNW4mAg
capJkDVcvnHZPIpQHcKnm6hYYIXYH3ya9np13idoQw+z+yVeRVSdDRVV9EUeNkS6DDKWlAcol5+S
FzKCD61BE/kS/JRCM6rD0IHVJx4MQa9W4D5JyAfDm85l3+1hOulAP9+X4eWMSf70YWvbFl0b6IJa
kixdrNATIQMHX0ONNe2nLyufxj1Q4LcsW4NeBcL+LKu80gO2K4fHhoQxc3CCwP3rQ7Q2YXqiC/JM
wjLmu04WP0DlEWDbBYP9GK0fiRpeiCTsUMXns7qGOZ2WPz3WTFID1hDu8JyUPt1vrlAcuMPJcUZp
fY94z2cv4HF+zgRG6fkQiofbdkt5GEVxEI9zMmUR9/XGdQD85HaJhqZtYe/Y7/Vv7X2UVRFn/HjO
yGz3Btvd5dfBrvBrBWx4VNqiRH/rCIe2a9ct9EmCG7xIcj93NuI51YFUMkfSqReznSp/ccgmY+2E
4RiTmdWs/Y+7rTopyvDwrVPn+72TrYG+bOUJLhRkZ6RdCwrJc2zgdRZ/lVFgE15nRzrArVQ07WWs
HaH/YEatZxnDlrwnTDXy9BU4OJKcDRhyZGlIj8G9gfuv6srClzLBOiBf6RTc/62Hl4z13C8z3QzW
ZdyYUhJamf6pDy5U5TSYyRsaGJDggIUcvvM4OY6SGn4jQH0McBx29Crj/8FTf2j7ZP9zvs0apG7d
60K8zdMkG0IkQG/Ec2rIWkCRLlii1Y+NmEBR4KpHKTc+B0n6XRL4HTMYPyZdBXo8t7xh2T5+97Xl
bTcipun8StE96H0TogvIiokdveloZnbpHzpfZGkb73CKfiebvQLWZvujyNI9v0ap5qsi89mujZXO
+/1H5sWZDrq9dnjjHAGiBt/cwoBJPbtxDuBx7phSaMVUGLGQj39jb4ldNGvBTvqwPvIqQHOqNEbA
Bvs2dU9vJNY5GSX+4rqXD+icVdicndoG4XmrhOIFvwqTPiKQASKwrQIuFMlP3NAsj2Yi8uG6RC/j
7JNTjqRKzr1jbBD6Nb3aPxXOvKhHe8YSpj0Bpy5iWvafOwYfqHnrjIiP+gz4DEupuZnnxaEQJBM1
7fNduzfF66nqKIhJBiGeZgUt/buFVz1Wo0hvTFN1kuR52+KtAJIzAZnC045jSLxhuFgcW8lXjnP3
AYy4qMK9Z/7Lq3mutFVxCneWcjFbiUWIYGCKm7pwwSFLmP0Qaqc1MNBBiZK6gj2I8iCr2rekTLYe
3S908rL8XWEw1sHQwP1yeoXLSEpiYo8kgdqaIIXDApImcoqEfr7665EURKAONUFN3sXvXliITgsv
g6CQIoOb7iE/WQ7EcopHnqM7GRBrCtp+ETzX+XfegLx2gczYtKjO+pnYhtZkGPTjPd8YmK/+Q3Xg
GXEabqKfSyyqsA1k8etm2i1cROZKM+6YayX5ZVI16a//mdj7EXtwyYi6yFC2oBcGrJWdYKhR1GvU
Sooz33Dkb+GyHvyopYtz/HnnjOeoTt8rWP1Nr6SVp+KgYkY54AALDmgfdPAX9TcGdOfNLn9tZavc
mkOOB+bX5N6SgXC37KnIlu0TAG5RkyIWNF7K4kulnLHOYMukGtEsubBWXewftjHvlEs/Iy0Ss/fa
KHj2VHJoW7+QfYJ4/0lQLkEBfPKt6PYBYzR47TUPiN1nK+mlsYFC5dJ6k/TI61mF2+fDT5lp6hFQ
UeqQCQxdtKx2MSEY9pA5A+vIxi/CBc2zDa2CKKJr4mDbb8ad+5J8yDDqko6QwAuL4GLUFgnufkJl
pvhQSP7Gj3qA8IhQjjndcxQYPzxOFcuBsk3OU8bu04wy2xfU8czNqWAtgYftvoDePVBCR68tFCIM
5wYQtJj4vLUUworNNqWsj56hxnhSQAfERowP/bVifSkSoqUHG3WkiqSRC+nT/cpbiCe2Pz+cNXCR
CJXmg33URbCsA5Offst08g+FkhF6obCrpvshBCtTombLE389myiE4sQdRa47UGP+A6MFDRzLf+uh
cvjjM2mZOvB1EWwLClVdJFqb5XZLwQw+8HEJ6WGu6YmLqbWspkWcXzFg149FSpdSvMkkb8FFe4Mc
WduIBwAI7D9JjqbFfVKl3WWR+ClBuYEpUE7xjtlzMrcOTjlQ6GcguhKma4FtMw7R0Ah0FxX9qPRO
HBfZhY0Q1rzVZDGCOMuNFsw36CquAVmvXO8CIjvlcJmfd8wk93L9qYugDL5xC7aYJ7n3V75Zmgsx
Z9hn+0fvCjcmVgvz9kLy48ZuUEnhnax/Xj55dsZpeFXhpIyRxzKDI9sUA/GvGwYeB/b6k2T9iGvB
OeOm4aaPXpCg8ktMU0kgl3ZHd8sD0bhj8bcP6QAhNRslBNER/jMxrmVxtZwl0kOF1fbDAa8LvuE6
y1emInmwSeM8NattNxXen9ZSb0M23/VZ5AP9lkW3kN/oqlzeOVy028RD51m/0wSCouVNrg6JUNFj
ouDK/O2nqp3su57eatAozuAfExl34D8sbi1eMpLZy4jsDMqMWNVXW9VxkA84eBFnfeuPOwqe2VA6
/UT6dgAFaw1d9mWT/j3YVShqBd9pokwvM1sS+py78D3zORDwahLoT7FIKpWhESxEU/vhxlSYEjtU
rLCAy0VRjgiC7Mo17LO/u9HXxfZ0C6NtCacsTbHtRWW+iPuBcUg/9b7wU0DWq9FEb1RMJIvzifKz
msOU5BhRl7aueWbjh4NopyRSALQse2GxUvxYQzTDNv2Gadh/J0rIOfVlFn/QyqfXlmUbRzu4f05w
+jhXv10LXq9MvEHYgnr+mKVtreTAhM8HGSUwvHgzqpLAuzwfHNu1Qf+JE3jh/6ZmnftjWZc7cDiB
KjUIUUIu64TM/ea9kKwrp6gUG3tSbPwhe3pB+7EYm82OmfNDoGfjHlu35c/OYZj8QHLaFF62pSLG
Zp4w4o8RmVR6uKlVukIJFAIT2gdglX9fb9j4z0unmfd4QQ8TWpNw0IzqwuBc+N1r0iY543SstnxC
Og1ujXFcsIrPArSdWztsjZVOmM9+qd0EoKVtiFKjmBoppDpSSjI9wUBj+mhC5clT7i9nw3cUngtg
ApKHXt9U4AKnHuLHq1I0qN3Q3rEvc1GDE4AlYG6k36seFx05lToWUXOUVQpDJcZctWRuJRUhFUOG
6wsihItVx0sy9L8SO5QRO9vjkoD9SgdbuM8wheLLFuZUSM+s4efdXQmBBSkOFK/jNzEADWXzwoIW
ViTLC7i3PV9HempZuLJiKE2Gluu9FYdKUkfT7+qAxNIprL/5wTxQ/UistJ0Q56jyzqgXXnLd5xc9
WDyZzlw9HmyOgDHFbbf1mZVbHrU4TXn9FHTexMZ0vNsHX7YFB6Ig/CYayYt2q1B/eCOkj7bNNEmh
6rPz+UT5FYmbvX+Bvpq+ewGT48KwU82slM5A0CpUkVqzt9LkJa/CWvyDZaoSkT6d4weukFPC3TBU
ZUWe3AM8BqIMG4aM0zPxH07kllsH/F3UdsRIaCis9pzVIJystL9UJQbRoDV6JFka+1sivF8GH2u1
svUu7r0AZ25D4O0C0dbLo0656gwr7+sEmKuu2tV6IXCYFWKKZLOjAj9XpWa8FluFEiS9N0XWpsGh
I99h7lqptsVCt0+0KyxZekNECRFeyY3GX2mRVMbcqD7B1AH1kicMZ3rkSYwyOviGMqbCoSo/5stR
6CpCVcOn6v3NuMEom0q5JsvgrhNE5qdZCv4JNaATB36fc5vaXZ5BedP/NeRVptRGtZdhmEwTJxws
ppPFSa+50cu1GpO3NxlNZN6WfR9kAerCCYmrR1JFW3WqM33c+AzhJ3bUt9RTk72auravOXvWZIkg
HwQHt7DJLEgJ8D8GAr3k2tPYMrI8ustfm7qL7QCQ54umbV0t+SjdRyfTL2ZKSKKdzldGb509wq3s
Lo7KGXyX1BGlbL93KIlnZG315F+/aYwCLhk+NVSwNuWCBnPR20sfF0I63G6Y/ZwsybMBBK/9jdSe
1hBt7bJRS20EFwnk6J8Id2hD+WNMy6bESl8HvFZqwgFWL25KhwnDpSynrdl3FgojGvsKRqUVkuUb
pXCd5IZH9Cz7hYGWC7fpVQBCnutUWfbvm++0CnLZz/0retamFYOnVLvuwl0rsr5uM90Hx/7zyRnm
huU1G+IBIlDoGGOfJLVVfWSo0+3QeQuILUlOs4rrBu4nCO1ZDymq4nz+2H+v94Hmgor2zYg1fnBj
l6s5Py8frgIJ0DyIcKNq4m4Ky8Ol8aYKl2CacDz4gSD5D+JSYNhPi5ye1DLeMmDddzEFRfplDEQ1
ps1o4NzWCVMNduspyxWEsmPPzA1hLjVIz2zrwiQThr2pXIXiMs7RtzjTd7D1jBHP/DIpSZEfOru7
sgO4z1zu1QepF9ClvO3TQ+KUJkSXAyyfyYn+LAy8ok7fpGb/+QwGt4gbozyVqDFXh6g+6Za9GFCR
gF9t/kfHQeNCSmgrgs3llSeaB48/7FlkhnxG1D2hdn6raD45LdwY21rLBhRs2Xn9Fr8ikjopLxLe
dhpEUOvUzJUY79q0YiGMgoZ8GEO6AIYPZH/mjXcU1Yegj7ZencWgMOpHAyVHFa5/7oa1m+3ar7vI
/Ykyuxkyla3KA+d0cTVucii+DTLK79fsxcCRuA71bNWp7d/qGx8X4M3XaoU3+a35AOzirQYMgSt/
WVRYTJED52Ia0xtCHDf/EYCaX8xTFxDU4cdingvBxBdMoI+P5+9P2ExI3lxKs3z6fJznJWvFK8Vx
UFCGmBnD7uFrpqKabjdEL6HliIG1SxK7DLyvZyjZJ0wixB5JwlQBUXYxXOewXMybU6kIxf86Uyxr
RjLfVjsOi3Yi2dZPlG40v4fjyZYoTKzJvzC9yeaIJdRhaEdhiy83gjqvoKyRdSP0eT7WPirv233M
ARVhiLh8J392+U5nsrexCvVe2/qFdSnkf1gxGsvI2dfHd8pxvEIG/Snua7QIAH9drPYuXTBSPVO+
1UY8IAZ/REuXYCjjE9xMSd9IDPar9sOHJdq4yWknJoEJkaYTZ9HW1aNDYax3MVMBnOh614zsalrX
w9Ep30zxDOiyix3MY2o7JLnb9mllYw3LwEX8b4aVuN89ECjdo4hVt0xi3DYPAFzz2BeKk7HiU8UZ
RdaBiRPhq7rhcf6PBDAnLz5M/3xmacxuJT0oltga5luxvHBfNZ3OH1NFfDgQAE2LZYheKXev/ulo
Gdj35GwLS1XOkTNIpbvyW+Yy/o7mCZeTxOZFPzj8yYoPJxCNI5cqdTV6MOhJsraBdU53PJYq8Hq9
azZ7fDtElBpKMyHorK5t1v+iz6PMo2Q0rpRrH7W5n5sIOo+o/tHRw6jJqrhzg9pkbvbK2ozxVGX1
UP/PKRumuGk/ELCQ3hohcQnpTNa4o/DyN3PguqNztX3DFNmX/x4YyRQE9Bs8U6r0uLAKW7MVb4pe
1AnPzBmiRuI3Z32Nc/WKqgooB93cCpVP7F7IRoQ+LC3NB30FT90O05oEPEz3neX9M1Gjind8LqAc
nqjymKT9A5OQnw6gzT/SnNAFiRUNmr9ctks1Ots1Xz9rgtfZ3FoNKgqCH94MDjDPSMi5qYaGFnTV
0/a8YKjVWW85v97HMSIh71lrXq6jo2M356iUXonZcjNxT+RqshoiWlftbz7ojJko8ymAZagcX/uz
AvHhz7eWMWqzLvXj7bzQGGwLEaa1DpwEY0yiqDJgi3eLrJfNwt7As0yrwMvqbC0cOhFcI9S3q61j
T37+JaztXWYPxH6O1Iq0oGNtNk420wGs0j2xzDyn2UxbD1UCqlGKro1ZkVMCkMh9l+E3KBOsrgja
E9WyihcvPJG7N3FaAClwwGb849i4XDWBXFgjfOm/H8+nJxtCiwHMATOt3NSuHP6Cc9V3aOkuTnDy
0KvUSsaDMzBIj+TMAjxaaG2jfra1OUoJC0FWH70Nmpz3FChqI/ifI51brIgIv9JOUi+13snComos
sYK/lthgLUpGEEkuaWQcC+/yyC3A/0wU0qeE/UZW9IUn2MZNV+p/aggn9eY1dI++iMrAA0TH5BBZ
jEeVys3HcqEw4gGOWQtbkeCphRoaDyU8onb5AykZwBQQIWZTFQX3b+eH3rOVW0z3Na2mzAn7VgcU
xJASS+M0RdszNHsn/AP1rEG1SFJcgoyGAf3RAMf2fETR6FxnrPxPOaF/flFRvTmAht3RpJEKo1bb
54kCfOlcoA9QuqvTTiAjZvjZU6llZNgQgvZAfA9GJFcQsEQl6y9ZCJrGM6VF0Xl20tJ+0GpsFGUU
rmCJw2d7Ce/+Mcv6N13SMmPV68j1/zkkf76FO85SaDZdyiRVljbVlTvnQq9OqKcbUJqpbrUCjisf
4/QK5vxppJ0LMEVntEGil47bWMNsqdoPpEAqiKldYDqICqSKKe1M1AmMKaDMt6fPHbOqFOIz/98q
TLY22xeR/eoKJR8/UloUQ9GEHr4HNX2nUO5b+cPebqkZMZqu73cyPvhGZIywXIqlz/oPlVzAybZ3
tkmNyCrQicFo9KzXdNMY/KtIYCAatqCU8Ig2zSiNT8fN76AMjoslEUBb8SrNAS3BXRxc8567A4dM
NMxbx9yl+sU8KCjpBlKNBWQ5ihxq20PN/xRkYQbBBq5GJJP36rdt0khg5iSL+UltUJj8M3jZJV4M
Ulk7YJ3voeOjD7O2WMRWEvJHEIn+BpiOF2lU6KJzaxgEmjRYYJJ6Vwf4lJSbyxYXZLCg6QomT/o8
0UMAOOtgxgHnEMimiBnvYT9SK5641PsoJ7v1t/gX6oMDr20yDs8Zt6jzfneWxhL5cD5UwU1tSkMy
lOSJ/xphTVTJ+fTIH/+YONTnyc87aow+GxuNPQzIEhQypakMc9ri17GqMcnNGJ2AbFVbMSVkVETv
8rWu3h/o3PhJQHv839GYoMTNISVZlRugPjU9b1ZzFFsCDLxnmAy0x5ahjJ0Jyh9yCtM6mHgUzRNM
lS4OoklFEJ9VKSYgNQG5juTVlbLGgWm9JOC9k8vF4UsxEe6kfcLM2C/YjNxRSIaovWnyWfE1FRmw
hSHHEYRYvL5j7oQCuFFmvPa8svgMFWU8++qI+tyJbfgXdhf6C6r5zrQ+cmhFvUzRFVE+DVhOkvPu
c/cosBhBhhyk5hYJDMXDIJk0+3lJW0wvYcpx6+r6j3NsLD85d87dHSUoSjG+kVMI6wrpbg8bPQvd
HcnqgH1fCaozXzsW5MUS2GPbvlnA3cAmtbuVbMUT5ofZxTzp9XUsgSGf4wlcd6rDhjKOHTUHo6RW
i+NuxqKBn5Mpf0799IAckquvm+5A/guo9SINdwATm/hg2Oi5ES/360Fs5QQwt2c3ZZhvx8X2OeGR
uMMMx2KDmCBBySoowRIFbPSm6ehubLnxz33VXA9K2BZ3D26cdMZK+8VoMARN8srElFGszL5FHcq1
9n0nt/dZIz76ITh+L9zMMI4qHUD0ONvmRIr+GcNJ83GBEubeKLJvRIVx+oRiZNyUFvYnRlKMrtYH
0USEehyOoGc/4UxOQEaIgTsZ+TNsCPm/0SeFyL6whj7tr11uoXVlXQVDrwVJyLzZoyMdcVc+RuIz
DlB2NTEK/qqrf0Q2iNe9mLomDHQ5q0dN4JFrmIv6qTvMMSEYCuKqk5AuKVuEHPQkb6qBnS8+DlpR
Qr75a0jE04vaprHbmurC7dJdt1xJlvjtzODoymLtiw9Z1NwZQwIv7FLgMJ2qeK+kRs1jbDC+zMQ2
8997e4o3WbwipjI2OsC095DBBJTE4AZUQodEug0XNjOYfO6VJb0dwQrfOgRocY1rtwlm6auFEfoZ
HssdOsg4NycTDBf2RrJ9biTC2DN7/aWzQE8r9kzP5Qb76mjhoHfJO9LIEhQ/FPyVNu1fXc4HvyVs
vtpCPEVpiu0/4esVzQVYTlxhYDvabmqMYeJPrpohSvsgqT37TOBOgNOui3PR109CKqCKnxGbeNl9
FZ2YBaLLMEfycOSK+B2yxujwwXMRQW7ZDVV7AaxwkARLN2OzZ10Bfs8sJ/y+hjSyUNcYQZS5lTFE
x/I0ksqAIvRgLYvhs7Ptgo5JzuvWahFD9NLKQP+h9z2fgn/F439hvFS1SQqefPhCPyCNOqHe8PT8
1AYHdC/kduG6ji9FKAEf+8ZkUht88z2V0fQ1NourgGPZw8Jwem67GpNDNDSJ6XdFAxzhi47m0mQJ
x/D/Hwhr5DFZ544stGtPFqvR8gkGnwYpuTsQSi4HA5ST4d7bYA8p623wCez6QaFnQGrtz8wFXRSv
21t+br7HCisZ95MvoKkwPwitI0a5uCXW3TLn2/YVgj7nwrFx7phWJBBur3IsJaAmGiI4+lukcjQo
fPX6W74Fw6qgD0DMZv6UApuDSVdSOERFw16rEtSGSDSfho7vLU3tlKCeWz67wuH+Lh93Fb2osfBi
XCLEFg54w/Qe4iko4U5hqxszbB8lMb6LYi/E1JR6csdydDi8y7X9bgYOayC3oHrsFWfa0pN0vNr6
K9sA74yVx8odpNTHZmAdXr8T4lB9LtX66I1eJ11SZA54lmDsW/6APnAiLEzFCoindffcFOl32LaK
T0c9YVtpLA3Te7Nw3OjUh5gNmqJtQK0hA7tFGCuaclhP2jq7OtMgvxlCu71xV5OSUDW4VaRky2Rg
wLFXqLaVDYTNGqxvw20uF9k2oXtdsIQi0dWFeG7pzBvSikIucEoLBuGlx5hiIsaWKXBiwGExOcT5
+AzhLzZCxj8QNph6eMW8FxQoFwWfID4hYZP5RqYSj8T8ZxBVu4VNtsdpnD1RiFrHcMfcQWF64J0c
zos3b9GakI7cRVo+JbIyIkBx3sTXGSG52783EOo8P7dB13/p7RHf8eqHnvzXu/Z4dWHevxqneOAe
5Cs9DqTqomwbnfsdZzbYp+otrR0NSpX3i2EYJoRLvW3BtgfGXtThUQ/jjANaqvl/shnX99UNxYnZ
Y2tW3bh35S9UTOepA/K5Le2CkOCggK05iZoEk2lZpc099a2mIsYn4Z/XaFobm+Mvb/lFPeExKGI5
rtPTh+eZ1UEUwQh2aop3iKOrPvpbSzebxbjcqQUIDlRSCDnAzTVTLUXO4usf6rC7zWRmILLwkMRr
224p7/bKRjWIsTrCHOWTJO0ys7z1KNp9QBzV8xkQYn07/kf0F1Ue1OLaZ3fZWf88B6it88bHTKw3
/6giWvlQ7DxpbVElUW82M4UgC0mkXcKt9wIqnE9YG/YsS8vI96bUQ5h62GqjTdfufVprSSeUPqBk
tdh/Xc4vkpYFD4ts/S4Pou23mNLwC0AWrkP3aIS8JMcUv0VFuJFBPY8tBXt+pOHwDhMVqMnxsulC
SaZDbRo2r1iT+OCy5fO1OlrkgL3r6zSW5It37v0xYzMQE/D7F5gaFSWoOEyqR/t0qvnfh2PxZoYo
HftrZwBksOHhTWmwrCwFJZIPT7b1XmoqaIRUEKyb4jLYefnkCPzzKhe3yKs/R/Ui68n7yXuwDE4U
d5tRiLB1VwKEemszbV4gSSkkZ75Ij0gRMN/Eu/aiPL5Fh2v3xY/1UlSD/MaCsoHnPLObtrnvIGnN
Jzj4H6bozf56wcXAG94e+RxJ/8Yk268OAIISgGM6FhXGNQYCBAOeIAzq8Nmcu0LdBxm2AYYUhCTa
1B/IPHCPIeIEQ6091EWgLHDg6grsjtzM/oiOdP172QAc06UskiAGsLsDMPkqDgY2TZHziBEKT8A8
9FGObaD8t6+iUcio9XeJxAhVP5KSt2OyjBteJ5C+F3YaaABtipZ2UBnZAmYPYhxhg4kLLdgfz/dh
V/HVr7moKXwrc/dcou1pbzbnOK9PIFNWUbWYrnC1LeUMx4HO1mYPc5mZKHvTz1x4FV/SZwe+4sPr
kVrQJAb+EOZFVdUSFuedR1JnyTqCpAk8cr5UqZlVI7bWUuk6qVIbJa6bETi0i81NNrj6YGLsuN4M
fax20vlxE71upFNH7eMkZs7GFwwrjA705VMRu5m5UZX8lwlfiXMDnPXX3t6qYANWoG6Y6vQSFKjf
9Uy2+5i9S0SKvHfOiRP/eQbqLUTRwozKJKtM6T0pthqvP9o805WHOA6mNR2ZnvAbNlGktw52nJb8
KCAvsWzoA1sZIsyNeiFNO4FmB66JJhMzpNK1oJ86kqO13k1WCVc1Hi4u7b7LN1RYq5nkw1Ng/FqT
HOGy0O8HdNg3gRKWLXocLc8qtmcNllQdKIiXgfCE7xoY/vUNSNMmGqB8d5shTjALgjdAIvDqTPdW
jDrlChzX6tFby4cWLx4zD3zp4ntYeRgAmtm23lxAuXv06yrVE0rGKwj8GEkUI8TGereW61oNyf7N
KYhkC4Qd8OZMoTtNSQ5AJKbKOmQMEr5IBq86fQKpzQyeScgsZv6p5YGOZ8ZXE/0iHgfMDwjdVgkw
8OqbGmFXWy+e5C/dT5EOi7NNEUuRwoZ4BztTkTKUyVoHoSMP0KlRVWpTYodOysmyke0YqlTTXDBx
gK+vqMkX3m8T3dxe2phk+Viyb9VsEifaPNsdQUWuu06B1pjKSyxB6MR6zbeUJRo5upbJoc8ltj8X
qhz0yH4L4ElCH81OakbBDHheVx4g8IzNrm51flQQmLjy/2Dmv6PEE3MtOIS0X8PycJEVn6WvACTB
3VRA3DxtGbxlUefnpjpQbX7ePLAbLCwXIOZ03SEB/CQAjLf0EwVAKo9GfDO9LT5U5meRRI6hh5eh
6YMTdccdXUWg9fxKaLwETehl21t/+9YevtK2d/ODWsYYqqGbtOdU4xeHpLQK4tL7SdQNs8b/wzRP
BTsgJkIi8ei8X3PDoPrXHtw7+SiZKnVYFukEk4NEFRN5DLmUKMI+ah8+6V5MpkZg0LPoKwsGIP7O
TTUSgE0FtaoVsiZ3Kza8Xm/yc7cV7aSusorlS/Qs/9XVE1dAc/sVbI3lXU4Mcu+Ek0xathZ8F2uL
XzlFJmtFUm8TL0itIhEPZdPQ9V/F9uYuMLsyhPFOZnFgl7zqdBuhWuLluyGnlnu1304Da0UhvIvJ
x3FHXg6sAv9Cvs5N2p3DB8Au0oOwAStWVfvxlGecwRZumCPV80fMxgGfSAzNjReR56jehyyBxIZl
W1RUmXmePFBQrsLCa0GEB6C6Y4UnWSHTx+3XrKzuw8od9lk1UqRh01tlQT5kMqjdzUK+vY5DpdYd
9WcLtvel7AEdjixZAem/OdWubAZD/Su5zkL3r9vUZYy+Ipiior43wga36kIWQvNqDipUbP/C1DrD
GALuo8HiIRi2QATeJqikVREj50c7kJGRVxbmJ/z4oVodY8+2f/VbpKOQxzycJMUGKKbOVnTPPDct
4TdL0HIgZNRxP6Nl/HaPqiSvN7aWP+Rt3jRS+Dgv4Xmk3crmJcz3hlBAO6mN27rBXAFNIgEm204w
sH2UsLIP3+T6l1mBTef5ZIW1mzRGV/DftL2ovU9DSLtV/jeF0mCUyAoqw4h58MZjpj50pN4IgoBM
ci1Njzf1gx37w7pNvXTvSXHaDPVOVxQpVy0U6aJwiP95Z9C/riR3wD12v9YTLQ51Cy90P2406vzS
lMQy842oI/0+UtD2Wqr6kJPsNXHPYmbV4lvz1MuBTpWkVvjMNVoiYhxf5W4oJG0rAv0j7+hu7HJ+
uNPYa1cB/VHwkj9cJgTJm2H3aL6PuLaQK4qpRIZc9km7Eh/D9fPvaNeABuAB9onM1Vd501r60O2V
pr1pl98oQhAZaiNcmken5iNMznBpDEbEyqwDFvmAkeXfTjkFUN64RFRbTFXfGr6s5V6VeglCLDZr
YYvPyK/EHPP4I426AV5JZicPUgQnccawNO4Wu/XxOnaT5EmVFgTMBpLOHFYEPhO+ml+qvegnrYrf
EauEbQpJrNd1GBTK/3g5/a2dX1Wd4sGfZ+OEl4QdRwKi153RetBg37zqagnuV5gO+fYZxBgftlCb
LGDVAji+lt/17VB7235k/4jKItzWz3Cresftc+6wfjj1N17IHFtCmUhp4RjNx9QDVbD28VEclyJi
STss3qFQf/nz5wa65SWKO2ql95yZaemVIXQBktLrN4xM6CAIgZeQ74KxaSsFwhyoy50/E/mPw0iQ
BHFnyZwq9weZyeNNqw3kjE0Q/tDfTPhSIVw3Zyn1iXiehrJC0xIU2lDkMzezTcCuPCXKSEhf4Vqj
5gqQnlsNxGLrznvlViWcxhmr8aJF6Ump5pwGE2xLzwRgXPQM4RSDB3NMpyS4CeNpH1PYOuZXaxOM
K7QBvYJ7Y1/o/Sq25BuXvhvHZy7Eer9U6JyRbIq2goLZ5J2NFo2hmZdPQVxwn3AolcRksrjFYRC2
3BlhlofZi5azyBuUUzQ8Rcx5nsrslnhEFYNeMq4/94IaeCf28yuiLXFcnxFcUEeUm+toxiNG5moW
GET1de/AawMzx7a3HYJ4wh/Orj6gNzQ8EsbuKRtb4ToidxuC2MGjsXHNfqK8ed++Sx7AZylBjbT5
xfZiWRAqZRPgq0uJ3Im+nKDoNJhBC6ZqS9GVwSiwBKRlkfD/cudFnPe7usrysupGMlN9ZQisMs7u
KNDQfsewsoN5QvC1FC18esRKfPU0QfvOLyp4/kk0O4ay0Nxyb6oloXUJVVA7KKQ13AZfIRLBdjFG
61BIpK2VDI8tNE4IbGlvlIjscG6JSYaQkkVQsxD9XdrXHCo4kxrYVkTMF2kQwQYiwrs70JLwWtSS
KUU6r8MH8wMijGaAOBi6W65zqy5ygDmfGy16xFmmqiO0FvaUovLCgri9PnB90pv37a++apeiuvuo
fdy1xKi9YdzP6Olm+z3X7M92yAqBMvr28omcm9mOcKyBi/L2tp5Xt91sn0e51D/dbPmHjaySprH7
rCdw2Gkvo1jH/WsrVCJJD3IxzWpW7PkYHcfTFjPOaJsNPs3ZoiV3rhhVkIGjNEOA4EVTgw6IDBwJ
3sqEVQIJf79umcbTmedPmK5+qfEP/3HsIOL1uAlM1kKHmKlBaYs33eSmm6B3kznHPj9MQh7vVcla
Md+T7Gny9w2G7oIJSZsfjl6rwWr7B3fAYmNEDN8JFLkaqVytBvi5h0bBP4cXH9gOdAHbwDXkyZ4u
9IQ0nfBy0kU1h8t6z2OrfF2ZZfaEppgeHkaj7+J5721iCUgjlXgqv0TLy3M8gHt346w0iWRXlT1i
QC5mvwJn0mIjZd43eXLHNhlrU6bEu5UaJ1k6PQT5rG8V71aOraxOJOkmT0B8Evq7Aj6K+GbsPPl9
niwjTaUz9HLcMdJCnqlblJ3CPysWpOGxpyaQd4SkXj99gg6eLCyKZyK/u+OP7BGWJHAiH1DCWGzr
RA2SQ0lN7C3tPJ6fARR28FvABBb1kbNB7xPqwfY86IjHEvLq8tp2dLc/YK5q37Jv+ggrIVrhqz/E
7BNic5VF5Th60CYqxONC08F99ZtvD4zZhyL/y7nLp81FkY2bTbFhofeTbPVlAp8TWkSRMWdhNaih
MihSv+aS5vz+B6+HPAVLfGd5GBCKLj6IObBMxOYoqHpa/66pIiVcIcHxXIDdPlUptV1Dx103sXkd
16Jarz3BYOmxrAaEpuqbO4po/vKhHbvdxNGTWqWsjL8VIgVZSw7m0RJRbh+MJAThJ2db++uR9c3V
G8nlsL4c8/KLqHHIPyi0wGy4RC60PuvPeG96+O1w6GC2DSqLxr0lQiC/iLCiDmo91RQkz8ve/Xzx
oO2xpMkGiAhf5GI+1Uf3tGaQjQFnHFid0oSrruGEHMw3SmTJscuYhOe7oX+P28ngMzQeFdntwJ7e
eWT0IWARcKIJq3DZx/GtOSWTRX9kLyB+Gw5PPCMGJHYE3ffT81VgIC6KTtpOCZbq2368d7qu7ShC
7i4zY2gnEgXyqwDnhtS7TZwL68XI7r7xHsaj4ihw0plNTUPeIFKJJkk5hNhfC/NLm/e7jCPWEFij
gPyIsP7/1zBAdJZnS4FJZLZK/Qx8JBJy/5ImacwDXBOvSQxCEyIRuQT4qDAPhYCXQcSq+nMjTrPQ
tXhi+xleVWqCjly/z2HNRJcLpFjyeQ4x31ZTBHe9kbqGyENPYOXekqCXrQTJ5aQ+Yh6BpniqZbxw
zkY8lgp3xfAPQUUUZbpU4X9Wgt2dtYDaOZ+d9099XHPep9f7OqGKWwgwTqkiS7ghoytLNVrd4zhh
D4ZM5jYhSN6+mrol0SOOZ6xTlm1/E9DeVJHrbD0rqBJmoHYqtcIfM9a6HnrHtP0KafI5/W7OpUN3
fyI1CRyg4fHOIIPBzYCNJ/HbkFR2q/U8Op3h+k3d9eH+f36Zpy3weeLg+7trn3frbWQelf/Sxh7i
iJs+QEd+2XxJ8XPCk7DQUzaVWwmZy9x/fDM38O8eVbgjDpXVnkwP+syapzO0Hbhs12FioZbWsI23
HuVsnhvYKDT56Xcf9tnw793HPDluaKIG1BpFTIOVwlUt7RclJtDLLXACaLQYQpUOLWZwxeaauDq+
bQLOge/tl9Yud7dg8V41Nz1Y2MNIVC9C2oy0tNYApXCrk9n1ms2LOhFKn04BxF4vSW+CR4LSWkeS
UUlkeDPSysUQVvVKWS9QX3wPmTLyn2bjoc0nKhzOJwoNB2csnJZHG6d+4By3mDxUjXDs5JxlqH7b
9zPduGDZxslinF7H5GZnQ0C1CLyujKjTtz8R/S/sj2A/POqZWqiVBEmD8Go67JKV7LpPvN0hlJts
KXhYFvkYncPtghIgCZQfcMV+Qp7DBSUpvNiI7dICw6ME98rmrVWJ+ezKbTuvjYeyjR5T09PoPfbK
kSd2BWMkEf4kj/zTIpBFG14TgsO6GdnMx93ch7L79gXNH9P5HpIgPS0Edl/iHc4h4/u7/BAphAIK
EzoFsddWD+gmseAwYJBQhM4ynLQAPO7d3UNcRoQFUc2FdC3IGOOnGpCQJXc7IzXVwIcvwmYnSdJa
rFgJaUipHGUZixfLc3rw08uXi6d3JraUUrIFvmUacz41WZS8KYDUpUjKxq7lL5wLkrSJvHUfemaj
OWSY7nt6u0FoNdZejWxHr5kzpG/mbbkvMnyK5oYl/ZcrVEFbPDQRMadh1lM9a7rTaqOK4Ffis9S+
lxt1CXYOCVTyHzHw3NTu9ja5K0zP+8c7gYgBgjV09nXGsv7lPhOsD9ktzd0JHN7eJrDWbOVoVEte
VpB9x0OW5YIeQgYtXr5VZn3ND5LIKh8SPG4m60xw6Ubtq2AYXge8xeuSFlFU8G8zoPnGfksAxJiO
h4C8FFqp5NoQZEUwzCwrwgFmzid7q+DGTb0RBBeoOsirhxPVfkE2vYHCrevCBtHTtQika1uE/tkw
Jf6wku6pOmfhDFxsEpRFqNlCOClmHGgSSxXQ896ltEN+QK6FhVft07pQIhKonbnN5BIEHoT4QOy9
DNeLvjMkRINbblHOTTW5UT0zowx3cFlkd34RVOO51h0QAGFUtKHq/0cnGzMLv/soP6hriwIhrfvH
r2TlDOzFlJDcvTj6DtpqsI5RM3dziS++r2QQAZncpNEE7fhZawKQjeS8CuEM1s9LAOcfuY8I5HsK
ZG/sgWvmEZS8Fu7c0m68Wlmwlnn6hxXnqhAm3gY2gJRq8+2UukEzKPn74Fo4p+Yo+X4hfHlZP+0d
7nsfSEQw8CIHG9QltobL4Lm1uiRNzXfQ4gw75EoqjYRGXbA3yHQVk4YXpHeYyOGltlpYf2nB9Jp0
VuO10qDmvCqCNPPa7sSKcGSV9+HHMPkT4Tl9v4VOvfVAgR9LJR5qdz37Za6NlRTssjA1DPYnAi6E
zgjXlM7BgqAGR2mqOrKP75AjGi3vuymS9vUzph6v6YznlV97J1JDFCHBe5lpnG0g5QP5yoZRRbgC
Y5YGapQGhf/tG2MYTpBVYEvE34E+xqniBQV/M6urnVX5Wev7LEAR/GjG/OOc418y0Izz4hXTOx48
mBodx+g3hEdMC1Oied7BYHLnRJB1sAMrS+o6ZlKvteGieHjS4zuFKQHsiEuv+3R+xRwuacH6Qpso
Vo6JooAmpOzRYfu+iEpNCdE3txPI5Yf+iZRk1EGj6pf/vgwIxfneJHwpgdOTVGOWcdX01QB4mGDw
+LhNYKVE9/9vSVLaaUoZ1V8cq6VqOJpBmFt4WFuVjJFO33J6v5s7uygOKosb1X1bZXqS4tbd4a8G
XB6IgGR/4qiGNsB+GncuXkLi61v/tun+4fZjbfPfqeJ+u4OaNdwrRoAFngNSVyACKTz9wqhwJdbT
/3XhfUgp+I5A+drzoG8CQAi9JyOS1PLK/3ywj6RjVDdP0WCXWBKTQzKE1mya8+1wjRqiF7KA/fMr
w3HqmeAk4hADzZxTY5o7fmTZfomGjxFEQcSW9usIQDa3832shL3CPdwES6htR8bKewMWMUnc8QO/
kwRtfouo8BRBK6EzlJAIB0z71QLRrvh8KTEw+D+0i6s4Dqt2y2ADyEFnFaI6TM3kyU5XbRGK1e2x
xgYTPQLO6g73Mq2A7mm2rWMlXNsyDFIuJR/bjPPGaXEOvLdjH1lrbQaDUPJDdhfQpDfHU6Cvw/y5
Y2APGDD++bZcC0/ZevP9uFMa0CYS0nP9ORS2Dpwot7OJHLgDYGtVrevLh3tUBqi6I+JpcHK6FlCF
raS8WuOyCtQlYmkLE7bbxmQzp2qLcH8QTOQPoSf/iOJCvO8SaodjjJjagEFEuaLybabKUqA9Heo8
8gMhKKY5GC1wv8+BpJ76f+4fcz9RSJlZ+Otlr0uLzmXnTt3LxHrIhOfegLKuf3BYZ0gzCN9s795F
eraHIodQTJuwBt9bpXQulDLIIvkL9cf+6dEqLKyImPNFC4m2F9jEMSNDsj/lv/3lDOPRcsI5sfNZ
2Jq91543iUITQNPgTzlEIXcQyA47tPek20BrROtxBbYnpZhpYkyWI2em+bMgOkHhVSuKAud3Q6uw
l9nk1Xf0LYPo2sSxpsC68qPwdqTuRMOmOkoTxoXeja2AgaeK7PTumTxV7rKOwvaa0IEi7YX8Wtqu
a+vBAa9byppyfUDK8+tZxohSwkSJmeuI+YTNRLbnfvxCl+aRWsLDantarF962w53sqVxR/aP5LIG
2jPq+tf+3FoNe0GYQOsuhoPE4chQVWOoUDkbDCeLuoFO0UIYvQfd8c8Uwg9qe5r+p77QphM9XyC/
SzZAnLm+q3NuKbtoQssl9AUOUOhTG9n1ao46R36LXbkhbPknT//8HAUamOwa6nuWc54KPuOAN7ta
1ICmEkzKGeRLgSF1MdZyXNVaxu3cVVGfqunLDcBaLQrdYVXYeSBkRgeesm6LWZqacVMvIH7nmKRl
ZMb7qq+9ewAoR7KvFt1JtF4K1/ZynAub4hlZrGHunXUWipR+DB2CVB+mh6UzdKNlxaxDOCVN1CpZ
LBsY8wgQPql7QjeV0R6i26No0X4FsS7zUzrSsd9Ozw0saFFS5lQLC5dpwrU75xGh2NSoo6jtnbFu
xjvLRTaTq4X1+z1P/6QG0JKw/DNokrhWIJTgh+KzJUoankhvaMis1IQaM+VDQksoCAmOaQMnBF4M
nI3xNr0UiXVZ2bzmV5q2yorer6wZ4U/Viy3NKaSzL/Z/0Ul5J3jptWthirZAGyJgzrkj7TbHu11a
KkdLnyTzJ5EkXrrVZqGtB0Qow6BzzmeJlYcU2kAmgQq7BdMKr6eEwwTDTS8M2EiMfA0SpXJ0uTim
TQqjXuwnMIMfKyhKL3MgqxBqVEtqCAvMdTrW/t2GhLOi5hAaMNhnwGtY8vIbn8xxlzl6VLRjdh/a
VuIOc7zHIuuujXLyCu2rZoraO6BQbD52X65SiwwZsf0N4nzJIKAzaq4yx1Ga3NZlnw82hxAcH3T1
JxhJg9OLXmETyw+Nh7D65Ab3YTlfulktYqB408zwdEjDwnOUWksTyXmzwilZmbf2vFoV0KdsPdKH
UkwbR0wMTMpLf2plgO/CZvUgFBX84n3e7nPLXjpMDq2ROCvnkjV0jlhzhvQKQ3RsSohRgAoS3Uft
kCCoRq2D2SBcrDI4kXy4PvIzIYzGoO41enEQS1ZwN4GtipeBSVdB8IKnA21SVPYDAuyZ0+7n7dnn
kjaw9fAYM/lZ3IY2E9GsqEoB14278d+ecN1/lQXcDDRuoZ/zsqtH0VWrMQeuc+t2xdCR2QY2/xHm
iLOESbXn8CwPs+V/O3AjD+CoKuJN1QjZnQUrqNZlYUEeWH5DQH6zdynZLTWuBvEH3gFSbvqO4LF8
ELHkw65FDH9YwpOn7RPCeiqYPaQhaPDkjHptldK7FPjDfm1xQlC8nIDL7bumdoRWDC8BECuX4GQi
4eJaSemleTVRY+nsvM8sZaSNn0sHI/OsAtmMmRktZ3OZC8gAQVQmUwsJJQ2trEOUGObWGQiZ0ulo
13inDDCkbIGSZZi9rFICqDf/J77PYMQOtzpZsbGo8N741FnYEuYi5IXMmoajyJSe6b1LrR0AzFs9
ukd0nYnJfYRYqRbQvI04yaBE9Up+9BnLeCwqydJpWcE+MdtDlcfn8ChsZywMy49AbReeJLnFYk48
Izg8yIl6kOWqdOwf7AHpa5ywIUsTySMQWCFM4x+BZmsdCDSZr4hptFuD3fKHAEKQpJeC1Qc867WI
DmqF2m3d/3Aqzk0zP7hZhvK5tOKM8XceONCHWsFLkiRUOE3RTCLLPAD+lsBwF/1T7AS64dKBopvZ
S9/0ws9xYbwaeMECkKaDnPdUQsAcRjEJ/mgOGc6hzE5xrPvYuk67g4Fh2sWUApHmIAx0AeZgZxv5
9gjvX4KZWOT/qAXDPH2U7Jj/WkytKH3zLStcBnG/qjYVdbsApTBJNkHZMVLeG91IFWGV/AONExQo
TOrXn6k35IKMlI8rnFVxnRUv6WWcAojT45K8u9PYmBA79MebR4ngBts6Vua3kN88ABKApq5Dv7/L
6Oi0hCb8zm4JvkWQYCOnnwCsD48sCtUBheoV2RFfg4kK2UdHZ10R53wX6NDfuJuPv3oCvV0cpp47
w2Zdu9EObh2wwsCBduX4i4SQ/6xRLg9GFgGvSbK6PSrpYNpwnany/YYEhNOHQtNIuUQghZuv2Fo+
B9WiF7VmTbASp7zKi+dXkvgqqxSjvvfImYaJsCyXZzPO9d3CWyC6/WQ3sbIvIRf/t78UBbQ2KUt/
QARp3rL99uGEbKRDP8gTeQPNPLIRUNmpWBfEkWlNPv+q5KmlEDImyJR8mxU2bEaN+cye5RuftOzu
9iIfVDLeyudnWavKaR4TkpgTHrkztE6oSCjHw1nWh4z06LWbczYpoXGjGfSLdsWRvNZeRlE/DSI0
1vzk2SjuyG1nZieUICUyBiYFmxARQQQEz89hFlN8WBuxuWJCP2Xkh3H+W73WxZwWY29GOZmsLf3v
rl61MFQgGR96noveFkFuVBURuD4R/KLgluADKQ4933/ZrwX21NwQaxu0oN6swt/v2awg52fvqC17
2KOxdwzuky5A2jcQDrwTUef6BcqPU9mlE/PFo3jTrrzCcAGGXd8rowK5Ezs7xONsGQ31cc/aq7Ir
lyPaHrBOg6AnQp0smh7xFuIzu+H7RUlDpyWqkPq53etG5JjGFWeTJ6BvkPddpHIiFd12LWEv35II
/wdADlsiJeaEP5kcrDR3wD4b13zUwQ1CK37403BjUzsXa75XyFBrW8SCGFA7JNwakfo5KrTz4ySg
CV8obcMNg4PdArjKl+fLV9YkhKKRf90zgwJbLQybcVS+ItKu8g3lfYfix4hdCFxT4s1u9iCDhIMs
wxGoeYTM1PuQ5xSPyro/5YM37hQdaEXXeHY8OqEwLw1d/B//Xgn+ELEilSP+0XWM+j23lQgx5LjD
3OsDxTyJ0p6hAgdfjYSHa4O+IoANbDeEQWpB4ctFxE5sDLpO8V6FunU0NA9ZovryMrnO/0u03he/
SJTo8ZUcenQOell0Wb8M3BOgMULs+JJoApRjEJe7Ag8E9UfWthsEqHkw4nETSWcTDT5aAdnrkH9f
liuXi++spFRuRSqjUGzNr6oJxYlyIpnhz4s6w7y1ThNx5PDCP8JDaAphqy2R+rQoDM5rEaBtsoni
W5ssG2IfyrysfB5vqS5z2a2b02q9+Xwo3fmoWa09/C9S1EMbwdu3bITsBbRKKErw7hAVImZZ7EvM
Kq1YcC7MRKTnigfe+gFhCPnqUEWYo23Jj4CXi+JxHPi1KJ1BvcTm/BHZ0ECmBRYDZn+bZbSAgYX7
kEGEpdpQ8c8znUrL2JA8epsYDvlkJaZNGLxHmZ/LlFux+6ys10V+/4F+lW9RK8VXiRWNBnUYBDIP
77ZpPScxfH5THa/y/k5Y/YCysi+aILzWZxGpD9CiSVtXocgfzJCNPt+RIFuI2SntG5Vwi6SyNp8l
HN83L4CIQhWhKEJnbbaxUPJoGQABavRHnjkJHMKScI12VFyGmJkQAF50UycekvYfQJkww6jm4bw8
xmZwoHypPW5oD+KE+o4wEU2Z6S1w17CdQig0z/xs4gdBlGq7+9Ed7cYqOEBiaNzvHamEPRWOjOUL
8/VrUCAIDgu1XqD8e4He02FHIpuK7vsbW6r87nT3qr3R4lpcdyc2mIlYDVcJn/vyxN3QUX7YOUzT
1iEpZvzWyIPCeIwmab10jm2aU2tX7YDWn346iM5oZfaCEy2pvqxwS+BWv5AUxGdNAvwG2son3PoD
BcaG8eqP/1Gq6V1wcGBIMJtiDgumuoEQb8ea1Kw6/PVRQ8y2y1qf6mH8k24jfuppBmWdo6XBBZ5n
mZhK1fabflGYNgP1mmQF+CmTwdf8BdIDh37XWJWb8IB0U5sPgBlZd8jyXavjcLeq7uA+CtPAyhWW
taZ2EjXRxwCRASjmD7uA47lq0lraS9658ExxJfdmU77kjaso8ONPmUSxmS/RFixJT5x5+nXMAyKB
cv6kIfOue08naF9InVBmHOLY2XtYG9fhmN1/mduuUs41Eka9//BZSnfA6nuevZnmd58JDPkuz7dG
aEFKdnpWP7M0Cm5ftXcpp5O6Lj3+KcYB0pHqJ9y2iEU9MngqPpUSJ3p4eHZTfM9GWMtKHisykzcy
7NgR2KVTckFJ2Hr+M4MRXjE49tNXDjJI0bi3sc9ElBVahRjXmA6uP2I4/ZvJ76BfBH7OvgWiM87P
4E0KK3qPnpco4RxZir7lGDeVmP8k31WQerDy8qpFwscI6n5seZPdKi6MdXMenjXZHO8XBdHQ16y4
RVqZWNzdKQX8DE0K7Dqo6tEls7obqKHYMDnIR3B/hVJBkUkz6aaJQjHEoorr7xVr5Wv1QIir2Tnh
IhHX3u30iuSbmLMlfis7v6b3uZFg7/nvlDIyoci1AZKZmayzMN0r2MYjuooRAOFwpQI41abH6VHM
o9CEKbWZvKrQkN7bD29aGsM8gDzOfsELdCJG/uvAEF7U6caUtBRkTSGKnkNq8rs+YvkAcr3SLbG3
Z9KDg9rAyPIpJOUQdG/rvi3uYI/bCezNxoRy/QUP/3ggu1u1WB1+ahaS+WamN9CTyubirI1BK8d+
YEf452FF+89ntUq4QQCFJcm52+5arpWj/QYAREYofZq6FKq+uZE9KxczFnbPPK/QwMDLf4hv9rmB
EkePKH80YBSUQgZpZoHnI+Zsu/Y6feQwAAtlZlZCdE4PC6KI51qdsKvR9LcZUmtMcEW0yA+eR4MF
Nd/bcYMZVN4NODgdqOVC4JQ4KVAHMRQHuz9YBdrkyb2eb+2KdmfYoZc+tvu7AnWC1S+ID/Qv+k4W
qiBscNAS0EC4yWtqywM8rgcQhC72p/sh+q02vPF47OtWHfCi8RlyBXGARKY/lWNFv9PD6VwfMPv4
BNWP2kxXtAEyl1bNp0x/oI5pup97O7gF3nL92sAbAmxlyk0S5JCjnOjo7GTpP9fUMDx/GpF3VcHc
2IuJZLkmqll7taQANZ1JmOnTSAXqNSdYiRKnonFLD6V8as7Bla/4xImxkI32VhbybPczEU8eUt1A
HxmU2lbPlqkADTtK1SA9Oj4cXJQzJy3jl2sSnyVgNthekNV1YhJTLp/AgSIZVDpLaS2BJsv/WWWV
ha8/sHaNJhJYgKucf6tU2hvHxe1KWvCWhoclrPuKhfIOX53/8wHLqB7TvUQ3eTXx+kZIyRrcwvKo
/1nI+yDGEkfWcZTJwJG+cxWtiwH/jnxhNOls05AMcYkfRblmQ8u3HFWqeDMXBBv8xX35Hm9MlMIE
fl/zD2sDwxODnh+IOnQvwyvqrTBMWg+TH0qZ3fGhkAHB8Fopfnx99t8uxgmSYiT6corSQ59LOqJv
92190SeGzJAwXuX6LnV46x/c61EHdSxwu9GaGAajg0wZanNfeMXbDOpHPCHIpUStuNI0GQa4fGTR
+m/9k1yDPJArUSzdiGV54AilVlmoNPWPGli1z9P4uHoiDo4aEtgberjTQMpKsnTpioG73idqlCyb
JorXQaxVtGIE/nRBm4xGXibYQFRMe7cwnPgKZ/Y62Jvvj4U7BpCMBINKhDBwtJbSlB9UixMJSOiH
IpYVxh9CWlYqGyhUE/7h2lcS+nYNMUqBm4SS8WGg0UFPoeBzb1MLwjdScUEK1/yhjpO/rUxM3JW7
niWp9U66BdmajXyRTdjahnSbv6iR48vziEMTRk2pg9TBQ9c3fHZ2kxk4fWf8aAybm/P7gCeH1a+Q
dd7SWSZY7DukHXBDtegLoW8bqliIMHzf/78kyCGpvfRexGEBmWW32DhGB10Hn7Wqg2etMzbUY8vL
GFg6CJWXYMCRNDhEYAK9l+SbSq3zY48GLuPt8fR4z0oZWv40rZPJ1aqfkLUMlXkf8/vBme76z25p
90pybQc+Ogzm0kxg0LLoq5BH9t3k6c29XES2jueJTqDN784wqWTIejxEC4tvcWN2O49OFuzb7gZW
SPl6fYyMZXTtspK8/L16LT2TJBldLdocdhBgqhLhLakrS9a8toM+DDHdeEZMVLnVFpqwPkIVSyyI
ne5+8WGMXQ156MpSURfHL4fQLgnfYcolrWm1s3LS4+/jhCInUqxLk94O9rqM8VX0n5B/+JXhHi+6
LHv9t3c1DJBfOVTLAkyzzhd7l6tb8hKJMcj6SmI+DKb/zNZ/G8wBYkv4VwSuehgYbgToZtwJFcUF
fkPqIJZIqmaGLiC5YN7Z9Q0AJWDPGNvhUVQuO4LRcqzfz5lBPyq0Tm3W1DaXMVTBktx6ghxkmi5c
ZbsGu/dXs05eQVESEI+0y5kW4qpNlqSvx4M00GNu8D2WYR8DWEED35x/MJDIYpkhv/bWY6YmMdQr
vaCzspkVKjMP2V9j418quh7QiZ9+R8KKrWvKaf/u7ZdJW04M6jK8rwFvLhxztXGFuGTxHihGyiFl
LlYuVQvN85el/EMb4x8cc00XVlHYaV1/FoVr94TpVMGplkliQk0KHYY8UKvm/oDNGyYNF0dbCaf+
0yuiam5bV6xvhJHDmbJ/jR8rI7VYlEhF8BIeGaFfcqcVuW/UGwRdqs8+tNb9d3DFMed+WrDMuW3s
rzhuv2DVMwXv5zjpdz3H3/72RfzmMCmQ+4DyOJdxzofPmrDU+E7rQKv87JZUtrIQu8owJoFirZPw
IBusCA3cJcwdYWkxh4LjO7b1KKb5L+OiQZHDj1W5yZNupF9riuFPPoqVrg7iYLHEz/4f2k1k1EHs
YUoiwNeMejTdxsja+ZflS7tq16zezQH4xGjOdoP2vberRkTUgjNC9Tnkulp1lUECf25Fx5CI/gr/
vFgbx5OH9Cn94iGCl/VnXGqGVlsuBFe6P300lFi6RnfGtB/tjPeP0dDutUgaKV/0CMVGE3ph4Jdk
SWAvWQ0ObSMUlWmmSsVrssJ/4eDtw0i7KZTsAqglJQZUT+VsSQkdxF0dnGzdYzPbX5Up9ulpn4jr
tf0i68lhnpa/vIFq2a8trP/HXUEbM3+Udejjax38B1UmVHkveUtq+72u6Wm0AX316hmHE1HgpQ+Q
1dBx8Z2mnC5l9NCN8Z7wp4HyCWKWvjCXKrOPWxwSnQavn+P7eSzDR65SqMm1vDBuYEIJdxeRG8ke
mCzgeAKQBYREFznst9AlEQH0V33iI+atFX7OOmL0wXtz8nHT8VIzkEwIiFOVsFa/sIFPow8dsCZ8
wlpqolkAZxRXEF8/m7PacCzCS+pMKn8bXRJhD9QzOVLNGc+baVP1wwguNi9l5hV+QmMw8k+PRSFv
6I3giPrJtfMZMrOJnoCr5M5UaLXGgcIvRxTsPXQvlKLjpNKy5b1ZaDjpA7NaTEK8542cRgqHnvtN
bfApoKWC870drZKkk0H/bO07zDDjzXmNpqu8uVXyyf2jFJL69Jl9p7w9nbGEesxGIcLx/fjThssv
a7dMmDOflSkbmVlQBS+EUUi6UNtEICd7590KynhZde1W4josTT3r6UUwrUOjtz54B2hUeQTWPNjZ
ma2FFrVjEAaAvL+W0QU8Hg2rdmEFcZmXrqpUWPsrlA8mp3XAIQPJGfnk58S7uCYQeaJFAR1yiKnz
tIxc/5lgF/zlnIztQj+nlfq4+dpzjcL0WG3npDyis9v202UvXY1xREEwFuqj8+qnn53ETjqHoffT
wfehe5aznpGhDxHxTQ6os9l1pqlPLr25bDowsMUKsiMQxoUYJC/hCoj0zX2SPfHERhXXOZGN7E45
bH/ey+T4n0AYeLtYncbtLj8G47zrDbg4nlcs5G4ZQLb978rHrQWqgnPHz6GCxYDTlHYM0dXDORRU
bvOSwea+8ftBftZ4LqI67y4o4Q/X7rMWbtWerlbLx03o/OKi267q1BLvfGGrgPWy3xmuLm38C3My
f5TS0oAhJMvEz61lsRGn31LwYxEtEKjziTCxcV6mJOjyi/5gYbZQjwnKIKz0mZEooCOCJs+58OMe
7wo6e9TsI4jS+acwmum39P0liJtP+K26JwSagLwYmXjXAiYxnxvKVHq/3cQMA/htO0XfhgxU9Uj9
yWqwcZvVXd54z/sJR/0nC5ndUjddClu8ND1vPHo2eyeH3W3DneHymQ+pjUwys5t+gBqpkx2tTQhM
ItVj1tDBt9VTaxozcJeBZAy64ub3cz2BleuMuMVTPxh83uwKORoGfZWUYo04GohGF2kol+ZfNN8h
mhjMntNBWTt3jx0dJXcgiIkikxLDv2dVQNJiiKzVQdieNcOUqz0IcGevrYV6a3ufEjBh1EupDpfJ
gJYmp1Kl41rJaD/vU+VJ34wDIxj3tGYxuV/VKdZXD5L9dqFy5FTGDhtvuNZdVIjl8wrmhmEP+Ahj
ufcQ7gp45Yope/t4OPMSdDfoeH+qbuNqe4dWa+9P3s9LjZfUQkhKvSH9a3uzJ7BHNqVZ+Yfn3bQE
KEM7bI4bloGqbbc5aW8EH97KVlAuP5EGh1II5wK/HxMNZl8zWFz+vYg+//5XlTDybHlm+4/g+TsB
tk7xgSiHLChoSmNs8zgBiXUOti0FTDeSTGwmXbNvhmsnbS0Um9WNRakNTkJHL7kAkKFknYjVxKOI
/QZNC+mzfq1iQPqcqHDl2NrBHP0a++Vehj3uOQNti/tiiTdw0YKDw0GXRaYg7p6ad9ZNP4LcLOCd
3/tK0i6/6iru/W07PU2HJFv4wMXB9Yt0CcmZL+Z4wSSbd9dSEAThdTfoqD8crhyzP3xoxisFav9Y
Apab2wYqHdebGbqFIfIt7IDkNhkNdXqFuM0wM8irwiESX6yojDVFXrk2Vfvva/3JwDoJKkuOWo/H
zH8Ga83nT0UxIYdlgw805pv3HSWfGWVHWffInizivrLPRZBj/BXtZErfd4ZcbAV/h7lecO1vzXDk
mbP1E5CAWXism3BScUw6bDeHDOdFQq9GBPParY8HCIn+EmHdCFpvkkKAF8Pcs8rvn8FZDQMor/Ek
uvsM2GkAH32Dv1SwLXZxQ8apprGpAyBFpNKRDgseoUVGUc+QQwK+kve4NB1SPhFpxvzToSvHDk5y
j5DbJDKByRD8VYUm78dOAs2VmBPHczLJvgytr7F46m7/LsTFys5h/007KBmNvjkT2Vbiwi3q75Xz
ALuszfUcoA996B0a6+ArAFjRMhjkzilZ8wwdOG72YY2Y1C6LSLb6NPF2m44KaLsVKaStVkONF7vy
NtXGohek7u93EoPmhZSQ7matxjkt4sfSosk9dZeEmE0RQCGqKBqStng3IFjgSVXXkDtAC2v7LYeA
1L7t02fAX2qOeNUyN5DyGkTfHgPtpYXGnU6WDMg2wcN2tF4bEwQbaRv0r7jGxBuGP7NJ3u7MwdNm
22g58yszaFgJjX1TbQyndi4cWdwrU2BT3Sg4n1+TteMqatyarqlvd37g37vYPbAV2bVXozoSaIhE
c3J1ARGNnE5HaSVq1olxdnn9XRX6kYhBhtB2BL6sGMf++4eaD/54vCcTWFryOaPv0ok9n+OYbR2i
S87VngNWQEDCajmGHJXWLNAfLyRlPLaqcXT8Aifa1zSjS5/MbVtP1EsOKFF54Mo4PKc2YILncUqr
fUh0rnX8IGwB6M22XvRw59Nm1W24FjV6LUOiCgS/z8OHkWAOkxSdyG4QTcVgQhDNpzt75mnvzBr5
wcatpp5DRjNInmgcQBI8YG+F/hSoKF6cVqK5sF1Hme4FcOKRFbhlaDF1EVwYNHSQbE5hs7Mv/Fox
cb/GM1BlAE6YzgF0E9jyXeF2Z8NkRl0A1glv1IbyuwM3vcTNQocP72pkM7sTjYWYUmL01UqW0NNT
dfJrUvx9SQn6wZooQ3AcEdWKbo9DwdJmc55n4IPjFAOMvfyN0L8Z86jw9iqnNmzHfg/iGVW9703d
A7h+fY1eHqGGvVrlbD7eAL0TC0m8ppcA2rem55xCBdJCLTFZYih1jqG8/1fn/FKHUQJjhcTBEAMQ
9Gi2grocKHBDeNJvuXzcH5auPhbZrwumeujocGrV0AzbBuvZywaU2PF9SUcJ7qXxSNQqyzdk9LXJ
Fu35RGrl8fwCRL7VdlzhJ13v6BKAsIby8oZMB4Z0pPjLrGRbqN4Z+zBBzHx9r4F/RoPtlIP5UIH2
XRlhEEprtREgMSUShq3JVo8ETesGbe2+OpQsR4NnDkcxMzlJ5U6l8iiqfAwxIHI/eb8cTCdYZQ1X
J83nJOKattqUv+XFu/S8nxNQRJNiHorzE2dWWWc7K7yrF46MPQvlZBZzs3IpeRC6ANicFN3xcjSW
BUnEjeqKYXqV0wXboB2xpLIlzfUrdwKL0fbHyCQOxclI+d1zlPxdhM1grhJH3KzJ8F3/k0Efz1jN
DmANTjcZcVkk3wWuxYTgkSZT/L70Fn2xWY3sF/cZ7hI8LK21XV7igi6COlmPVKWxMnbuK4dRo28Z
6/litRVdymjrFQ8MDBipx+nTzWb6yPfQUDlfMZEaRGxBs/PMsgDuo1emAwv+J9z/F8XBFeNdcdrZ
fvfIE4ytXJqL+FUhTlQrdPs0hcSddEnOXrS6dVfGoR8Ol0zw9UqYoEI5SBiWhH6rfdchcl/PwHfZ
oNSmnXBqfMoZ5or8m9PpqkjpV9x7WpZICq+6dhO9m3NhcBbcVnuSD27OpD+Mc89i3WOaSdQNTDS4
rd6NNiilsxtm9SwUBstZmXTjwAiKsFPlxmuHO7zYEb0WKCXr88NWM1Ne1AH16Lp8W/kgc54PYH08
FRwa1H8ah5/cBA4vvfMPifHubjHiSz+2H/lhWwELP+5cSgny+HzrlsAp/1dki+8wLBNPqVcDxRHv
aYo4j/LVmdAXptqgXebTgCNcf6kspq5wmycYd4zHlpJe68Q1PpistHPXD1uVAQNoJLiv1LoJBfow
ZHgt74nyyrNwDiu+RvM23DK15F/20mm7ozcANzbthI+fsvCvqAHSHB+tjRZV5vx8jeMPvwyei51r
+5Z7N8PRqi83xY3Q7FHLltsuat5Op5W5q0m0YhCIolIJMMxN0oVw5sJ4GOEHzbeg1WDiMtLJPt8x
1q02h15l5j5I1VmB/GWu92Xi7CMhFMDl2LhOF2eAc1U7Cc6twPIuTDtEzylEVgHhTUAyuOZZZqWX
5XXqOhiPBoWN4sK5CeJUMUWaPc5Ooee1hznjSANG0iUERhs59y3JWdJ0Vs2VRJhqCsGGmZtDRPth
kmjGPePFEtZZlhJH650HxXA6PX8gyUf7ljtVHnzDPS56Vpiez4dW3XOOsIJSQZLGR0fXa2WcwHls
RCSr4w8Hk5Pz8U2rDjatsBZzu36px5v44IQsN751DAZNKDrPlMjbekJTCt2424UJtjw82rjBYlC6
A2mQ+y/AHjuvQFXqYiPMd+bFC6hLYS17OIfMmkMSC9cySXgczxmejBZgGRfWYy1LS7qWinYysm0z
PtUUGglVN6Mr4hDnG9igjD3LdyqV1PQyLr8L7M59TOaN1vKanT5d9pWPFZltPJPOwj0zg4NqFdla
35F+w/uI9gUhnR1sywVYP6LC7iIQvJL0nL+EDD1PoBrFSiHwLf6zcy/8k7dB9xzqrhWQD6oX3Dmf
NO2yGVk9PW5bc8AhiOzBi9Qx53rD6edB3owYeoZ1Ynhu5YdEY9vsLU7bLkWRsgY5kGlQEsPA+W3w
zQo1k7CiBzz+Rig2WpBmuvn7uTJOwyuYRXGAZfQikDOm11p1MzV2pmvhglGRKTFCwheIKsgxtA+p
yrMj0lImN6zHcbq+dGrdx2BvIjdXDIwyxMHvblVAC6qGwfwn55AMcoxt2bvqhmdttl23mi2tqsFo
lAqH/WL44aQ5xMIsao93sm+SPxz2GN97eUW+WyRxOhn/RNXTXxwXL/oNMs1OvkYFSzHIX6G63Jo4
HisbheGLtR98ZZl2VDWglocKFdZHXHDJD3Bkeg8WuY1F5x9kyuwFCYDHYapz0YszRjRDs9mBoKhG
+NPfIdAUdZ4pMzMj77Pc9O+3qjUVk6Wy2WNvfJrJaRIas7TPrehmu8VCntlZAK+9uKyQdxPsYj+W
rgTWvLT5w4g4e8biCMAKUw9LVjH/sr7z1CTb1EldqAm561xsLbB6O2xhhiZ+ZO6H/JNsfIub5mmm
AnI8f8XMXaN8tkkBcqrBhTChAvUjkhGpCZc76JXIcDbZZEQUTlmPxm/GiDvgYDn7TNNpc/vVjweL
9qxBeMOPk4RoR477FQ0Z3J6C+cihRSO0/r68TUPNR43qh2PFxbjjQefxBGf5nZAVKvBGrePBk1cA
j5oVRFqBxwQBYlrnXU3Z0UMm8wvYbWU0AUEAHXo+VvWWE1K6rQVYNj/1Jfcva6VQ07FDF0iQkV5E
PAEZNMYxoHMDVpMgAq/4joKXSaeScijLiNiYV+r+0kfbGtFR/8kHQQR9o5Pght71PTuNtB3NLYMY
ZArZj4DfQZU67I4YXYMKS6ESzYZSD9RisH4QMGKd5WJ+iEcTYDiCx8GPl1egCkwxr535j3jR/hKp
fgb3vl/OwX4lUh3Gy1pkgL83Kbzr1IB0m/TiwrCDd9v3yJyHtUGkzUgBrZZTqT+sfn6pPvKBJOEk
ShlIGON+Q3l/MZPGXN+PSJAVfDufV2goGCirVEcdshAUENaI3fkx2jU5XIYLFDKTFpFOvQXVcPSu
5ib0XQpRHmmHDX++AycTwnSXDRLc2R9Z1p4M46O6z/SgKgAlla74axV4IaDhmiaSuIV9fmJEjoyr
gdt3Ty7idVl+U0qewxA2Uhjc2D96Jbtcj/b+BqsiEX9o2PubeadR1/iyMo2gD4Vv4ctCqYafbhMJ
Qi1WPfbymfj1ZpVVqxHbcYWus81wakDWType8DjpsXzPsMy85519S/yVd3DGh3GwB7rWuPTIuDNC
UZ7/ShL7PNu7GkCwhig/KIPctU4Gq7zYyStUKnfDO9JotLDMZSc57M4WmObQoR9VaDR1Yp/Ob4fg
a6ia05LCPwPNn7rb4f4aATr5inozS75pOoqCC0zFue1pAN89CWUuOhJIXzqcdM+6LyQaTM107L8p
meumE+Xq1e37Y1J87AKYgc8N2rYzPrNMKYj4hgGm+hILLWXmPH7Avym5b8XL2LPTaUSZZ7nPxyXb
k/7W7TeOto3xMviEqrHMjftlRwqUlERToL+G5tBV2j2ISaCT+n9RQ7gKZ/UX94aLpA5ux8mYeAIa
ROKd7bJTzTMqQQ2SuOvdflHgTuAgXKIr7yCO8oGqwpSJ8an9mZ5l+yRkOjVQ2K247IllTy13hsm2
nmbL4lMMiw0iMKzXhCHf4qnW9qb7az9EUsDQI5r9a9Q531K40ksZz+EAsWzaR4UWg0Ib5p0Z7ysX
qNEXE584I0agmpzPI0TwTCz2RNww8wLYjmNWN/vtxRHXYNiEkU/Sh5Hc7AsgNEBr35bDuTsqPg2M
7T6A6LfgAH0Zqcapm3PDT75v8Mlni/3nzCgyUhtWUhKZDwX8C+NROCsJPHRkQ19I2qGctn6dQnxp
Kxn/ZeQ0kn6fMR5uGTMUrPhcYlflcGTveecS8hI+rNmxGxmvIjo9rXcv65kpdnQMpLIrIORA9G2m
L3oqNpJLqNioDuIsseKVHzhDbC/C5cdVGRC1/TZEcGvGfh4nKCafNEdWHsPUCuuGlHMkbrmcfoCk
9cyfQIpOa35o0YUQy5D+fufRdwwlqR9zENgzHE5X2hy1jkYvJHWVVR2y72rahbd0a5MLCKw+i+xj
UuRlf2JfBYFw4B13UxxGGI3gdCI/rA62iTIbPY302z4lcWqTn/5gPrKrMP0rKF3iq4srUp4iM5Kl
MwisZJQhVyJEMsOl+NwuBAEY1frA1DtrFke1p1fHvsPnLB5yl7TYm7RxJofbXYsvAYrDWBiZFMpB
TgkF+KLyEN/cAFQNpuUIACWFCoNKnYYqhLKlOKERD1ZzKHof+nuq7xy2Jppp5n9rhK1uZOBEXC1R
xrA0f1KuODnpvB5fcZLt6LPF20StVaVyAYcuZqCrMn6WFBpKiZFIhiKi/32v4satJiYHBeglccL7
kUgQpfpSv6mvwaRyLm7SDSSPWMrx7ceon4smHXzeupLLNTFFcRl5NPJEWbK/ambm9hCKWXEOIClH
fLqFljs3zzFpq9mWI65HZ9yykl3q/TeBZrRFSHe8Wj879uo+PR3tzIXtKomt0BDUAd7HIg1/kXiN
/i0qANnrltyYP5jT7G2VTZ9hzNSN3+2pQKb1rB8FotbzJ/6+bkTx7yuwT/b8xHyZOdE1VfNAKSuO
rFS/JjIUeRzqRa/Ld4LxfwA+qu2MW+rXvnwEU9oSeGQo7qpZl5tVOIXYZmCM+mipLM2djBT20eOq
OAYsjeM2inLRayoL2tT8WAgQAL4jO5TXkNNtB1pvJoqWS2hkUDKiV0zIGpg8nBLia7f8yGi7aFFU
8IpVVI3ZDb+FhtR1O5zcYGhWFjfGZFcDppswR1f3fpPKMGpeJQqQdGX3GZAtlBsEl82yIAwCxfct
U0rpCew3F78gP31MMnr/FMB5YaMGZ9mxxhomp2/l7hg/m+L8efcD+ez5o+DzOrE+r8WYr8nuBWAC
faXP+OqcIcMfNeFPyXLkwHUKzMhhWqYbJBwOR8wckAsw+WP+KkS2tNjbNeFlSiwcfTdWfyIR0H2C
NZI0YcFu1O8XU848Sdp5xzSj4hVqiFEQjuADhxYYnP/ARWQe1xcPakBeLjlVl8qe/OqjcPdn+kqC
RZjGLZgCm4Ko+MTSvrZx/N+NAm1tH9C2/ND8aOgj0tugd9YA33iKPw6cUSsIwknx6Oc8vHLknoQs
gZP229lO5rVGo/k/Z0AGt98TP1bmq/TsPf9PPtozrOOhTZvkRN7UPDrmKskqCwOKoC2bRxLHBZa9
9uWUwfGpf/XrDwxS15b4/gX+M0W9p8O6rBVKBe1i1up52ixBIEcLMNnoYrNdgFTKgTvSa/SZIti/
r2NVL6EP82hNeGCHym0/iT1/kBcjkGeFfg3shhcLeVjlellAQmeHI+rjQLE18Y9xnjKl2AHRZnKZ
Ehyb4SxPHZFulWK48BHxcgffGXfANObTlLlIiger/G84jaWwMHg090yZEEi8SzCs28VcDCypi2Ok
613vnkFTKAnypkl9nVHzjmSPLtagPJv0Q5Hv3Nm0nabWAjgkCpb2vrv82v6CWX6zQK01Ta+M05Kw
jCFz9QV/clQmN0LyPz/YVysot2xo3n29eBezm9iclRZXddgsvcTV81zeL15TiU1cRwlevO/lxZey
4FS3L1QtAwS2YqJrbIfqpA2UZw5h68mhoK75fmX+l+QG7hhGOldFqFhaPBCFUqfqcN+hQ39Yy9B+
MeKlKKVkWKEtWJgnWTRYABeVEpAW05a6RmiUCLVe3fAcairh+foH3kjeKKGsLZp6SRtoBG/3xQW4
QbejR4HbhhYeKNYd6D0QWOGHY8nwwcTJEUHf9U0ifWao0Eh7JCeivGkakyZz8jQqad3u83Sg/pDv
njsYqEz3sLWQW3fB0GraANOpyf2/M2dhsLpdg/EdpUDyI/FTCOTdFcg4nBD6hzJVv3Yum3FJVCgk
fH77vRKNVr8KqRHlUPTBvycwzuqWoV6yxp1a8UmGdKH8EyR7eqezDFPpzodzRUEfWWtwym7+Xd5+
oh1cqrxAFqydlWVldRut/Xowkji60MFOFNedpCh1uSSmojzxCc092VPwahCKD69NZXA9kz+dNO32
Pe03YISNEZHUa0dmC8uG8TfIvG2fSiaPL2/nkgrsSNRciEpad6fM4CNm0g3sTcWINUdj5WnWBvK7
XJg/x4bKgsxdRbFLW9mAtJ9dMN1u8BV/cTqDllpzKTJd4tlenAKwldCBT634+/eBncokxJ18iBTB
xyJyYSIvXxY76urKrBGgLL3dtFvnYR0dMkschDc+p5FJ7Ko32XvHzHTT5ybbmyvVcR/8gzVAlRhr
y6UjVgGRBdViKh5sWxAgjD+cU9omU6bG0/EzboLYr1F2kQy3ssV2P8akSCB19DFCIvky+5MWNyDl
iIH0LkrusKqWMSUVymVk4A5Idt2Wr4z88CZ85PdAA8ioWmZhO/okvwHqtv4y99LA9ZJwjKY6jrzd
0HGO1PyYUxpgoTNuwPrBwoxU1RcLodB9tlqGeJUVQd7213ZIrYY9HfO6irU3oChwrNtHzQrRqOGy
uviDjNR3JYQ6ROk6/TtOeIbu5UtFO2uvdnuk6As62krE/MlIvejSQC7yDYHdGoTzsnflgjc3rOkt
XNocdnzzB16d1kgdegp3dGvhD0TbgmyhLM+Zd6dTSTuyei2HjMMZf0ZGmocgxbm4cOhW5Zwl9PdR
1Y6HOeAOzc+MwikqsYhkGYp5cVhw/ZPE3uuIa1bTHMxe8RE37daOw1qE4PTRy+A/0oizBOJhgNW6
O9odhAqDl9n0KXfCuO0KzL173Pr9JaCzAuJoS7q9P9luH9+i7ylHi6hKA64nAbZ9gPtnJ6rmjWJk
MKKzIkGqc9DQUK5loZYzo0o6hlL8pSvCTDsPCsML9I8DKfGKuadUHYjf/5gGFfzSfH8DU2yWOx1b
OGxIEBAONT0Q3iYlmlVyEzAk6nNA1HNNJICI7hTOKaRs/u8e+D7v4Yj2eAjDt92DzrBYfopTTaMM
uRY4wJ6i0ieY89/sFEsf7X+g8PcSFrQ7K/dEMxoEJR2QGrPr7mRyH1PjRHMLDjnIjeOtM6PydMCO
taPFrycGNfjzwDy1fl7s8h2PmynZZ17kdNLhjDQnBrSJhL8y2iIEKa4Ya+SsLjLEjMYR5yChzrfE
6bOYO7z+bYvaPaxIjc+MHzJI+/ZmgKa4GzmsfUgtcY+35VRWTi1CLS9JitdDTjBfF2cL2Q/Py3Hd
bFmnRL4OF/NRoFGA3pzvBYKAKc8llAHCeSuZyu4zbGECz9RGQAcUXX5v73PNQsUJ5/RRK+zl/YlE
Yxa0q+FgC2Iv/SFoUI8DU9/oNYC9zC8UbFxXQh303itoIYldQ7ngEDONOKEVp4UsUHjkGkzX6Z/e
BlVDEDTmEjTjFwBJ6YN+QuhgR1k8r32I6gnMzfKUjm7v5FOU/ybMKcmqPDCYjbW3t2jac4BrreOk
J4TN2/dVFlmfCpDvFlBNVwb2EW3OVzLR/0ob5XP4lcJNeUzjLLBIT1ONFowkwZB8XmXK7/lCn/G6
JC73SYiwzTeUJ1MWxBuoSBSqqjQuLP2EDtgiK7g7eHOpunZHLJNI+OMC5/kusbBV5ic8kKwqRbag
eaOSaK7J0qjy86HakJC24mhpcc7u4R7mD+a/6Nu5dFc2C27agStI7pbULwr8kfaQweCHfSav70NW
9E6Q4dXOqoivJ9CLBkoeglJ0K/URQgy5ELfklGxvN9v6TjAN8pwEzOnBYDgsFkYhffIM5JkSrhFb
nFhQGlA7iRBU7uDQGuypQ32yBiYr/Uc67wUHyJwYE/vIeS6e1yx4dVOhB1hPpwMA3cdtu86YsjMI
oW25OZF6Ga/ec143r4/UYzF0MfSR+wjKwYANRweHNORwXN+fpo5WJtZJM1oi8X/scN0OvH08Sscc
bRl2bERVADQggmJQweG5hgoB+CoKynNbTHtkx4LrA2jbU84lm8mH49/h/stalqddfnQpg/F5WpaK
1Ma/fdyhrBzgtq0btiqP/uJa9LNATcx0C9E6U5ZQYFaglUi5xvGdvQxXgMkM03yhugoFSnVgtXue
irm4LgQUcdM+Jo3ILmV06cENlUttLAyrp9leZa2L1/CgtYG7EeRGk9ppPr2/O61BsXLXuPUZB1sF
YtTrpzrfWfSM4FzSlf6BFcDaC8PZv6ge/doesOQL3GZK/5YKGBteU1yAkx/Nr1FRWhinyBLLUyDq
guehbvHiNRm3E3ywd8m4kd1YjAFAX4SRC7xdmY5t/EDdFSa3PqzEdwuuS2ZLjGXnfx46PhUvJiOE
tCCgZ0ulqx+w8nw5R8Azg0XQRsNdqO6WjEmG7Ql7NbvvnCgY4eUoVoy1P13LkjMTH9bmRGTg0PaY
IeXnsi3aw9krJeZHb0rfwbqV1rnrtSR0xb03ftDhZCqseoXVf69XJ9QObhw95m7+5krJSr27pNeZ
Xb6fNFhz/TC265/nCZFO34UM8ubI1vm+zCk1XsJwMC19Px96qz/2fX3tEC1NkKcXG5y5oyAS+0bc
JcMAVHCxUzcc1IT7k03DpCK5uWr6L4QDiaZTbxJnpSTOwtxpfEhm8YJLlnBn2vJSI+tqX/2kISRV
avdjYN+ik1qPBgaDYnGs9bVbiYKoVHmTrFZtIaG54cN4Bl1Czwk/UEeHzcVTBSn5HD0vAizaTspq
kgfzLG6KUewbhxSUCbNXv/x0FazeisoQzBPWn8CxiLhCsOMkUp1qdtd1m/lws0u6Ftk1ZYOjkkYN
y7OKCGZFtRGuk+iIV4Eqde7WO9tv0xpanbpLzX/qVbdyJJWxIlg3zuTDhIfA6IMjnm1ywEzYXXOv
MRu5UwjYDsAfz8fWMkkwpuQByWa4fyj2PvTX7oVfyrs3Q9rNO7YIJ3Fwm5SQW0EDgIDZXL1mJHDs
8Rm7jSj/wEfTpjOIoP95ysOlYlaR7nmBI/655HjdHQ+YmNk5o/Fka80f4jFwVPxHU5NdPH0uJqBR
xMLfOtrpmL+1zSbikWqR+wNilsswoX/eU1PTSlAjtb0jktkiFjNqHI1HDmO2yFgXXWCgD9xK1u68
oB2hq5HOxxP92Y3fordFawPZb/cvJ8M7II2OUC/yWkfCGhjAzpAXeqK74QfMOBnQzRq0rnhbCrQ3
+3bsTDmh+g5DtVjyamoG7UlEKUUAsgayBBseAGS7kdGD03mrX5P1Qe8DwcPVP3u0iU3LP8fD0aBO
A2zfQ5btLV9idolo+TahISWbvCFAKQUUl6Gdc2wwkw9sqjpq3aym2lqY1ROM2ANMoO/7k1JB33ez
06LpCfpgufMhCw8ZcT8vOAxzWaIfwL0As/L7oc3ZJKlGoEKhFs/aKLs4ZsnIHO1FoMA8T2n4Pei1
x1B2jqEQbklwqVcz4YOKDV+4p8FRoHhfStiOEdtdSOXPnD76qlAgXgYpxoQbk04j0XMtaBbdYGRt
m1zP64Z09vGi4mlzOvvM6tCfjZ4/nn95YFMlsiB0PqZ4kf/o43hIrma20e0ZJZ0Itthfo2RIQc2C
0/qR00klGiIYQhWCSuIKTaDrOyHsfXA5JWcYZ6HeZxEpaC0RGI7HRUfkyHwQcEUCL8yfAy6Z8Z8O
7vmCD3NCaifRgc2S3DgejZZ5V+6ccNqh5+z2vO0jkZjea6ooDKtwxq8jOlfMgx09FzX2ch5WVB9+
QgzSfjTAyBLvBKjf0/+IyrD1KXzaYqZ3no1XLDenu+fs5fP7jDQbBPR6GSQ41eAfEe7RECQOFkOd
POBbMtf6kJCpBStvQTXk/SW5XWVxqPqvTSby/Kp1ySSYdhe8IBn9pEijugtdEVfclfSiK7IUSVDX
FXCPxI0+4ov2rUPcJc+oVmaXxF0pzqQ12A329jnvCFOYYoWgSwHvw3gzLewtbJ8SRlrGBUr4JBK6
57FJe75+eFZ0KbvLeQrDxWbm3SUJtsO1kkzMMpSJcPC5Wk/S+ozz8sREbWXZph4ac3FDeOrtbxzl
MRBIsiLT6LocFJLL+vwwGQ4wnjfa4Fs+iBDCf2yq73Tv5ZVNO61sbCw+YGn5WuiRQ7T8SrJv1/w3
pWxAznbvIeK3Oaf30BCQuu7l8Dco31TY8Q9xUaOWyDEXEGT9SYsSnmiIdnW9nyNYkJt1LmCizFkK
+gwJtikzVjTav9ztgw/jAaJ0Ej94/tdgHDZxbve5TYeqEs2Rol+DwtuqDmk5DlOCTz3PAccp9LIA
f7ERq8T2YpjgOyLgAmrX5K3Z8Zzx0tk87QrrtV3M9iDn5x0RgPr3O/o0w3KejSLLvaKsmqUHYaiw
MJdYZO6dV+1V1XmtLHIHSdl0LCMLPSg6ylazZXPihNMGOfe0fmsT9nZfsqfQcVVzJ0pdiT7uKZFX
r168cz/ZX5i1Crr/+zA3snsQo9wgTjhw6l9rSvTuYYUpr1jspx8b9vuL5Yj0XCCI1WZt50h4tPod
gDtmyzrC/esF6hde+xVJhTWvcP+x84Bput5r0WzxwA4ot/xNtCcuuSA1oIkJYiie7lEJbYL6vSJR
4wDY2jnQKPbxkvMJNXFF4ePBYwe7UPe9vKisHr5+XgOgjl9gkv2nvVZvAtLXQ+Ob++L+S30sYOIS
LtArRK/YHpanusvoOCP/yCV1rCOmZLBfChFPsuW+jN/pu6IVPGiyF93byoi+En/p50fTwdAEB9Jt
wDKo/WXxB5/MS5PdqCdUiD9T0PsbgEfk25Dl9PhHP+Sla8DsgrRqdd4dccFokTrKEJfMTaO1LJc6
UIdux2LWqHbiNF1TK6nOYv6ZrsgeJRhSHA90YhggvcC+cSI9GR9yKFkJLisLCDbCfYzIXUFCTZR5
FntiAq89ca4d6RoR8nqjTglXnZy3uccoFHIJvrVN7B7k+1RxuvcufMwD7LguB2awDyNDPWx6G+jg
Dp/SJrWKcIccBYCj13ZJa6EfrI+6HhldkD+0RljTKmEW1qJ3jwoYviWO61Gw1VBDtXVFKvFo9vQY
/cbDUnYtwU3Q8iOC2taWXRTU9jgLQN3zDDbDccrCLtBn00zJRC77Wu3mYCfkmOgjGwg57h2T7qtJ
9nbz7c38AjEgX5swhJqQBYXkrcBOLvAuYzv5TfI2TqAsQ5TSuwQhvs+zJst3Ycu+MI4HR7X3gYW9
yXbrDHrWAmdDSiTsML/wU/BXfIyJVgAKWOKL4bFTV3n/X6d2CsaUO1+ID8RfCDcmH+bOPnR+J1Lm
/EyVpD6eys61wQ5PuYsZe9bIlwzCQJ2K78tLlcu9e2M4rsVOaG9g36teTP/fa2sfOkmY66NHVTYG
pWpEfyHcQfa833nuCx9S7CbwDcFPkw9xv8FTfxTC346vkt2HrhIkzfXFNIPny6rehTG7R0R31774
fssi0PpZ2DnlJv5wgV4eNB2Yj/rk69pKjwvJtQ2Lbgq9kskQ58MwvG8+5I4dihwXNmcwEq71w1Rg
rTu70oDQXmR90kvWZn2A4Twxu9nVWM6qOqoyiNSDgKy7sthIt2k4bVNSsXtnQY3ZtO8/OUpKJqFI
PoBGakYqko1IcoPNQ9T5L4hNuBFhRsUHjpTMqKnxMFx0t5yH5a5Soi3oMt6BthRE5Nhiok69BtQg
7y6W+NAEVJFRyiyMD732rLfhUDihJUYAijsQPU0UmUlEhfK/PtZsiYxFtyUds2bKf6gFhVkkBfsc
LFV5SgIZPOwSS4kragHg2IytheZRZfRgbaV92ytw8puKn4WRPtFvoCN/DtBEQJ7oXtmMbYXyenRC
MQ+db+rhOCcy6eTsDh6F7llGrPifAyJ0E6ju9qK/C9G6JImEr9cGZYskGKjijq/GwMmxEQmMEXXk
Gs1ulivYkAxBfcJpoEdQEDRIRYgpgijU0wPGyqY0PbZejD2dt7xMDRtOE3w2LzfPPGTJxRGxinZw
cMi9hdXw/TlDRXjqbjrJl9HgozAyyvNbYicX6l0kafYweJS9HTUebKNfjJih2zj93GeDV+zKqTzu
xM5I75VAIju5XfCtExeIoRmQpautgmRMeYzRXblGJON/jskpzUA6ODwaMTL6bhZvan7eC/ibTUq6
KKM83K1/zE8sKcFUixLbOaePvgEQFh+eytM6uMHbScA8UoMqJ99E4bheskaF+hDXTZEfxKi1x3iK
xeBvchqTe5nn3r5aI8NA1/jiAtTd19DG0C8xgg1TkDNOOPju+xM3XdDlqMUAT0UK7+lhrb3p5S/R
I4h447yNVojxK2/QJOqE7nJoK0NDS4Bpmhc51vilAzWddibtPhokJfb7gA8SwUAe3ZQA3vYmS7Iy
2L+5T7MNjMmEG0lPYP8kUWf2Ls5bhzU017NX6mH+lmEy1BDGakIEs8cJD/KuPV/iQ0jKcRzV61u/
j0zGsGH6uTEgzfjMZtLfv4qkycot8mAEN/EvF1msXBGUYCDiAHiEpq3+lCAYcbzBwQRqq+tA1lk6
xOpK3mXcAuFkSsZvmEB0x39IXA5hlLvrbdSWNn/W5W8desD9xzH/ZwINbs6ltOWc0rom1GqA1bD9
W8vMmHAg8AZERk/9dxQqDKudlUUlPD137w+92NiYmRH7uDT6jGtILI4Vp2tflCW2wOQ9nxFpDvc2
vrA0uB5sOF7kff60j6tvmowJ0RD0uuOn6fB82BZr13RqLtniawIuxXqRNntxnS3a+yNp2x4VpYYr
iQyUsZI1Hgwxl24B+71uZesZYxhPooJmuLchnHRvpkPEj8Ux61Zy7SOj2rT5rEkgr+QJdNd7hvYA
E+82e5gxtBAfGLCEQBA7haJ5F1AOhNpimloDNIcq8EHBzwTT7ZmJAYJWaHJJLpCu94QQmEIOZbti
1E6HTVD2xgMed6olOyrZQQ4xiL40c0aqLOiRLfIHbVZGC4sSeUUEL7CCHHEOGvPiq2Ga2/M6snzn
PoRir+HvzBGkzwlSH0dy89ZZZDj+AaVcdNzweZBBmBlM2ShGfXbxRBD1g/8kwHOrZTzI4ybvRdh+
WTeLMpnLkLhpQtfUiieqI1mYp9YPZSMF3kbZlnmCNvmpW7/wsC2E+sxGIwbSH6hJ8vDSu+SOncG4
ToYtcUh7VW7XziKPE5RseMLvmPlKtDYTtImmlM8de+lYW3Oa+RoJj2Ueho4tHkJDfsAxYFcy6QPE
KAzDMp3XoEB2s8mOPs2NNdV2hXEN4ccWoovq+0blCQ4B5Q7z1ScYpBmluW7QRci/6snajKkEoMU0
q/4WifIDAe7D1a22jiO104HAoIMlGwVvkMWX/dphmePupStFEpi1GPki44n0qxYdL2ZGYx24UTmH
2PIiED0dnLOm81HUHAxjzsZM3BO7g69Wwy/ZloLlT6ekPqB8kLnY8+Tax2IbRln70dcrdF+YnFuV
JCyi7o9dOrkCH3ACocvJlwGkask97T9KLDg4afgWgKzY2RAh0S22n5iEuOdHvpi3pNBevRxgAvJT
oYs1ZFFlIIerSAhTc2DmcV7N5TJ4eBkoBVJw+Kv6CiFD6fPFENZ/h6tw6QKIFM0ctmpwZyaUYPeq
k0R4SFg6ZFhFSFhqa8xBFB9FtbHZNMmR/XBqO5J/dxSHdrp+K2XKkQANqVR0z8zDgXs9cYJ3eEsR
930l7OaXw5IaEy3Mg48FlY3PFxXYj9o9V9z0dzUEAFJoIXctrgcynzcTeHHEH1FHwrDnnBFqW9R2
eNAC0Wnl8Bqlt9cW8b6nN9SahrYHDUWNArm4WXfei0D0k8Y/H+KKVJcuOsbebqKeHH2xNvkqxmcS
nemdONZ3F3SC1pTM7lZ9Cu8xm4oPslpDW3LEwwPLJFUIZvq10tNGRgNZpTJMHKA3+EnC7+N62+82
pSZmR+nrIIZbvM2ShojC+CoKd7KkB+faE6uFkfM4IWqPX3Zklaizha/TpQNGfmriN+9jF0JlA/8w
LUVkNznkZFZH9jqrZ7V3PIz1ZQTO1d+rLY4NSCAbm8P7TDsHmpXNjWS8Y8iiX/kpcoUvIerXwE8+
unW6osi9rFhA3G7yYiaCe98Nt5PT+/xIf0UIFg+FLG0lqsgCXSXxst/dTN8/akR6DU5jV4+djwPR
p+E9eJtMiM70gDHs5AC438OQ5N3IWtt4WO5KVec7Fb2+iDMs4BhzHGRSwv7TcZ6SZ9z5TlgLjbYx
3b5b+7MdTRcC2x/CetEa8vU2Z5kJ72LOgl2YlGJICyTtzqjJp6UnTOaiEAlf/3HUyCILx2YlHDKh
88HZa8cnHslm3oYNc3Yi0ffzFUbK79DySKXcwLhHSaXOtSakEq3FJhhAuMawubkaWJeFuWQlC2Pg
NaxPT2qPXDo6TqQRHILhl/jdr8af2GwoO6/J1KcQMK6OrEwIrPaaAs9sK7cfqs95SfuaTxX9m/kV
aVeY2QkxEcxO1Wm5Jc9udcooyDeMKz8vVAhJtqgjm6QNYGKGurtvhsCRujbLM6VdJvhDa/zdIbvH
eCdtq4DMbrsSoah8siM5YZ9KC7kAeTpf9A4cH3kOyN6VaVN68UAjqFRS5JgyjI8GF08z/Sbkyvlg
M4o+/LJ5XD9uAqF8761Rey+Q2ZIgMoZcVKAH5ODdFTLdgayXylARsplfp+Uh2o3NKgonetqnp235
8IgWA2qNCZdSZ13lyvo2LsbHYj4nZFI9sacdDrMk1x8qaVGKbrCgU4Qb/ISPtomSdjVZNNgwAX6K
CTnV+jroii+fCfTMgUZ/T0yFFPhHL9dkZkls/nVbhcyKnavRroDi581XKmmInP7BWhFn7lg8x0X7
sQNcRUYYCkRT3wQDNdDxkXOKrzs+eFsHsga/1qZadiG8uhvrL9GYxUhywqvYcczmRAYGZmPsb+Zh
HqyotjiU57fWmjTWoadxWL034IueBy/Hmy7IhIEGmOm6JoNaJ8FmHJeigXRc147tk6nHecRu6Aq7
ySpE+kLicq8mCyViCWeHHaJRsMqSorH2iIjQ74hc9B1AAkfX8s+ipcGoahQfGY+huOulNigrruHY
ghcNdjQXvcJyb5SC5Lwf4PT3A34avu6VPD0YAI7OQvzvqusZe3H7bsy5zDVLD9cxgO+k/SJSlaKI
aRRqjMmZuJ7qAyL01tPLpq1Euao3byEtBu/x2Y4FVvRwpqxVkWxa6gUq6J4Za8TsK8cOZNmhJ5zz
ZZAsHYsL4rIi0fvVezczcU4iAkiV468QVFnSRH4kx3MJ4aEcMkGdF5+vfQuPCUAV4pYbEL+7triS
AjvoSdhCQI0AO/AePQH8HY7DgUB4pLLar9SFDrd+UHvUAh5JiLWvwfZUtIgKy6SEHteEz6IVyMUc
OYOBdFyASKAb2pnRs+E9QpBZuxJYYk6sYubiQ19wUQTO21PcZYwMJvvRpq6pX+OV1s7wIzWVXM7b
hTDbfI4pQ3A3Nb64HivukyQSIaKIBRS7t8S8rE34AwL6UjRHbT0vT/ollPNQXySPAw17Av2/leML
nleO+I9vsHFvX40GqfdNjf00WMtDP0BBJPl6wEH4PKSZxz8GITtOEeUAOoOaghUETryw8tfH6KEI
CxLBsjNPZEKFvwbRVRGhsf7MaHPliCqPNahHN6qofwf2GhWobQi20C4Fs98AqBNIQCxIvP34+qmC
n6fvKGkU86ZSwuhG+ZNdpyGW5v9/WML9/CuuXQqzxlNLlUm1B/L1asWtVbcrEX9g2rsRTWJ7L4Vz
1mv9PWXBLnXxxF2ZuXKAGZERJwcP8M8q5+9aGxvgQShidDpGxFM1cmmROeqW/xlHqSo6vJkQ8P/I
KV/I8LSmNWQUVl+T79Tj4tQQDt4t5AsOWBuxg2bJ8ILCIBhViY08aT9THAxb+RQzjF052unQ2mEn
8e8rSCMyyprZdpZ/1vWRuXAkk4tUSmaF/wj5PfvMWQ/r0TYwoVLm1LcXz+rZaWbuRUYA1le379mI
/6oNquKjmCOr8knuuysfKMUKxyf7NJOmK4uUoLHtmmEvC1wFnSNKso7Bpodq1wGPCcnsZSbj/UXa
vMSYO+4js8x6HEmHS5I3VB002sZdlfu1beBJxaiEmBLhTm8YmAXcTjPBs1+XTVayMj4E6SVE84Hz
FMvgms9FREYz6En02Ie5IJq896JUe84X63Lj841yOeGmWy9lh2nN/fPPb8mFjxPHXo6bZuUnh8Pa
KEJwUMyJme4p7foptqnuG3UKshcn02QFoqiQ0eH9GT9rnbIC99TFa4ZCYTMODp5CmkfMfqJ+00zx
IrNuAe4ROdn5u9oxPg6hsMOeFKeMoFIyi9lMYA+JmNTI9jFSIz5Y6gwA99dd6kcaoA1ZP4Hxs7jU
SYOMD1Xorscl5xx2BzIGtxJH5nuwgpSBCT6Em+lF1cOlqN0KKna6BlTOgokpTrQgqx0WO5CqLaWV
INsNwjYMEELKtwqZGRPH/alARSIywJ3gKGYTB8sgr0/fXTgov9ib1EZOT9LHtIFGOG4VND5mtTw0
64o4pwZ+FynWd4sxbb0v5XyYovvpx6TxjHAb2vaOtw7GrGuUUT2t/dH6sNrz1pHjylh+JVBqwZY4
Wrof9673g3o1kFAaJ8rpPnGU0kX9BkIUHn9nR6HwNqvL1Zu0+oG/gao/MC4HtCUf/Ykn0oGOkyCC
T79O/GuFJZZu/2vOH1omW6pBhSBGfzMuZkn8Pqz0uBpc748QZldul8Wb2FhRyFnrE2mNcCllEquI
8E5CrDSz7C3FPRIrx2hKpBwL1L4PKbrKtwswd8yS10vPjfyXOVStOLDUVpp0+HzohNCJLDJamlrp
eyY+QFkFPtSk5z7srT4Q3Xt0Qd58J01PzkzolZaOR+B2jZ3PUlIU7tr13Zu5ghDgYfb0vDCFKj46
e6o68W7QAWTGbye9u7uVYIUxw/2xBAYm/BwK7dr+Oj+icHXKAjp8vrMfdHdpJ4Jb4+sxShpGDa+C
0QDKJdpHQF/E/4jh5eIL6pMgNqPPjToRKHLpey6YnOT1kl9w+EeJ5SSUrXBq2EzW+Gp8/EekOF3x
EnU/rRVxvcW4/PP1HTNObim2KOvjWPZ7Z/bIlrh+9vQayAeYq9HdRdHQ5TOoM/wGY+ObWHBWSKLJ
we2wrBV94W/qz4WB/3+eEaePNBoeXGYOZGZQ7zGyIWFgrY1RmxMs/w/lFHX3qiAtrfek3S6dqERG
9gqOTGlZNnDjKh/5QyYdMrM0fFRicZDxSBlrF/LqVs40ExTyf4g7uNdRzTb26Cgdvnr5TXx3wZul
T7V91TEzz0nM2SbRKaVhM0ucuJ/wfJj9zMhGZwuFbi+3eaFbvsMWgrDwONMnYz4AhxpPDuSAElZJ
zXmy2uJxzIRLy+pLgz1CTzONQEGQK5cXCO5PN1ezku/FohIc1VtuuiiLuL9Q5XOy2OgPqU7FC1XW
M7RiiWXT/2SXioF3PTxZP4GXvcL6dgGMTTsQ4WcYmhYSrjS4bA0aI/s8j5eY1kN+cMyVNJByg5Lh
RvhBHBDBFAdtzNGUBNDH87wDZ74NKs74elJo1YSDMv2b7klRQHw2Rc8+uQvCvpuYNxGmy/ZlNXGl
MXM1BYBY5j4Ez/yvG4F2G1ejIrH4F8LwcVjoY/dxbzUipM3RQ2lvNmkbLe6QYmRAU15hoyCY0U2H
nZuOBuBA8ee9asEeI8FnAR20qEMU+MF93r5N3r4hf6ewrQDs/LtwWtJcJhn5kDYnmj9w2hXDxeMI
6qHi50fQaKtw1uJtzVLTe+4ZYDaO9TryNR6+pWmAg2oTQZqk1OZoY3tq2PGZMYuC4mOu01fneKxf
vRtNMKnq1kWiMw4pjbPzpmUYWvMNqalE7Mcfc8c0vr+sp2NRtdFaCMikL2Agzimsjvr/CrQMrWWQ
9b9xYpve0jLGAetnv45Iz29qGtHebrsXPhy0wbOM+VoaKrpBR7vtFwEJN36/mEMOMGGY9hksNKxC
YDpAS1zHrbBYNJDwl6oM6ZfCCb2cUUlhlw9b7RfHvCNQtFWci/kjmXDKL+7005CM47ESqgnxrz7K
rvlqkoXb57EkT6JoNOzjXUdYR0BGvvwqOFchCVhdRWj3cGQoI9qrrIqwTOIKOoxWdheqfMDJLQyi
SvKMzv1o+DfjygUWbQT6SgPW4Z0d4vXyHTOumbSthjSuDcCHaedBF1s0kPxgXzOpfjX5SiAPU2n+
gboiHRucS2naDDo/t1BsRqcJboeCxCrOQoTafe8XYfcOZ81e2qu20zvW1AnSWldGIfNuqW5Xqz5J
/HX5YohX8uxovPkyWu3yE09oeq444DtogTiAGxmcV8hHXQWZ/Y6zYDX0aIur76z5PblwXOnkHLHY
2dPw7b2r9qzGaPQpVZKSi8w0daHLCx03O17ny5UF6tsXoTNNNgc83PNX1Nr/VRou/aLQ5yl3zp8T
Z41mjAsnYxFUNRInxZMplVlEoD6O6zhbsEjbRUYpSMxC2hmgQJfABJgl19IYlVdeafev/LsX6nl+
9nfTVdXg5t3h5qsnFkKZVjIOEuLMYTv/xlmpSMqDIr3i1kKypcJkRbFyV0wWyEb29eg9GclcumEn
reI/+uHB2229FrRWxHb0flnhbSpbOYiNXxD/ruSWFwPq7DdFdfCqn4SgwG3efmeC6Aj03pQjt2QO
MFLIhShaXl3vP8OwtOs6CBwbJ+xav8N2oa+6Okd0ZfdK5kDIsJ59KWQp2TqAsUupWXzPHK/UqeCL
ocwhCFgy2BdYGKe76zFj1u9vxJyO+qPuUr9soGNbhpKXbeyo5Sk5rYGIBKnFSk/f4UCZhw2bBYnx
loVNUeDgbkTdctYlKQcvUGRHT8+xH6N3IsggON/tYDwFK5S+/TzV7mkQwfIDayF8lnODfn1h/wUb
wr0o1t8d2Ty6LUTib6A7RESTZYVcBTEtal1caf2w0OEcf3BFteNWtlAPryT08yu2IMHHEqVf4qFY
mXQHgWYZPOp2LLQSfIrMJFIhhr7egApF9HJFoMV9mTz7FHRLREd+JviT9/fTEa0bluiQjXE7vEUf
72xNosOVudHW2k0dX5rxkX+XeyLnWxsvIyO0RrtnPXdyoG4N9+JxaN1NeFXuF0bxGNYQ/mHFxAT8
fBp02EBwd0NH3D8TA9Ldrsc/aUMl2BL/wB6D0UYT3XQGhDTtwtE1A4Sxi2P6ITLXx7EZORJUlTOq
3HC2v345UIEw5PywB5ETU83tkPF6OMTjm8pxWWjrtsRkqgVUIv6/YG6P8cGQ/NJXXhntMnoAWfVq
MEzYlyQ8E2QIih05LvNDntqxRdFPNlOLB6EpqdSVYw8a+U7ZapB7vn0k3DFIDvo4PQv+orvW0Qi7
fJD/fxqL3dw5bCxvJ7Z8SIuM5v52KqQ4EKUyzlqK8jWlrOp0ZD3WwW6kaV1w1NwnbgvC1JNuTX82
nqOX+6aC+Ib0OiIbw3y9g7IEFRdLvlG0YPCQEC0xtECNoiPydWVuybmtENquTSJ9hyRBOLIQKwBS
eN8RuOpb7wd0+k7kJI8xJ2llSf2YCYL5n9Q4Dahav1833JsOJGHg2IxbS/6kvV+5K7O1u3jKQF1e
Cni+hvbETcYH6ee0cFS9QGfnzukDvU4yvMAZ+Cv2IWE4mDoJfH4w5CLrJESyhRrpRX+/6n7TIQNm
ak0EOF9YJlCmOXu78r9FQx65vK0dYoI4VUHUkrJ0yCTWgDFKEcZJuwrfQ1EWgHTL1fiOj0Xx23Oo
trdJq9mFcoYS9zoGKMmYZMg0WUbakYoq4ov+4iWZTMThhkAz8JU2W460iRiAMDZRwXC29zfNIqF6
HbcpET1xetlniVVnDVKZT7zpx199rh17DeTjuPf6ZGmIrr2vd9ITqD9C05MOogyKh/eFLZzmOTcX
SlVdAtZfxnLq3yPKU6k54Djl+0LpgCHpT8sZh6sVSkUQi3a2+dpZZopL/aLetR8zVapBftjmAEEX
nNDw6BmJI46mTY9qJMBosB2qtKakYZPLSuBUD91mN5c5OziJhva34VBohQGkwRi5rSa2Xh430nLp
khw/AWNIeQYClSyg3EOoH0/aJ8e9wtcnEiU8BqA1QaJDJMW2EltZBydPfNit1AVEB42itjQZd2gA
rjTqbC1DO0yrE6m5ZrT+RAmQHpb4ci7vyOJZWCi54cCBHarwGgHyE4FlYQMgukoVA2hA5pr0CXwL
9xLlZNhHAaD1zZf4z2HC8CrEwQYwFs63jQtBZNGmcm4H9/X0Bd5Kp9uKh0rrjuLq3q+jXYnpWnwM
c5I6+QjfjU7ICeE1DPUkekdAtW05x84/EWgeYN5N7pW59qTugbnzwdGUyWgd/xjmeZZMuKsuRI0h
yJC1LFwWKzV4SFwotZgpZIX1+V0+lZiIiuOZfNn2Aq/FTUs2gQ8rYq9n8wPjCZPZG2rmyb3Y4WgJ
IfJlNmHIQkiI297xqyYgpzEH6Szo5EswSnWEX970VD0/HkS89OGfhqLQy63imErsska1ZAAjNcqL
M459mHVj3h3g2YTh39cyYYsST3HKFG9hi25LRhLFxFmpvlEbA/+mc9Z4K6vqf9p10QZh36q+g+zl
Be4iGV56Pb+sWEj33G3xoL9qiyqusE2B10UP30QxF3yfST083az0qFxBC3O/ucBBnLi7BN10j7ls
7te70veOkLasgbUU4mBNWOQ4cWiNWU7ho2t9Wsqfa4+hdgJNytQyvRkXHODrFXDtG1owBcsW6Pwf
N0Dx/6/3DF61woZyyuEAKh229PYmW2N1sakRmpgsJSVagAgwJjy8zB25CA9uHWStfqc022aDEiL4
B2JTtTnTqyUYXcdD5czzVPJQ4KPLBCFmcZ13bDPt84iSugCwpwkmAA9XksnV1Vc/YUraE9aHZLg+
a4bTtr0usR4cU/CDO3AsJ3rAEXtms6mOhn7166kXidQr9d7FBDUd3WgkU+lO9CtMCm4R/UeZZJyi
l6VCizyCV7hD0TatILfpWxAOyXiyLU4MCJ3XrBheAa7UxRMOsn1Z9d35ISebLac+6pYC9yt0ar2k
d8CpWO9+uUhyZnFCFO3mpczIboRA1IaJ8ZvR31GG49wai9ncJI6UF1A4Ba7hTzW13cooWsxI5t3m
ZpjdKvYyKshLO2rxos08XvwmEYMpFhPVnjCq951XGGI/9GfBn15RzasTOyKd4pAYSjUS4jH855wa
kfR6P4MFxjDL2dpTp+AkOYLx8Rx6o4Toae3wMr+3TGP1bUbkSjKVwwY2mViwPhYrcbchEJxJctBy
ixjXvLChJcLJGuUXPac4XFdKY9jZE3LvvKG41fTHvvGPX18j91C+YsfyRbpjq1cJloywAZdohfdv
pJ5fmx2X5jiq4MqnBq/Q/XucqZ9VIaeqU3a2t2C8sdIw3rNhxRWBSasJVMKMRFq1hU600Io0LfBJ
WNT6znVVPCt1gQtTsPiqWJju/l+EEAJax2HufDM85PbIqeMIDE7ncCMG4CjtZVCF7K0duslFp/yi
OncT0d3cXRCeC4t/fjtqcY8xqqPAKKuCHZ9to9EbJkbqP/SUVNw63r3qEZvkLn20K2RwCgcvZlsp
ul3rmAAIYRdUn2FwYrmwFeKvpA9DLXB5sO9YoArun9a9Mdqzh3U8xMa+zryzePZFlAuGaLymnfYq
Qv1xUm8CR+Q9Q9oEj49LZNCOGTesTUwtsuoc2Gj6njOYIC+CdMvC9/exwSX0kV/6tZG9BwVT4K8h
byiPgYLoMOwl2hAzwjmapxBOUFsR8Hbh7V0705IcTL5QBfWZBQL8Bw+xueSpGrlfbfJPyncFLYug
Ky3GLozHKtXks7X14knvPII8lC3ZrxWpWR4a8QwQsnzBvpwiZLvwlI/SxA/2NNmXUrd4xoAo4ZN1
E/crv8JBEXeg7KginAuKbpLwuwmjZPcdxJpEV0gsFh4ZIDa/tT0yRjYmTchI+14c6VfdazrWRvfq
kL7TFlPtqel5clD+4ApphQaeRSzMJRW1VGZdd40cXOoe9hUmsOEg8vdFYtY+RkuvN2le8sYb8D54
n38dvoGnCbFPUfobcEGxeGaLmsehjmtTEhccpD7mtBphD3pgxxC7UtzbVnW/VDuTlfFuxrhyUX2e
Wvp9cKoagPL2SUNNVcRwHaxO2NcHG5JRIO0AsTEXWOfVFK4w3TvnnBNl7qJF755TMdWbBm/F76TV
EupDpOsIb6I5VgQA6PFSsSAvSelzutZd0F/pHE4iohwrFxeQzQkGtke1yk1areU8ZD1vx9KeHU/2
l3TDZTOnXWKf0noL/Ur8NdI6tnMJ6ZmbYFppNErKY7ie6MKnei/ob4maUYdWn+ZQj5pLdqs7qh3a
dirvO5O+wjsEAz+rJqAL0exT1GpyonVxWUEXocGktBHyixEEKCdqWkC9bBvBk19HXkjRhFu2aBhx
aetjjEKg0cq2wZoXucNjb/hS3N1oAqV9Y2dcIi9EuXXSBc9MpU0VDBHaCOtXFUr1BloNdTMAUYWt
pyKKMuVI97vyXS2aj4DbJtDSIMkv80t/I9LNFrVfL7d8MyEPSnzql0R0q1DlO1iEAH9qHxCtdP5W
EpFpfJnQr5XnWhGnfNWdhEjO59VZHFSbKCl/W9Dtsg0SchffYJwvHDveGJy3uH5e7gWS+HpYp1Xt
aybn/GqmQbHS9DlztXYDPCFBRTd/bVDlER9uxfsu4tePl8Sf/oDce1KEmKTDqt8dJ7MGPHpACj7h
CmMkLCtpKeJXvG6KOWxErJdzKHblsIIjf1pqc1XZXv9iBvPSLpqHvxsoz4cqQ8+4dLNCuWlsocKs
kXytxlOHleUf/D5epGowZvCdtHhm1n62Sp2UB1Ow8F8BbAk/dvlgV8FLlGEC6z9hK6756Q5fBlIK
HDg7J0pacAR+xqTfDTQ17pxJCeS3HDPOCPWtTioKscdAc2Lu5GrJUiT0w3PmAMDqMEH9/fiHFMpJ
Uh8uybYnxUePDWudIQHfGUQ0tj7LQcUXAqCztIAY7DhGqKw7Fq6bveRhuQNo/cGGf14r/G+ZFswd
pHC6r5gH0H2QjPW1qUV9MI+H6lucIDTf5AR5iT2/huVUvEzNZLsRCSqa+fkBJmGaCX2WEowrpKyb
43jzPr86OkaL6DPjZJAkBhzidUELzXt3/PexX9acPUlLkyCZXWPun0f9n4RfhCnZPqs4raf6/OFy
mfI4/y6u8Flbsj5ftnR089ZA969WrHmL/9PgFTpekYz1zOtUClrsVNf/B4Z74z5UirpXHhz2/8oD
SAMVM+1ZP/8OK5sF3pWfLXXHAsEAb03cIte8800EqoswUKyP/Bm1OyV8dUEc+aeNjquJnYJDNVoW
as5gtLHeW4zJfeT7dVOJd3Mh+qHY8iwcpR31beDi1uzFhO26c+IbcKFCQfzkdsXlcZYTgW9g1lSU
CZ2DttYjtkUrOSrLQHJuocccaVcPDJT/51iJvl8tNrHYBgzHwLYedo8jBkiuboSEsIJiFywAoFc3
mK9Fd56Pv6iwY+5QWHiud75+Wa1pLMSQ3EwRPr7VwLZVWHjcRMGvonoI9Y6g+THYo3JZp0iqbB5g
xcRnKQ7Al2CL5OV67rihmDjX0OuCjyrphl1OCInsH65fz2lStle2iadQun9B9649yhr4ODR27lqb
sed5Imlu/wM6CVPAcvjV0q0Pbxl3dYGUT1NXKYjsl/1IvP56rlON5sFejTttK1XaW8C7ZfW7f9f8
OB80AWhedqec9vyDKxiI4nlat6bUaNx2Z6j1sLMu/uv8YonrgzfruwYuu6gftJJx47IIkWU1mbuJ
tziXavYeg46XCCh0tq8ww48DXiXzRlQaHLpQEGmU9ohyWAM4UEDR3o8bpvpRLuE33/f9sfH3y3XW
4F4vN5gTtmo37fQqXvFndRp6VqVRApQFPy9Mk4IKaDd6EHrTt5Yl+WIrFMSjLXunupK9FK0dl1UQ
mObuO2uiOQLIEm8tOJFv3eiKDS0uPO8UL8nNKbm8OorA+SAXKcMiZlAOyzHjkFatBf9Fbw8qtM4u
D5fzcXPVYXfZGuipzGhD05awVfTIDN7CaQggy8VUtQDSaqV8+yCI7ZL316ME5Vxp53mTQir3Mlta
GS0m4gpe7UXzYPeQQhi8Vn3LDIMfFn5hlmFL9X8gwshVTpkh9G5wbie26W7uSwHs2RnAXTMrYnyU
SD2V8aJpweH/ugWHPQ6nTSqcHeX5DwT7uk1fN7DfNlEWHYFp6gp8vqVHC1LIjkOOBSTLiU82Vsyi
BtMBYxTh/B8TvNG1UDS6fmJIFEU8ZooC/de9gxKWDFccvhxfoG0rjZy978j4D6vk7hvAQkyiMntW
mYq5dBZEMEzDpF/CGIgfAy17x7VY8fTHbVpXqCOKidfoshbH1VyNgi9DUvU+Z1BOFibiVDZ7WjMY
bn3upxrh39yqRweMG2RzmIXQkCcvQfFplEEkxFKdBN81nZ8u2TmvZKOTUIVjmUVP0mcZuzqogky6
8rvGuq/u74WnZgRZE1LJwtoeUPhh70JiNHKlgjbsk1lVJ+ivRjqJO8ScUvDZPHm1X8hlsRXoCSpo
K8Ifj3D1Oz3dD8hEzpUJYfjorLzk0NHjQEnUarFJxRCqRyY4KoPyX53JIODv18WgJIWlQc55YKfV
yGHIqazIXWl9pf6OOZG+gtEa3MVCyLw01uorVoP1BjiJKt+Urct7uGtCZTuplwhuLcZooBdY8TZ5
SA+TkSgn9fGhQKsTL5q8tiDjoMzo+qkBNqwyByV7rmrhE8WRsrhCG0FbecwV3b9BPrJPspx/JSXx
QBFIitj5BLEFeWahqdpTMMmZRIC/4cZmS9sv6v4YEpliF9/XhJgt0MvVfais9am1+/lW2TCos1OY
jvcYGMA4fJgEWb096HBIR+b2d+NYAhfEAFgqmQpa1Dd9A2zdaSjqUIOHGt3Bymrwa+AeqXBsZSuc
5QC4PP4XXcGsMTbw6YE87T8jcocp8IE6NRAYa7+vdeOwhzjReFzLCP+LgdK+AeY3l71fpvga71yE
aKyQczB9ELC2Q3z82CaV8vsqOTPcdhSRXkQwXIU68/DKbN32WUPpQFLu4hQ4FrW+IIcibBng9GeI
lg/urX/DG8U6Tmf+jvWqm9YQrNI0z9fbGJK6Plc+ziR3RTHn1QyRWdrQVlYuxEUlUJGvQpVyBgBs
qEJKIROrUpbvMVrQbYwrITTUeUR7ri6qDCTfEz/K+TRk4Qy786SWP0DO5bZkFN0ytDL6EkVbzG3C
URLUW39PFoE8iqdOmqyy9JJRYi2gp5KRnqrQgmDA6ioWyuMfUJ8878WuyOCI9s3s5kTZhcYeSi4H
XS+998eWZ0wHVdwjKf5+iqy5iy+Xw47hJG/D0rwbJiD5sTNTs2Awf9ZpUcaZ+IySBXtu7DHNgQ58
6tFDe4u4KCYxQQXmOUd0GeGezQv6K2LvI8e26KwXkqCj9FRHK5FemyuDRkK4PX3apeTpqE0CJY5q
2Tsl904SJ3XWmsAkDupW05Kh3OlNAOoaQon6rlVYhhew+RST5BimbBi6f/EM+vqTdUQUr2LcrZed
0wuuH2IfKAwCXOY42QRe2bpaRlVmMqOvRL17CAtiE5kTb1RgnK8+jwwJvnsbU7NNaLXRzJ+Vviqj
kBWOLhdyz/+YAmUjyYKoflnjoSkGIyKQdC6yjfxgaM164iXU3ZRAUU1eskuWgBXMKp+NzmWQ9LW/
rr/QWQwwiZ9JNXH/3Nryzea8o6Gbz68MSwf/sltoQ640AcdgxaDIPlpkQgPXiLZpiGOKZufYQ8L4
Tx29z/tJNpOXEM/VTRERbAm7NihZ3A5D4M111ESWNFlwFH5vqHYnDALq48u4XsP/4t0KXBvQIGVZ
AJ7hor7/zDKyTfyz1JB8Bz//07kRxQQzsGEgRhe44pGBqGePRRoyox2FT8b/YLhtcNEa48bKzlZW
toO6fMmv0PBTrhZPZc8sVy3pC924p/qqFaneOX9Ij8QFv1aS8QNwH05AaAmnaOzcubTGJb327Ndp
s0T6rPLFvIh5Bx//5Evz7MMpkakySc/wrPbI1cfdcQmNuw26vuUwyxP8xilAY0Nijt0c/Ssi0Mvs
NBn5bbuTjmkc92uUvrpODWxRNugRI9U1Ym9kyWmmtS+VKlBkCixW/aSm1rEA4+TK+GTdB+prgVo+
GZUZX7VLK5mYGRr/7kBqbl0xPc6TTYagKM/TV/NNqfRUG/devMKnbqhRVILsRdzhUZpsfOhE9m98
yv5K/oGJSwOEUVKhbI2wFsnatt2OcJ5PIYEaX2vyjWqX4BloYBAPxuPFlODharvi5Cul1RWdng3e
NUKZ73FU3+MBKrJ2fPHzlL2M9m52J2VJRXOoa9FuA8WkPYHuEYGLsxvw/UZdnbHgGseTOl5hHDtV
KAJ/eWhwaZk2IvO5Cd1nFz0NKCAnQiMcMEPFXqh/p5B07Lmx1Wz4jXBBvte68axhXYlancpbISuC
v0wMsbx5XkxziNwjnPOL074Q4aRCIxUVIppNKmiOa5iNXEsGqLsObkoQqX/WaXA3N4WASeqh4lAd
Rq+9FeE/li8UWqKqGPo0t1ewfxtBUtI/4MHJiFc9jMlmCqK1LRR5M1YA4zOZrB1dBHwuJgPV+pro
IS3gfpdeQPmfgwJBEC8KdLlxOFKpJHagHL1+DVNPRWE0uiSftcjo33Ui8hs6OmuMsP7v/B3UhmiM
TczdPWWR2Ad4H8qCRuEIGHuuAwn6U3YCAUeukmWook1+rRlgJWGD+53DkIAQDP5MfkQTRFSX+OIp
wy9LGjCBQyRjQiOS8sJxCIShlwGbcwVtbFfCvHn3StpBHMNuz+XZDlR80xo0AduAmJorcGsjj6F3
wQYFNluW1lXfHIoDS4BkthcwKd6IgJSKL8zQOianJN/p5bINcX6w+beuDMtbeBl+V41F2BUeNzjq
CO9AxkeaDTszmRoopfP5LW/7DBnQ4lKS1RiE14blGIZEyVh2107ALC/W2Z5a33XH9uXPhzoHB7I+
3Rn5z1hvuDPQ83sH7hksme1WoL6wBUEj+tPTj5UYGqB5c0INDA5XgUsn2vtWzMjNxpzc6yL3Tdzc
MLXy/7voabqUEeOTp9HSQH0grU6INZHz1zaTX3Dh/sZb8dRIgER5NmIanyH6v5FDiBbY6Ru3O0OD
TFknFDXXyfYvhYS0QWBhHMIBDOLWU/2ZnppEZJJm5zxM1HSwe03+uskWND9+AELmRIJskZkoWKv8
p7+y5lmqmRUSGOOoJuLmK7vgDkK7ACeHLXJI8pw+EdGMaB1eVlxYOQExDZMQghPk5ymaOSuhulKs
cO7UcCaojyvMGvo+pAcVGvJXXw/IjiesBjd9nEaCQNJg7U9b1inzQIif5/lUQ6hW5cYlAA7Ktp7p
XNwkF/tAN1ZX6KfL69nHDyGzJ4HLc2QVT/mtD4GI/H79L5cry7E1hnYVLSMCMwLLJA9Y5rKae9oP
SPSKi5ZxIKPHETbOpJnhuEa3/quaC4gHyGdoZ4h6IBqjFt6ThWMbknbSxet0Tcbb4TgqjwKDrWR2
K1ACR5b1/N3R6J7QIbvcT7p1aqatpXeBz945YzpUvzHHUTPV6mxYaNvOb2RdQzcypTFDWwUQ8q3c
jP7q+YwbZGEcqOB5L0CWiYX8caHO8OKRMsLfuKAhMgib8tyD1FcU5bIt+A/Thdd5paeDtsppW+IF
VdcsWfdKVq0ALYILoe0CuDKfGULrWRUgeVqjGxViMkKqwFUToL3LvBbbFfkqfe7rYarp6uJ8ce9q
Lh3SVtGpume/kYfcaWn01WOIcFOK3bOl0F0Ioic/q/qM8L3gZmytD9eCYy70yGXlHZaqRquEUXUH
ZWNc6OoVB2EyeuyvddkmWFS13FWkF7RoTpqgkFOxLC7BS03DGzc7898Fe7CsaI0e/XM0AiF9W6xf
2WagKmWLVCkp0GKIGDNatUL0AMmcUk8ydxsjOWR7CFAqVWtxSDsab5PMgjRXMkMMeE3isf4tFA9R
7O2xCpQmAEszHzbS7wH0kG5zRwnwzPvzVO1zNruoAI6GstJ1hpBGIwvcf7HKzdWdSKwRAj65GjNO
1bGaszY0SjUwd8t3nbmafKR2LIbs9k/DQsPHu7hzFt/0b5Dr4PpbRjTDs9qWlTOnPz6yDi9MVcoN
TUcyOeJ1+oSLZFJ+RcUoacFx8uk6xNB0arvDLXBvbffBKA9t1b90Dv7PgFYgUu2g/p/h8zIVPuIE
OS857F12YbXviQ9broR12Y68LN7XjeNqQBWFmySPARngGzMQhkG3gGV5PRxVBhcvGVen3uPuHTK7
evsL6mSzHxpDZmd+2yoj4Yk7GmShM75mzSz6YjBjN0a4bxZ8v4Wl6AbI48o7frrCiJwFD4LevQ4w
2zoKDfxIV/eaXLi0BjePGQiGsDZHj/F+k6Igp02XQDSFBDFJaK+25KFWSILro7XxS2NbwZOWKNW7
ItxlRWnNypQwsF5YxbpnAGIjqAUJgy9fficuTpJoLV1sR7BomhmKYncmAoV9OSulT8F0e5UxocsC
/o/EKRYzrwHokUhWLVqT3n981c+XYUAOnU3blqRPutRuLy7VGSbI/G7N4/EgQd8+1g7X6LmQYJ5H
t3pvYipYKnmwEH6apBIZR/sbJPyMjfoNNrpGAzGqwzhSFx8VpIS1qEJzVmSqyWYUq2Sml93r68At
XGJ5owTJZqDyFuAPRVeX4D90aBoRae5iWmTU9E8GSrGYVhF9o7RGISMrbmJZwW6QavMtwF2xDw2l
eNuQN20gzEcRltsqUWFKrD3aMLY74cg6Jx9OaYVnkjEiG7k2TbxCahxxYEcTOcQ7Ad5nefFxqm04
9gHUY94dLMwFnSB/JTLGsmu/5WfILQ9WIPMdj5jyGMNTG++/rpL4WEZR7oPcSXDxrjPdOWKmueqf
GLcF/0ZtWoBX+mu8L5VhwCTiRljzm01f+4YhUdxs5/g4aZ+oLVEpYJKT59i7KncRIcfqkvdpeZVL
RrFWWyodxh19UZ3wv7ndP1VrLBOcv80UUXul+bmZFjCuDpfBWq3pqSI7wHY/Nerc5tkbDZusnde8
oSV32HR262kv+gqlouYUCewlzfEElwNKVtkCp7W7kYnIQMW9upJE6MPKiN95B633aBgmlId4qYCY
tE3BL2K72q/x65TbYSVooZDhz86xwKk+dJajfjrOT/if60QKGD02SByx5g8RpTwEQDOgDiV0kYPq
87pJUA+zQSz7247gPs5qS320eQamlv/VYbNxt9PQu7ZLXAVgw+9+ezkciEAm18p5V+gJs9/o9n0D
DJ6QHDSHENgpDobY3Nb5kCz289yspKEko/zXbELpWRVOAtrv2aUncM7dzWxANnemzU/UnghdvgFX
wEeGRwmr7AIzgTpHsKD0tKFOz6aLn1QmpoHuxJhn8ibrVHDvDWpN+PM5viryu8eEAQI5hgNpVm+O
E2fEcTEGJlVsxZ3n5ncCYqzGkuqWGKe6y/o7WooRBszaA7h3eQVc9QTAdZuoxeMmQNOSvNWB68ak
CYp9Qi63OYW1V9iL/JRuK3CrcHcl9yfo+3pgebWyeMZft5gnSO9sXEPEFqOMbF7qZgh2mOncvdfl
ylK7F672RBDUK+aBKLRsxqjl3QLuoihnMP8YcNvPNM2B1/E1wWO3s3dqr+uIrP/fLrzWEi3W82vQ
1IidwiMzxdcXXxsfi4LNoV9jqYtEkv3oMXnvZz8Y8JpRs/URtd0ZFSlNLiyQ9wM514f86lSX8iIe
pKnXaXEESbw1Ik6pmc/sADCOwTh5Jq7m9xog+pq4qVm/9i44GGo4zHmtsXAlZOSropu+P2vq+FfQ
nPqw3VhVP9a9rfewDDU7HeQHz45ZsT45eb5NfepS2kY/Fggqr0ifTProjpbJUkCFPc45tV8z03Zt
zVX212BwR4nct2eGFj3lCbHDnosASmEoGWCrZ8qt8s2dU+kcTaokDNXJYxGGkFVw1EbtBDKB4FqX
y6RpN7Wgs4+BQ6RAmEeiQcbBta7HgHJACMvJW4dhUq60OKq67JZSweuyOdM+rumAtUJrwC5PwjPP
bImxboBJoLjHUyBMIudwvLRvG1cRSo92wYzHBKVLtd8W4Smv5K/UumeQKx8C4LeSIgK1Ds3cafrZ
Gw19qgGBTRfPmK1p/OH6L515SU0j4aZP8A61yIthJg08nOj8r4lU1CCSZVT8Q0uoWe7fY64E7ee1
rXulLAaVhLcHXpmt6q97AHSv5GVmeyEtZWMIHKmXy015wxcAIZWtHw9gzQc6zBup9TlBSNW9fLPg
WeOtU60G5r0rOTzbQKLEFV2IkuJTpi79hqLy6GElZbM3yMucbfCtOjWEMmxjKymViANxnOdJYPjE
wKT/Idrr/sR+/U69tSvndS75b2shSB5Jh5HhdVFTcsBnd6JNRxRVcuXs+8E1Z5rxZ21NCyMspLvy
Y2nFFcXKgjMNbgIiuAD6aKB8bNwxOtMtAzOihn3fW6kzp7u8wio5vp8/7vzf/6MNSSSkKOJ2+KDJ
C3CU7CFh9qPlnrcJpU7Qn2F4Bhk+aZBgnFhTtozUvJFHjV66NCixYiYWeOHV6bN9V6PbD2BlotFj
MO+hwgdMDcqn97YzMxu2q+dPCRBb0SdP7B2aifjeNniaTSNZSC1MZWUwii/fP8Y6/IUFtcON6n0J
6BtWMYvEqq/z6eR5Oy5sIFsIQ7nwmvfDsFgP+aCvhveDbXFY8YyXIif4ZJ8K3zt8vvlLdzFLrn7y
ZhSMhT5aEKhN/7SAgTUbgiKiugrVsqURWL0Hi6ooynY7gxgdB3jJ9Imlfq1eVx9Ujy6XF7OQ4Ywr
zBke9DKAKfKWVitITjVPUm0OleuUkMsNuuGeU5wXJr8qng4um8YqMu3yDdfrPRjFdXuK8YwUS0th
DbieJFdoIVIbORk0qJWwVlHFsh45Jv0kEnl03mqfB0yHZjV06y58j02rWisfm/+OG0t+meSPak15
hH9TpWLTTN6wq6uQKrswOhOyDg6MEtlEQgmAxAB22OtrgTr131vssOdDTO2g5FyxehPtwbhOzWta
+eTuplrEo/qw5uvVzWkwKX5KlgADmnuyERPL9iSvE2kVsAUk3WFG4axaNtWbkI5/ZQf12UG6uGgo
AnyzM1VO0FIjNoc3+4yEm7PxU14zzkNp2aSQ/L1tG1BFbFlFhPt1hk3hyJzI7md4aW6JN5G4oeyM
0ofwEIYT4cI3bdjF/g7UrQN10/8j44qYFZPAHbVjQG4N5VElwdQIp+BnAl3yFqUnBNnn1MvgE+xv
vmx1FSdR+T0LQgaM8opN+hUrge3jDTGBhtQ6BKq3QSSs/+quDMGM5nekioidwCVLkIjzXn26CKVu
mDzpLuMzGpy+k+jhDXLqbB/iBF3YuPoRFBlz0F9ycitE9wmyWEsl6tpalPhR/cRruCtv39kry4PD
pta8LMk3tv5q5IJ9Wbiyx0lVOmtlAHrCdsOsvFXJDU/wNTGSHRgkHmfreTQ+qdWVsRQLbMqFgWvC
CCflPeSQSgXQTYIrDqZRka/jayWFd/WWvB0YtZwgMMqBPmWe2J5rElRi2sVt1JZAA5JNUviZ2M4/
0z9nX7d0BC7JcyfnwsSrVECdVSUhUAcS97ZvGyRTOK8PeMdN8gGSe680moJvVg2ZQNSvUu7GHORO
TvIxZqzb9DxAn8NHIJASlh2n4zZelM3i+bzfkR9gKM6rn5KXPl+j9VKAbB4o0lWeYbxEUidElOkD
PyTj/SQ779xydUZw5EEwoK+U9hJ55a+e9TM6/ajXFa0pYXw9mxV7QIab0Okjf6OBcagV02kIrF5M
Irvy12zRE5NtU1xI5znep3IzOzfDOT5EivjtcQTo+0sIhOSskzVhmeEZTIV8wu76ivCQVUvHKC7P
sSMQ/mHmuu0ru8JdCrx/oT6pjuau1mqXU9ukna799f11x+6I7yrapMYvAp+j4k6ZMyx/nDuUrZB/
Jyj8n0asLVukx6G31INmmkaa0DFOGgNDqVBSgOMRr1ETs6SDWWgjIMCI4dYbjW8vfbKZICVyhbKx
hpdPqhEJBSC1Ku1XNhrLgJQ5I5NZ0uotpEB4XOUg3hPOAx9ODs9dvMC6091oWjXtB3FhSjNLjvVy
y0+xvBqeGesdkc1QtKqbmI2QBXoCK+XKa1FnEbO3cIxetW5Zlf1hSsf1dmW5+N2zofhY+vbcVNJI
daAqcwAebuEuoZHYOCNE6R9ewqv/02e/M7w7lrQ+Zrm8mDRkAiGHl6TkDL+RcFOoo9yFn758fJiZ
c0KWHVeITZbd/MWwvdfienL7QvICQwPsl/AleJ8PEyQFzNstV/FOsBKjiE1YOlcju1RO8xY2Ku4P
BrZ0If0XePxrr5oKp0Mm8+5O/dwwGZ//TBL+30s/IPs/5kfzQ0SKD4wjvsSTa9//wSLUn1IHI+vA
dua2glocXWtoCCzq/1OpWS6wecWWp9YAKERqzHRF+bvhbLpDHGdqO/9gPy3KjGFsxgQNBmwKI8He
cYm59gWtOdux0noS1n7ZOOCO1VIRT81Flk0t4QQuISb4IvIJTTXMfd1tGwJwmBMtKqQpWRI6vdwv
694qpLwm13kUMIUKxfyod1zV+1LPHOB32eCC8g1sF/odETSSp9jacR3T42BQBX6OOqJxsqssNydB
Mz3P14wJ1y7pCFpichITkHDfR1nsxBtiw/CeU/7Do9UFezL8oKJeig5Abpa4Tgddl3SKvRHMF/ES
FvUhT01vqlAfnnGGOyC1mrZQtA3Y7Cki+qrMACJFMSwf4VMop+SI9kDwJjifTrUuZlOERIavZ9hw
PYq6RrjtaXP92j4cV/5SKUh2XI+CFXW6UAuHBS5eiYbspyBFXU18ZOvt4usdECwCJa/OTySKGCaP
cbMkoXbu585IQy4oBRTJiUbdDwv9Hm2G0WZMg3ey4sisy+TioFcKtRTho4BedXc3963uRdXsPt48
9wBp2mvnf7Yk0MXbRdSvCCcMftxBCk6QUr6nchrR3I0+MnwQ8vgPTZC4iMGyu+DNMtTqVbUYL0bk
DB4ior4fCZgfgGQvZ55MauoTH+rOMcY++k+7AlNNXWC6lwrpz2PWGtcYFExNzKHizmtrTgkaOwn+
GWSTtL7yFcUnrh8qgp0sT8uO+GTmUXTfcw6tiBp6unehsdj9fb0AJsLbpRKNB9JYMHsKhPVX/jzQ
aT9VBP7u71AT33HW6NJWfsYQmHKA9E7jImsV1LMUysh6XcBU5HoPZXr7yT0SyuH3++ddFrcZ+Ttw
nuMcl/XHArL7x9Piwh2kW0xpr0wt6PRw0b2S258EFhE7auVtEnGYqIhrZTFos3VJJHEdfrglMh2b
7GLxrnwU+W3NMuOGt26B19pk1AMyTmrMxjL+/1lgB4Ku7AgxKEvwFFeR144CVjwt8aFw5QXFDthH
wWOndk2aHR6JWyOdX/sJU6+jPZD0Rfgfg0hKcqAaWS+NMSMOpdWVWN7b0Z0oOzjO27mHqFSfZKwQ
TQVuB7JY5WMQLPHNVj6NBnXPJTnuWYRk5KazlF1EOetNEi9QHBButlXVCzp74KY2wBFbnoSHTbyL
HnRjxXzFZipjuhAkqTKz66PCrBDb9iF3S02GJgXVZfD7RRH6WA0xGExR3nWvXalJNUbW5Li3ciIc
Z2G8WRz0DSNVXYsdTiI51DWAD+UbHd1kt3eBclMX3NrnM9aNCModt7HRuQWJwZUbr5+xOPd3zoLm
VBjLrUeIgtoJ0HNXirnwtbYPK0y1MblQbFAWkPcIKeUHYI8GeRg2P2IifuFLWfUb/YMH9im1Gg7i
w19+j3YYovissEucORXtv+1h95eksi4gS7jy0m06v22j8Vk4Fo5rn4+pwSK6Zu+ioB1wNX7896M6
nmXIeXnxfuQdYb3xCUQYJh6cBfVFh57kRQhgIMGNWf911vtMgkByE3m//xgU7r2ZhP0ZGGQJivsQ
t7rpmX7xUw/qYLwVFSCwj7jHvnOlpph1zj0FuG06bG1WJ716SbQo7k9eLYP8vSt0gXRlaD1PTH86
qnkykPn2YTT6nbQcFEkgWNq8nJuh1yYZ2IRFTK5PzEYPQ6CIE/E44t/RuiavBOwiJaDqLl8Metf8
fdJzA9oje2hoL1EsMuXVQvnGA0PNJQ6BMzzqf0NJ8B4gukUrLLwzqHkwED9E4QRCCVzuQs+T3Khc
EODbX9e7A0lx8v0ZhCeoa+nqWOS2OzGYOwUzvufVFC09X3Esf1fFnju73Qz88KhkxDPE/J05lP8N
FTYtptUaf4C/aOmDVf7pTVp1mxpVLlbviLps2W0cqWBMfHBpV1xpCBkX0QRdFI2RpQ9pEoZMUSx6
8aDoFbfG0ZlPdCCdEqvrYtVsLM4kj/9etQXxpeKJTR+jfqqjRDW4uL46gigFMuZDLqxeAfxgUi2D
1TgHu+6verQ+lXqQhYQ6ySDrb3k0VNThSoJWee34UnUzbvxQGv50IvQGQBmaj23yv5Q1EdmLX5wm
CfkcDukqg/hZUf7SDS58q8mh4b63gYapX4cCa/7kcbU1bQFj/4sK+pgId0GuT62s94m0PjIKLcP6
aavlV7pDhT8Wos/boA0rN/qDESKtPIzLpG23rDBZbrfpQ27PrBNLMlAUCHjlB5zjaw1UMj7qeok9
JBGgrIFrbwK0zRXcPlBVRPC702wd8Iw6YhyARaIXmoPfnDNE714u/ttE1gtr60hXcZXSkrjiAub8
1jnEHpkz8lHb5SccrR9OhbVFFRQHOY68uqICzikK6DL5sk19YB0/ODY5QuzsMgnVQvHGpl21KXkO
kUJin8ou6yqcojysr6IAPt7zo7mc6bTzs/M+lzEAFNqGLpHbNU3wfD6+EmagwAQRt4rRKB1Pfcjd
6socqBlAQUkGqWQMArshk5pC3zyzmTKJWVxfIzq1cSAlnnOcJjvLZ4eFo9Flgnf29amETNg1sPa2
oRZwNVb8guZuQWLTN0MSC5BN5fjtj7JbJJIppKgKam6+Hknk5HwY/0WYloH1SGD+OdnJHQR3vFQL
I0M0QiLFmhmZCyZrRNJJlja+I2KyIUFOXbbcXfvpX1js85LQlZ+negnwtYbzYtlV0bbg/hYgI95U
xvw6cq+syZ7fl68EPUqPzeXAd0I+St/GXlQf+8B+bixX8zTw0Zq+3E2r4AIYBLKuiLyi9BlrTRQT
kYgUxulQdx7MCAlqCvE08rznM3xa+U7wRmtH7FIl8XS5QkmXMjF8B/RIyG88zECeM9Sh1N2Z5B4G
brTMb32yIIfvXs2x5z+qKNSsuWFnR3Zsar2v0pUL5MsvvFNwodp2fCrENIvBYCvfNg8IaylBxTgh
BXVmDsq0LeMRO9MFkoNMgNNuUX4SQGFXDn4agnMJJV5fVaCovJvEcf7u5I8fFvlTZNlk3FeoXBeO
qLiShu9QlB7ce2ukExdh/93K8/gWS1IBP1WJceYVTieEMrShPpOk8cNoOfWvkYdodxhDsDkzsK67
l4Z+dYByX2u7uaTW7c8LtEnxB91YX273NNTzT9G3g9BmUiW9HHn/1kSOVHL6mIJaAYuQW4UfwG16
2QhYFc1CaEEzIlZNi2MkY9w0J7fBHd1wOi8YuS6qUMiJ+EN7HbRAlGoYZqG1c/5cDbuzr0927UVt
y8ihX0udyGiatAE6C6iLw2ISMHkoziiY+wagZknl/Re3cvTFYa9neXaHR7kiapXNhjPnDc0R9IJH
r4i7UCH1Q1f4VAjJLywEtwqQsL/EE7UPusP87oBMQhzOdUxDpQp3PAAfoQo1fGQ0tf6+MlbrJ1Sw
cAOOy8UHPfhJIQhF7tW0aIhRgdlOxzdKYHrVNH5ee102CN0dMFtqasqpYHFuz2m6yTYrhT2bJDcR
MaSe6jiCoHwPIYrCpGfSxZcExsOTKvpXnAjaYhkY5hK+Re+FPwMDmFl+qozwYF2USlpOboawXisX
dcv1N1JB6SkSE3Lbq9VC+xGrJx3utfB73nxen852IN0iKwZKLntFBuKC7UNP8LtKKlyNzbFUDxh4
6BipN8Tf5DT0exlRMpdq4Zk7fKNGG+3e8o7w3IcVj8vdpw4g4fMU5ZO7YbaWtJDW9JFsm007SoVb
Lr8dQupAnMRWCyNSCWHtvyo1kF47Tyad1r80xMqKU04RIDhGk/yrQn0elAoGEVfG/Ic5WIY6G5dh
HS/M9cRyKjkDL9Ot7HyK1txkwvZG0MUoISfRbzq2cWMlndndWWRSUALgdWuA1YO4REcXIDgrEuzi
df3s05M5wMenBRkBrYl4Z5duBpD0pc+220Wm14dlZWuZRJArkCpnZSIASyz3xEi5wArg0ES2oZgY
MJpfL2o5ANhTG2dlFPmkxy7RkqVqqmVYZ+THDqEFLpX2/A0nyrJupFFBJdfHX8Kx6HvXmWR2M/i8
obYVTJLpj/uyJuqNqkQ6j2/Q6PK41H5Z7L1pdW64fpR+oHwRJ+G+XnSEHYWq1uQHk+2QdZkRnaSi
p19PD+t3Owmst+hWLbfdXt1RajvyzLhU0JnUaSpFnuTwNj4XAOhJyH9AHIs4VxvoG6lLDfHKWuOX
RqtLQtK1mtOvRn2K7IlzMppjtmE60Bd6TGvwAeKjGRb6dLImsTu7LWR9B9zwqhD4PWFSttxl0nIx
IzawH4zOJPe3N5KhluWYFKQUNrs6uSScFqRo5o86CV3H4HU21rZpAAOnTxgXzgnbAbMUBLQYdFbv
aqkg1UFIDeqvReP5s73w1gDmeKXu5bMdP83a+xhHPJI8xhdoC0ErooOP3bODg+sOb2xuPi3SOywR
tmY9jqRbPf0y1NCnoWuVCuf4OWW/yAMCfQzqjalK58iVmt04XtUWjmJOmcfzecLq/uG77H5Tg1gJ
zp2Y9923uL7P5WylpYDVZazx/yZfEIFHO5uIwf8FOxEKEg79QTNlWs3kRA0n1zvOlleMyL2HfCLD
RXhozWYJiJKOuaj8PizHLYwGYCGFsitCaSIpUtWrcPmovbP59+qDeniS33hp9jINC9spEliL3eVA
ucGXMBJCe3+23zwr1EqfeJ/i0Vhc6FsG0cxqKYhizXPz/wwjtYdETtz0zyaaZuiQpc4W5gla6Oku
iuV+ymbDvfFhXivC2XuTFgMQqcI3AuwvT8da8vnbFLtj3YVp94FAfIfmHaXwtUhno0GkOxVqWSH6
aoxqrdqbf5HQ2qtWBbHCoJ/85JQWrE1J5H0sYBLi4zqYjLUW1uQLnxL3OQ2XHENf9Hz4PSPLFG4G
yh2VyvvsgsibtBcCR/FTBQ7HovDpSav4a2q5B2XYhxf+/Ui9OEmv4v4S7iIuB5sXMqn9i8HeXviT
VDp+xr8WDf1tz/BXWeIIPqu/TCymvfe62sAjnqttprKCcLdIYkwCs2Sl7GcjbSGGFOVPG9LNZc84
1R/Eao0CC8P4UTRD8LtlrNXPtBhZpnwoA9CUSMMK1P+FC2BQ2VyK0AgWNKEATvMZ0Pk7GUmsF9lS
nwl+tT07WTeaXGHi3puoreuCQLY/mQ4HyYD/P40rN7XkNYYz2NjycEVqWK+bwFQHqCWF3SHcZraV
cH/urfo/IXe6qvRgOFF0AobY/eKLClHQCPxqNUbTqAGwUWYoDgse3SYki9D93pxMo30O46ChqgEz
xrr+LT6bhUjuQZ1HfZbwVTVT0wlgYNSxrAt8ml7wkYmMSmZ/69A9m3hWvZnBzT57wheCsfEgkZsA
ASsPgxnA0y5y9o03dTxoF9FU13R3IgE72ntFdXf4kCRMKJuayxpzfpYCFbMcummkrDvou4OtRVCN
YYWCC65rvsj4dtoFLaKYZoqeccAoXRIKfbC34A1rjK9LNu3x0Z1eVsGEOpw96G1rGb56W0wSFxXo
iWyH+xuDh+iIe6r/KmjCb/FuEkkI7QVwa+nDKdsjrvjeDkuMrrizb2T3XIm21zYa/FFEhnrPbqcc
vATtSmfcB9EMmxo3jVttG5VgOyhgsNXKFMhK6tp+mvnqhfAhi4l/v7xHSJVz4qI5T91EsZhSUQ2R
LGS6Y651B2dRa1Tu3dWjZe1lm+l59vtHBfHWUY46xxnHAJ1Ob5OJWscp5OxTd3seXQnHtnDEAwgA
WVPvdnto9P6kmgbcHbezvNSq4cnPh2DNbWfNVrNpIPM5j2CL3QBMGe/bg1jjg5JEqia1t1sX48Qb
v5Xw4OSUdVgUilRlxnaGEACi1jSqlhvLtOX9J3P6XZNBV9rU+86siAV317vlDTgqq9/aH+fkEW/D
yXm5w61a5mGw4EUVyoM0lVvke/lCVw/lurHIxFtmGlyj9ew3S/8vkt2gFM+owQ9r8ldQbQQEzuvu
Oyo9RpkN1C/aI9EMaS8ji0ieoc/5gUmXhI5yHnQ2Dcs/E3IILrloADYdL4oj7IWF6jKEbmmYC29l
Tb76M4pEDHozwr0jsX8ttcxaxKFr9ub98rt2dEhZzmEyqmlIIDp9aNG0JqizN4oexb5ZGkCWCwlS
VPUgHtKA6At8UdQZjCKrvJTvFKqt2Hn914q51561fh4SiXMNwHEXpvso8bzf+3cjOn9JMNVaeXQ8
h2OHhaawUoPjKeh2Hkkwarz4zPOBy2Smijx0V2+kvJD2PTA/MY5EzpU6O8sM3JS3nE7cctg5x31G
sKJ6dOgpo9QeiHCyqLj+ohpLf/ZOVzOVc2Tz7AqOoDB3UT1J8t8z9mJbNK+jOYeufuiYtEUvxumt
c8crmJlFKlHTVRz9DGVFOnOIyVRRvUKqOWte6sivcTFbg8XpMLylRvcPevaaO1w3y8gLCyQ11L4U
D+Rgz10F9D0kHWxQ7N0BtA2sbbF19M7m8I23Fiiz0MvEe9wV2Rot4i42CAXgeYC3DoQis+SozQXt
wttPdEkeJ4X3wyKnHX13FKRAN4j2LIVrJYHrWwzEUEnYzx95A7Y5TeMJP4WyKj4oTaIf3QgX8hQ3
Ih+Xxrx8xoj7X7mIpWqtMuj+6iXzlit1zJOf89/9AhIHJdTlJ8NLvFFBwadRwz7MLtmydO3lvEWd
76tKZ88zJbSkkIwMpQussNOru/l8EQjSODQeYcAoOoPQ9h5uflRwxo42WkyEnuf8DvwYiW3q6WoB
lTMHR64ANTFnaAa5+lxvCL0KbIO2mTDQLgSTDyhwaKGR15FTLZqohX9h6luMyjy1galKC6ywiOcH
76P0BGSwaLwi8SCjLfqQ5O4s+6fShXZUoXftMzZ2sWHzYCvyKR17pR44drwRCyPOHvbSxcD474x9
+STtxTXqo1vMaVL/p5aTaCh6FlPJmc2K9WSCTaT9k6+AFfVNfKTadogw51BKMrdCNnuARxXFdRe+
bPsHjRjvDFaUm7AdaxgSMykhSU4garpdKOyJCtnp1KVgt2I7fFvjphR3+ePOrPm3qW6V1ZKl7DNG
ftNs5t4y6adxgVLkepUq6IEHvwHv4WhmZsQN1vkERxSiJ5VTbIGvtJtNxGnhjN2Axw4myUaPRC/c
BQ8NLc1YoFl0MGl3DeMrdPZ357ubPiFoj/TVeGDq2snupYaPAFPjBHHQBsr+iwM30Ty7zVdssLa6
xi0t2oPVtWJpJL54SbzA1ouw89TejtEx8O9bRjSCG9WVVx7vWcCjTaKV4Pa+8G+T1k8aTec0skwP
G1+Z2xqKp5nz7+9G+2sE94zk2xzQyo9Zwpwn5Oypn9BFy4EtqMGclpWua65fzv7VL9IULBZc/iXx
8EYv9wst4s8OSw0t+S08FGu4vuQCu2qCPXYmTJnAXSoiJzuKrNmQMZ3b8HplCHnEylrIyKYnRYEI
VklLo/+Wyf5MGf1J+i0XP3akfoeHTrw9c3hOYKjsQw87ySzyajryI3dLLfsrjjT8ZbaeLoCcrWxM
C4OKlyqyUcofFC40WfnL2jQDndngcUC3xuF+XbIoj62IeoM2fS2jt9U0fKvaI/dL4RX4SX0rz0e3
7joF3kn0bwCfSxBRhYxIeil6unv83rHmL5Ib4Ak99EdSyQjO7Xu2XNX9NX8OP2X94rL/eDSxWZNP
SER59uwz00PHik0ZBayxTq8rjcCHcdBQZurJyy09CP1ISB7Qy9fqhdvhM9KNvJXmU0CrlhXHqjMH
3rQd47pk/cWyZZ+MMfvovXV07brdH4t1OlF5HFi65uuGLlj1SnDilqiYRV0oxYQyiqNi6OE3GPeD
jG+vRXq6viwxkZpAMsnt1rQnO12+57MOlkyPQ0gkwco0fMM/Xuf1bhhzUSZrsIgvQd3mUUbYSLrS
OamrfgxCYSi6nimAu9jSYzEcvUxTipO7awoBr2MD6tKT/d8Os0WnYPNBIPOqFnLJJeX/C0l1KGNL
ChEXKsJC4zRewxPLmmI0GZBSZ0tPBqWH9+3Fqd3jppA7MFJ8301TaqmHebfXcZRawtIP+DfyEj5e
RSrWdC+7L8ggNihJrTBsEq7sGz452xcmts8jBsdMzLTV9P81g4BN0zK+BgStBnWwK0ck/XNLLwpc
we4XMjlDoUvcy/q6L4owu4iXkDNH5wpYXI2hbohdolL/W2Q1pRfxFW4AGorYjFke5T6eNMa25uKu
6kW6ahKWVcwrGc4LVmg7B8lIQqnkMOCdqjxKp2XddmbK664AiKN8oAuXhB81S4tJQ4SVU6e5IlN7
sqoxyzH445gayxueNev14Amk39oRoiNQnOYwm9T+wCY/RO4LfmxpLsGjdL1vBYlp22QNZ1WDl83v
szP6Bv13AIAPN5nDJa+Ouaw7RffeooWaXycX+FKW1qAa8ieI+yY1p2jU43B4Kks/+66ln4HueKXC
12rn42Wg16rb61cyKV6kxr0FXFDN2OskZFKiEZwAoYC3FylSVSvhSdqN9o70W7FyMHhtQfz3wf1w
jU0YDU2XlqJmXsEafP+sT/zN+VRC6lL6P6ZI6O7NvB/Vgn1yJVGeCNFKi1YWOQS93bPO9GCxabwz
n0KBBVRRvPVb+tpBcpsWFYvB/gCEKzZ69IjhiiH+bsvgjIGVLYuWXWnBjPDCx9Ut19STtOhzIVFM
qUPsco6iDFkY0NdCk5tgCsZ4Q/1N3zVnxkNjnvXB2Far90rF1m1rz9FuOqHwsU/BJAOPF4LUB0U8
ht0votw4cZeAiHrg6X4vnO9bvaM1kSjeTX74dEn5tnIgUuTTs6dF6IXAArftsXFM09H18a03vPTE
PknPaAF550ZjwUu6meXJAGFlbYJO6kORTMbpuS5xVhZQ9uQLdgxHdS0gKEzn5DlZyT7fw3OKgUwV
a4RwdQURb9Nmp/JkwBrkCt28mbqT1uh+o6V5IjOhMYv4e1tWuoLxM+l/nJxdO8/dTqGAmsPGM4UL
474MZp/imfzT6IJvJ2oWhSyB5ugLClGTSfASrf++jkfk91RAMa0WJOsLr3564AdtWewrQuhL+OG8
qs4nDMmABDb7iNdvBFzVxHYrdT8fuLwZ8A3Y3vG1i/DxNbggUNVyRQwPAy/kBZnAYpibW3faPVRH
ZVXDzHegRtVTic9b1r47I5L3o2tbb3pULTYeF/uxRdTedRrBatm1LLdxVcuEMNfJKrZm9ijhFkG2
69AwBz/fe3T8b8Wzxa5I8l6eUwbtod1jDOc3NxJu2rVGBV1iAP/5DD9UV8st5T+CA36Dy2PUns2w
SkM25b/7LzCEjw9O4jeHD+ZxkmvZW3s/F9VwkhJcwHxiQpAhuLnrJO6uQixToelyJW+unvC2qvys
FjFZUMKdzJll7d2SnxDVaqLGyNZTENKbNTOqwvHthPdlN6T60W7mu3FDDAKXXThiV9LX6j0Q9a57
UfRq89F9/HMX45u7Ex7L3DQ4Nsur/7e9KpJcgmWkHsOOZijdCUiW7omtdHzksnEtciCaUFvOcytI
vSpRIDURemxbSoy4EJu+6pHf/vJeWzjDv8ZuKAoze08HzE08V5/fAWE2Txfl5LSCA3EEvHKXk9dQ
ixHrwimcXPdRhHL3xmh2BYYTmH/Mr1q4brYcBHgC3ejx4Ug16OhZSi/vbI1+F+YOW6Q3n/nlKRxy
NtsB0HmlQMqTg0tGIrAKdllCgonJgv7bXLpYGOy0p6rLc5WFS9jHGG0ERdMhguIJXg5uT0xtPUJl
aGenGA5dfvGGR4p9va563NyBgNqlamiqbQbAeSVfP5bS57GLGJDnYAQ/aTEkWK6dEUH2kYDovH0l
GLWTLFP+08BLURtKnYVhK5vc0Xvp8s36+H4KK5oSneoAlVqbLAbgnN/6r1hXYF8w4V0eH1ls48O1
pH9RCmg6FrxOxUVTr5fYGzARWilXjnYS9WDBnL91RxkQ+38WpV183HekNiTCz1rZ40+CAQ1ty5km
Q3U3VdL6r9l3OTi3BZiHTE8u7TeNhd7BTQFn52gqHPnlZfYIa9jGT6N23+UutBKar6saXzF9wSx3
EdJTZKIPo/gJVeHUrwLTYb7EzNyluHpHYb7l8cLGWDWG9RPzV6oBpCmaHta7LlENPpYIjVX+gwHx
6raG+BH1vBGSoO1Vm9vRDS2cp8rMq5vxVeAmW9wdHNY9qpvmgaho3Mqk/J2GeNZjY0C+6raOw4Wo
JTir7xO4q105kFWaZC2UbOokVpzFVKpRUQgdGGu2vtT97gHvoSINebp/vIIXYuZaU2bn0db3M08h
yJAS5a14/hUgS5ClJHOMDjQammucoVZ+UX7h3bpLW/psEfwRzY5cVBepEqZaCHkkRjieaLZM+6VS
M9tEoOOfmlHPSodBo4b9YNH0FpOWYgfkqfywqRhhCeNJDpQaIjIvyQO2su3dYD7AfuB+0w8JyNvV
KOoePv8f28HQJw1n31Uj3mpfxgs4F+PsMugSkoSeLMeqf4SWaZo91HDZumMxuFiBSAk5Z5OOfGQH
oPe0rv9zUKjz3aYC05QzjroBq63LdFC++sadgqZm5MI1MMHp6IA9vReLDrO+gb/R0LQbLSbvSjac
KRGTBJ3ajGSPXXDEblLnV0QhTq5bxrpA9tVmJ/rd0OFnK4R2hl9WXWtAsY2iabdbman8kWrxtzxl
4KKEFKlKDceMFktS700p9XebKNEtkMmtOO9TAULHoyyhjqzZn+1h4vi7mY6oWjKzPgGY8puKSioW
r3Mmaro4t+waLAcRKFGTe05E06sWwF/GdwWefQYXUFYfyUIbrl0JYXpkJ1QWhTFObOJpOBLk0Ysw
nutAALwXgMe5klpaZ1eInNDCl+sF7j1ZBHJPGEncxWzICmRb92SRO0jPNia/+ibKMIXQF1eW3fmC
Z7fmJrKqx47Hst+eZrWcAf16tb9ff7GTZIJT89XPNfE77Z9S7ECwBOBL8JDgAy3sFM1vXc54xG08
Vv6pypfLf08woq1b8PBus7c3c+BF0p+4rbgQ0wLszRP2v+FHJe/uvCgZc9YV35Sy079RRNkuzk6U
FBGLoimwyafglhDlNfMUO3W2Ne+PqQSSg12i1TWLW1B1k4cCttWJxfg7NR2ph8wsKt1p8Ue6tVHp
Mnt1ncNs4v51qs3a/hq2gwJPYV08SNuyaRU543til86wz082TKSI28tx1SqZQK2BjSdHT68JUALw
uYFRfT0yuDmOSeV5T7UnA/tNthqhwnz4I+w79rk+iZSLA/SQuZm913ZlSxLiwkHPXfGHKd180IQ5
xe+Hl+uEFu84c0MFr7IxkHqQxxD1fjOQDNEJEQIXBt38ip0Qrczn1ok+FhcYoX2f9wyj0x/p+Zhz
TaHEcnYyyc5uMBbr9lr9DpULufju9dVGVaAGDS2CdwBqznCRWK+fAwzwPKX8K4ZYHtpzAy0Rb81O
PyKENvCXGpXNxOWHstsrZky4VL1yjMxmr1SXNzE0R4Ah9jB38KhEoxUR1r3Iwj+tnutKX+5R2tbz
EfOJZ8gltI/0DoT+B1NnIdJZ7hdzS006w7b65CEiwzgMZE+fvDcHT5g9iiQ9rWABvCOpj6B09n2V
mR69uY62jA2dlWAjejA6CuES1g2e9itfJgOZQ9Lx6BGS0VM2GdyW5e3ORCAtQW0tt1LzLSlFY207
oj0vBIHW3WAiVBD/Ob6pXcTgwJVQsIhclnRI05OLbfSM2csi684F58tyG27S84B95Gyv/Eb8ua+4
kOV6c3jFdFB8aX50yRd9WDa1fQGSRbNJDN7KC1hyOQ7CnkBedPOXnPPCMWzwqWbXCRB5beDRAZX9
HLp17mPFCUisog2ZgQo/qaXXjOLcaTVgPf9yTQLAyr+BVKb6sQaxYVk6TazFDjupufmfI71G2L0i
xK2oKJVPwNbE4WtGa7SjGGHd4fjO2XpamfANVlsO1+42pYnco04BNYXVI4Cw4m7OuaRpMb4bKyUE
oo3+aVuXXs8sImN8lMBdbZVOioPRi6eQSJmyg2Zcc2W5yuVl/og5OIGJreK3f8ECmVYdm6SYP6J/
296C52h8ehmGm/ZmUtzNicOoH1/AmhwnGbAwsjU+VfHCoz5Aa2S2dj7WU0oxxSSk26oYuTOBFjeX
V1qoi/l000InG5I306au7xihiJ7sVspzeRb7YizfeYBSVXSi5sKuuBnx4btjl7BcgUm6hxv2v91C
HpiUb+yozn6jMcHftota47lkzt2XdxpLKrOoJnfHxNGIBpjJkz07ETmlZET5iHtZ87XDfr3O3O7K
4wbQmKyuSf1H4474LDGX3E7gTkhLD+V7VXvhYbtd2FJ9bTW9eYNTgkGyTmwmN/W7YZxzqmRglTuE
ilQqIvMEjf2/g6foOUmTodX1RHQ4tQEMy6OuDCrbn8NBLJcCx2IUxoWl0/PQTPdeBVmXUxiIIncQ
wmvJJSNzwgDnq+SIiidUefFSOOy27k6GfNsw5E1YhkeCOGvuA5TYBQDSJBB4Rl7zTa6rsOOi9P0H
zVlEq9js5VLnH7ECMxIkHsoW/PvhHPROHmUo926zJhojNSXTK1y8j4zwlOGqGRe13rEBMr+ZpDoZ
VLx9foltoEKDLRKQ2Eeigwa96rWx7U+AxrxyEj3ZWx7AOdEKRlF+aoI7nG5umELLkNu9CA9RBLMB
JTcsb8u/0sxGES4bnefAQ3RlHYzlYOn5luFcbKDrUJIKIPfHG1pFRplTk3ctAtAFa1TzE7I++I9F
IAu+8nz1XQ4fcfcxhEZECkMSOCW9S/b5wUdsFms7z+yeugL6/HiHsD01i8599rVccq+9/ksL+dy8
fTLeNXwZ+Wkx1XAhTUeImjdduwT9z8LloCBSg2M7oT3bsXrC49JgKx6OJI6OdrR/fWDMx4Kv3q0e
BXeEPbiTJtXgaHkcZl8Trlu7OCGLOjYQ81sCmhB+LLKewAJst/R/VHbg+LgT8gfprl7OJmKJ0eAP
Xtf0QkNgAvfSFy5cdgg/MTSbuN7ka3jTf63Eml232BFMDnrSDwkR4USlHCKYQ5wqsv2VRciQ4+IC
VueNZ0fSvcnugv1pzWZJpX09374xogrN+nFIE9FLnL5sPfDboWtPLOI8VN7J3s5vup/AZsQI7cbi
zRh6WVrRvAMY/HB3sbN3cs6q3Px/6G7y2Y3a7GX3xqsl2Nx0icd1PM7uoKp0AOAx4N6W/0cQsU2b
OTZ/E74/b+iMq5Vv0ErhWVrQhel1zF3g8Iz9SXW/8fKF+VaKaVGD99wFs3sadFfJLHmN6RQWY/1D
gCyHKisuvmJJr/q2I6/CBsCHQIhm/OU2FJzWBv6WZC2Ldy296RNIAt35AdClXYhfp/thEVx4PUjZ
rdHUJjYxMy78+xtH1Lz+wTo69sqDKtQkaC0czCxDhD0Ul1dnXZxXsbCdzk/guR6cwmHlbvXXavaf
UCYRNkP9w7KjRYVIk7QbvzBXgiLT8O1qgF5OoA0utXniuFxzVM0bp9ttQcf0xoTM6QTwfV73T3z/
ln4tKKpWDFYw6G1jB/cNbRg07l8NgIeS5RJYRL6+ZV/qVB+BK1R1hXRNy86oHbA6t27hRP9XXy9W
cKV6e/gp1Nu04+7awvxfIbtGS5wghlxR6dqR002+37TVeLfWR7s2srMfXwBU786/86pZ93hQRXpU
jMlHLUab/2ZLSPqKr+QOimrYPhv+ER02CgO1DWMHctoECor2iBgcUJKHO6Y2WFrB3lwuVooaz0oU
frqV1LcxpqAsOwuldf92V5tO8luKTxPt/SUIPrwY03Q+SogVtxfGpma1iwy4Isy5xJH28oHY/d+R
voLZkZq7XZjdzArCHfjq+m0osJtxF0xfeQ+RN0Zv6lgHDEEM2d3qIA2oVM7p3fAQXKwXleLHASHs
SlJvrfmpFy/SucA3seDmcUMwoM2os9XUfnLUtDbiaec/3ri4luEIPkvUgJdWaJrexqSLhwgJTRhq
pLEWUBnQbmK8cbPsV0EJzL2LLXSvq3zuzvpjHKQBVxeF58swxfPzQ7IOaUyl7UbrfJ1bIMngz+wq
S1dwPEk0N06wqRxF1KYD12jHO9PXvWdICi/v1ra51Ly7fyfW6giVJES62VIUD+xafDTKPYsPPOzn
YSLgk3nQkCRCFY2OSV5a256E1W5PfOxJ6WifAnEJNVwtKl3OO4oKydtmYctwT8fLx6SY6dHjAfRV
zj56+St56+wK9w4ikRWiZvo6i/fICCBRQ01aWk1HaWeIa8+3QSHc7jrpBg7yDVaVIiJiX3zDL1uk
lx5yjar6YEKmE8vVtTitsO+qAZMQLKQRdx5xf4CkAamJ+UQyJ2v9zRpF7mcrTLS11BeTgTuNNEDK
/H+y43WyZZrc/2kUHlK2XQEwHQrwpOSoYb6xpDlcxaFtjgO62uzjCkcWvnml+yapFqcZvZ4JzCOO
+AOqslLBdQPsu+JnPCSR2FSgCZEPt9W/d20n8e/zhsiF1G6APGER0PaWGmfZ8kJ0GgadFIoNB+Hm
zqvs8+URC91ejbHn/oj1JBAgwOkcrTJy15Bi3jwqodQOXVDPzq+FjePi09Xhbh0qVddbeW0jME6J
pIlIMbpUCMmhwapJJtmPVZIN49DoGAtAVx88Lbfh3cMlOYzAaVYi3XGomQ+53h3qwf7wVShps0AO
2J1DLdt6WcHZo74MrqLbkPXGARkXEEo3TjVhKIb226fp44MCol/vjv/523GtDzWf4mZZw1/MGU/P
SKfnTlnkYdclm7lVpC6wZe6edAbtqPyNuaWqcjuzBYWIRSQdAEvlt2u2HOWYjkThJgbE+vV0H1DV
czL5SskcT/l3FqQHrpKGBl+2sG0Jt/2IjULyB4JwI/O4cp7cBYUoCSc1kAQFdNK0GMK45uyTNaDw
lXPJ1gOIaXw0ErjtIVbKdyGvOcRsngXaTVVna9w4omfiX5kKr9lkvQ07ieaDENCJhZ9I9tDB53Pd
1yuKmc1eiQOO4F1b3L0cJeMpchLpGDAWYuyXodK17JtODYzMcqOZsAyOeu2S6UpVVpd/nFBQOk8v
GBHm15ih5fnGxxRgSBwcnt9+AngG5H9emq582WYDePdB04x6n+ddBr8RDE6R7NTuRzCBSJE4U2FQ
oo1qiTRuvDFkK0v/DXsh8oGcmFuXV2T+cBvrE1o7YYhE75ISjc9XhCFN5xWl6EOFMK0inNJStzdV
mdWXb3Hm11sW6/aBOs7G1Mw7PhoB8ZK6rLzibJmU2TryEfdhT+un/pMIz3eiq7YJO2bcXVZel/Kg
NMl2w6vDFyPHifchMrwRPx6P8xhkdjiMx5m1PgEyi8imbD8KE73hM/SHLHc8AgVXrz9C30yr6kZH
wWpAIXWkkIfSRG5PaehRRUV4/mooq/NyGzmKbsDL7vv26aTDL0RxVGhMsSVQiR1/Y223LH91oh0Q
+T9s6M1EivFL++mbT3i4HPiCMMIOsKwqga5WszUws+wuPtSRScjJStxz8k4laVB740ula1Khk3CW
tXgTuU5nFoIERyo5fcCjrfh1hlKAJFbIbvDeZFNaHEQw4PWcHantZMZ2a2JWGn85O+DDfbaxw5Dm
Vm1WFUHpkqHeypBnkIL0yUgxqUBsWLfaSrc4q2NW8Z5PBZKPcHduwAaM93myH/YfQyhXW7tYMDLR
T4hXQ+X8+2dMO7270Cs9RMm0YTZQH0R+B46Xzh4CJz7Uy0VN+B0QbJQGwRfTPGAE7zD3blsNHhJ6
NihSLV0O3fhro6BWvU8xT4i8wkNo6mA5cFB8Ep6iaFf7Lf9WiRObNnUgL8NAwP8DW2yuNN8QfR0A
P0LfwP15EZ1alMgQA6RX5v1GTJ0EZQts9IdnRUYxANWmvSbTRHpnwqRCfx4VbLBgnKGHgoy8aPum
RAShwbmi7Kc13MlW/qoWwpmK6ZbMAjyDwUkGbkph8pdGbb3+5eNCDZ3ZZcm9m+3kwt/uEcxoShSL
9eQrt0uUJiA2ZBZouvwq5cS5NOXKjRi8voOty6JezrmNObwGpw6L1wyzKtuAm+leqKz40PgKdaHz
qQi9SH2XCs4aAhmbd3N989B1XAV06cXN3/RGkaV+ZCmpHKXgeMYiv3oXzGjWYl41056M2wDvqncg
uYcFd8DP/7Gxz+MjpFjNhuPlRaTGOBF6sMPyWxL6bhCkLXf9DG52GvSEu3nRE0o6OpnOBEWqatAH
cXTjcD88hQQU5VUthqOstqwsQbrTbcRV/eVwpua1/vJUH3i//xQE1zp37/+UP4EvmZgdHhPMmRLK
fLas+TqHFkqdLlf6khy06Q9vyx8Fz6X1mFvxgCSN+9gnA6USM4MC5qAR+ODrEr2tRfbodW9QNozC
dkjb89MYeFjNji8jMfINNRT6Fv0FXTnCfK9dQ5czqp9JwF726LYB9utGSFD3H3MnG6tOXOwmVtq0
D1LwnwSqr2zF7KgaBUwvZatuLuA7NDv3rpUhblGAP5zKc2LYatkbj3iZVXPfY+kQr+CP+s27bUgD
kk5bWuBZZ2G4ip1zGRM34NlUcVhJwWQCCZEGcuffS7Apl23uxzdoryowUjIZX0v5SvoE2FvJ1QrD
NTRU2sJpSjWs8Y7XiedVVnNO+X+Gl9PqileInK/8+GPMRA96FC9oLXVJwaJ8G9v5dvjHMwbjlZkI
KaMlTYIwuW41vIVYzhbZj6A3YHH07tgAQXamtR/8wdtEKpEckurbh6ShO3sx+IDsN9PVFVhscgKC
S4vNmPF371FBYeqaG0LB77PbV9vgsqZDz02Cgar+TAqtZbP5mOO8vhHsdJI8iyktcaV4pw/Rlt5N
uyKnqCAD+CmLmkQ+vgGHmPw1uPcxEw/O0SdCZ8byXd3hA5a1hCkbH7+IoGPfm5G1wJM+2quzlUgB
WzZra+BfHk5IW27ukJwbPblLCyDEktWmGydlBhrkXTwig+UkKZPmX6yNmV86MFbVnUXn4xyxjpGu
uWqxO4ZYfaw8zsrGeVQ/qjyBbPSdB3zHtjufnPeW0p3a+DLVi/B0fOGqOmXKPOfkfjHmqOwD9n96
SmN9VFu702WnydIbVolxxUQZoMsrXkHYyzNHPtR9CssAc+KnV+FEp7nqdA7O5pQapidqB64xPag9
XhwvEVflfpQ3xKfa/w9LOKiYn4wpLMWycRhWmraR6E515N1B5DrxSJT2tOJ52RCAbE422cUeEZSQ
pzRTkUQ/2dKub7IDOI5osUk7PN9ix/yNNDbNdNX7HyRtDtASePGcB/f0R/HuSM8k8Pkxk1cng/uR
fMdD/kKldNgTq7w9bIXsjTeVDshghJD4bzaL7SZblBgIYDA0ZamexZ62oC1/g8VFk+uLpMWyije5
xMXmG16s8mzjt+H3AueKro88uIr4mHKiUV2Lio5Cq04rdwcqp97dzIGm0twT4+ipCicNdnwDvTP3
C1yiCwf66dSZYwtA3rMi3U/F6pDewowYoYdZPGrlEttd5KCK8P1zxl8HWXujWhPJaHL3OPXLWpOv
xa/axBtxZ3hP5dhd6ANLXRPMjYRfijnFKd8glcceoH1Ge4KDpqnvz1mc1+R5czvP4O1DuYQJdBbH
rrNYXmSINKvK5BQQTEu+Z55ZmHGzX5Kb1b6BwKKOHetn75z1bZfqzJRi9F91vx+6UZ5CBPMgRXmJ
MX0wK10+vIzUv+z6UdI1zAXADHEHXfSn9T5xO8ksh6Ab1VCCmwvhaL7kyUzBzKC0RnN5OYo6rYkv
QYhtZm0Mb5mAiD5KKhuG0Bf+PvtgZ09rBBxfXTblGDKgCSzyVUl+Nw6jkD1RCzQmgzGp+yUg7Ye3
k6E92539fXVAgphAKx9QYf6ZYeWfMdgqj9sKgcafG+5rYJlfcMbMQfosaWUMy/G/oNHDh7WxsfBS
wT0Z19vpKy7QAE24FqDG4topHd9hu3CE8KJwLWXS4zUiBjacKMP7FcJvyfTlbMCZoLE7DCIb34OA
4wVKZqJto4WvES0p9/jkvO1JNjVF6HfCdgCKxbqWb7Gk91eaG+YqaSVc59gpE3wsQ9iLEoshA325
JidiTG/yERfQGWOZlfukick8lj/4e4drIbMFeOBUipsVs+ayFmoohng3dBlhuH9p6Lf6bL/MWtQ8
n6xvePrqz9wgXpE7e96feAD1GQqMNsyQY9pO7aepElCxZk4dxI6r06QHgfNXUter3tNuvTyjUUPE
RLbENpHdrKqOCqV7VXOsxwGcAD6BuT6okH/sGxeuVbLUdb4qWLTzBUltEMwGrPjIBcBOqIed/ye3
2HkxXe9M81UJxe7taPAN1UBaKibO9d5IZElOC/8wExd4J4aJ/+pEexjZ3JicYLFTA59v9bJ4igxV
h4FFQmq9+VDWdoH3V7XSsi+kVzGmacom+R2RvpGr1XgHgc1hNYiXwkBXqewf73MYJdbNV3eLlOmk
JAcbPNwLGMronmjyTqGp1v8rtmnXJAxT4bZ+6fiiIaCWHmU1kT+eL52QvBJDAyqEGDduO+bvg9RA
+K1T7COcrcQdDJBp4DkwumbhJSphAG2fp4+Pw3f8B4QyGV16IFMaRFTiSWcsfjl5Zv9S9ttbztwc
0jUNd1R/miuIwyvADBFKwSAdd/tN5lREOvipci8donB6cq7mbia3JTBDi4brzmtxhnZ0d0n22FWr
paayCj9DBU3vwrm5IcJv1NLs+P3K7zq5/bXdi56Gh6e+KjwawXs0O9aGX2wNvKOmuMA8etagjWIZ
brYlscGkNLzTdZhs7gZ9kyiIs7gKK2lST9LeRCJJzI0Ns2ogy+XZI9nqDkbSTlD4oXkqJJuUgTFc
n35Phk3a2/EPWOL6L92qPzAGzRjzbtr/CcPaplWW8hVG6ufGIJK+UnhSRfCputj8j4ZErE5Yrop8
pD8juyDj5EWgMqaOe7Pkt/kkIzuL0/VhYnf5CFPbG0AlOxsv/X2e25Y973S/70qS3v3pANxE59cC
vRgGKAGKQMXUNMncQMfmmG+TU+14TFbofThLVL7onXHdUyI8cGxmyRUklAqwnkfFHKIyk+8Lrjfa
sMGaCGiQJBnnQaPywQ3k7mS85CKuiGXdZUIgDuV0G1FjAlRBW/cFhyfz97ohKi4Z6PNA9omuiwOY
v76ufqND5aekBHx6+1NcpD/DMpTAE6M4RReLnYtri3Eox5HbMwOt8MimtbynoBdmiyhJO34teQD3
6cHZdWE5EMzHCODC1h3aGT3xNAQQyDxsUgxis9FN2755OZXJuuAt1aUei890SlwEOnfcz3WSnOk6
MhMsH6Q/Us9cuZOoMTaV5PoJwEW+aboRyLqCnPXEKRNe5qPHithQBw0zHb0l8LhD8ceFtrPRj5Oq
sUYX9MKRrQza0X766JrD3JwGOqlcVQQhtOL8iNIavdR4QTznHZESulkJkL/qQF5Ir3Vv7ixbwYyo
Q+0kiasgCHc5TRLPDmuQ7QmSuLR6Djva5YvNpt/wcRPpGGm68cIdBw8n/1R0ea8GXT9gwyRYju+r
O8kN4DSYcA729finnYzgQfrzimxv+Ku5QXEo9vcsof9hAI8HTsEzFuo6/QZMmndU+55mx0pUBcNZ
wsDET5qRw695kn6LuYtZgia6i8ekAIhmYJdZ5/NyBSM1RrkwM6C21GinLrx7TAGLZvp+S52KgZUp
5CDwJq8X/+A4WGzAOwh6XZs7zgTdhD1OvOmJug5OjYLtLRKWzhlM2hbv6uCnwv/gf2+yWUgmVtUi
kcBnHOe3RW2lzDNCSSsnWU5alJrlW36z/DpBMA/tQKYj1FzA5mf8/xxd3lsH5V1d4s3NQjo9kHrJ
NUAo1WaIVhaM7HKcWB1nhxoPy4GyKPQlnoq0u3Q7AmQ9PIjlVHKUHbiBMcHozgNde3uBOyL+tJgQ
zmLpqplQ6p+dTCN5P/ai7VK49n/yci/1G+/J4FnRgMK3S6bhewJ5WbBKmeItby5P7zIhnMGsyiy/
XQ7hklh6o6jVgb0UeiXl0XbSuxZAIOojv/CGgn5u7R0qDa0tOhOGjapa1eIpQi+6+aHck/JaO3L7
u9fwcI1+BBJadqZov2ICq5Nhm+JQHLbrYPZQfcr0mbA/G/HkHV2TQJfMgq9uEmiA4hDQauS0scGK
zQIXfyoo0NBUlJCvaqoy76gzmTPjB/8k8AsMlmvJ5kKlmzSwjFH/v1qnqX7oTh5nVolK1Vlriwsf
HYCRhM8GUMmWyVIWOZMxnqLVguph0h2l+l9ASROfY+Rm9fdqsD/2HDgO8Y/Ik7fjg4LEEKuvBXJr
R8H0eocC0JnB/iXMuYNWm3YPbCEt83qBrF/X2xqRiG9ETEUcZrmmjakcJv93lEC74DtLBjF4btw5
oJwkjvEh0glth61DKqLMDhR0cLqodUUV+nMeLnPNcp/qUnhdaOmv2XcmrR4gK9fg75pC7Jct79YK
sUud7pYrJ2/shMYKZA2MmmLTWEQnHHrNWJ9xXb/9zo3wvIC73yProSCy894dQLnBCaTigTj3IDvb
kqovjApmeQS6AU0m+/O5gaTeu6F2YzVN+PJ+HrXbFTZLIg+Eh2hye3183DfwM1Q9+QbSBIgAgxNh
jN3D7/wgiAc5GbfxC7aQwRG7sDjDsTLqXF+KobFFaAt9WqRy3w2+dRU0CAe9P71CcEj6Pj2tScQZ
K4KEZQnaZ7F1eaWIZML94V5x9E6pfdenDZKFKueTSdeKl0BlJg43Smw+njFkWj4h+VDvppQCFfgN
VeTrBwLMVPb3c/S5M5N4MtR7BJSqyg2afNNGB9E9WmDvA7OiXLWUW3Dn+sHsDmzfF5j0e333tOCo
tfpfuKhwZxn6WlgC2rVhhu8smrRfwynZeOd8KuY9gLztwmovCViZEWAdKidozCVTDLKTWmi3bOFH
anzSDZTWya+60NhFap2wnt4MU2kIZ0qT7UpeHC5GUsQ2rWjQHRpgu9EDHqzUB/BUiRm2+U03QpxA
giFIaae2oodJdJ4rnxLinw25gOHAaJpAVTujZaXWuJR2SkI3cq9wY9np3h0VbhTzI9Sei38dqqoT
u08YmiAweyxH4o8t7lnaoWiSncUl0EpxjKC06CxZBJM+hLR2nd+SLNx0HzXjK5mFrAY3MlxQmsKF
JGDnBbjw4zgdZJtXPtYIYqQrYC6ahdXVY9URHIpaKVeZFt3ANwfsIjutXIscmZ1YmPMx4RQ4+n5e
5NEa3qNctU61UidXDTCXww1hFqWNyn6ChQFvPUXOJXI9XPZD/QJGJRTBfQmqhvjFXVX4aCUDwj4T
mi7ofjDD0S1ohmq6MF4n9QRcwiEfXroFLuC3ZNGm/TbufKVjkoClxUS5R1e2nUoftrbOSwC5/oMo
Fpa167/rW7XwazbBBMUESvgGcOAcgs4mAbwDp/slcccRgBQmwNsSWAE6rG/Mt8qHKRp3Y4jD0BMD
MsIVH9jIDvD7RLAPC0kR5Z8ww6D2TTwNqss5tNegUf5P5duD4xVcQ8GzayEA7JWLvonAcRuKorV8
d3aAteXUBPsrocnQyBGM7AAlXMHskjDNsQNZSXK6jhjZ6zfDrq1wBxY7TKLsMfSMpzLEcConW/00
F1ZibQDI0Rb90770tnQ8L9uToOHuKtGJoloT3mmyNXw0HD3E90WDqcK+lwvJSyU3FbDRhngYE7Yw
XrMMHUJSRE0nmsDF2hy8+/4HxFDXCPefCCzKddDPesXU33ukteYLtpKNGCcQCJ9Aqchp32QVYZfZ
HEgzGcpxfD4ayMHNvs/5Uto/yCZvGcMNake7w+em7uplVAMJLsYaINYVaC3FgwUDqXhkfCAJ4hnU
xpkSx3KW6aJ8I8etb51C6/vm9T7El+Zwga275d/DCTw4VE+fvYfgF8vW95Ts+iiPqB2sat68u370
LC6I0zbHstfN5cOCiiJkk16kiW28Uq7Vknh3WgOitPI+HGCKoWhLQg7OACninwPGeXKJiY0r3HVG
tYI4BTomfPO6eGgarr33JcoIP7kbWJfuhVKqui9oeRG8TuO4/F6BreLRCm1tmV311N/G7NioQnf9
zUET9THI/phxrzlNZEJT0F1ajE8qPnqR84J3TtjR5fWK8jS/i1UZ95qA3SlssEQNDbPSMIbbuf2L
UBopiayi/Tuvo/bTR0Td9L7ZngoKJK+2Qh+ylsjS1b7X7j+gScePju2JIJEnw1y/fJdRynx37AOo
VAKvRgKbh+kt3ReC+8n2Ka3n63fdmqORVpqHe16UFlSlswit7KBcW5Sd/FbHTgf6toq6eR93ncwY
lI/373uaI+N4qlMhp2KiKpa23mQoQJ0OQkItVsAh2vHfxZmIHE6tCIWSD5JElzt6R8SKeWCoL7Q3
ZNWsN2FComLZOKJG4WMle4Au+hfjztaqTD3Ai9Xyfvfoh7oK+O9QxWIds+si04V2jNwwrRnyRSrK
qbeTz2X09AB7CNdOcb/7dIOvNxt7+tYwOZno2LB6notPCcRZ8K5iwEt8zVjrtHaF4zXX9BrOHs3l
QOZB6fo59Xb7NU0Uxot5SXumlrslJyWboZUg/foL2ubdrMO7Mvbh+ptiRNSMoaTmlo2lalp8vsU5
lhF1YxRu9Q+RcnA3qD9V5py5szrOg25ZW3apeOfbQ6ckCOAeZsgNjE77ZPiSt5l0sO8STV9Sj3GK
a0rR+74Ni7JsbV4s6PN1u5Otl2jF/O9c0CQU7qH/J6+izI19ZB9ny4VQx5PWC6OV7rP1lR+SN63o
kg5hTsNHsU/lSgmDK0VutsxrWTEVUvT9Dmwr4z9eTOTfW4QMzoac66Yy2uI+eU2WOl4A5dL3nNZy
Hx8RTM7aIR5C0mNdEg00p1n9MJl/i1CcDsdmhUS9HjWzQ/fvoIlbp5U2mfp5nJIla0oWcOKTcIVL
OrskPU7Yb7ONo+gyuiC3M3p9fpX/VVMmGUJrIMnZTGfn5l728xci/3TG1tf7s7MJXuu31EOtlWOo
Blutez/2qO+L03jkseRCXKvx0ALMOXxyNweVEURTrIfA9rd0wIIaSoZ/X60upT3ITmaiiohO8bHh
G6VLhSyc9ctjdIsHiGjNSwVia1cMAmKpiOcGiEZtyVvulds5ufcDj5zayn/57dwfcxs5yeTCAyKJ
tlrRp56dwlqKNXglBwcMMiv2YlG2Z/zIKSDDq8jBOJovwawADJ96VMcDlP4492X+PRPqQvtj0ngV
9e5yIJ51EY7Aifub0gzU05SuHe0ODuM6ephEkTsBOyPcIaHEGqTg89vmcvAkhK4Z7+dHrwClyBlk
3E5/P6g/4nVq126jGijK1dlc63M0wXQe1+HOj+DMYCqabxT8wX61aN8TT0FTfRITA9F9WFeBPFZL
bHyVPxYHgCcDGNXSgzDISM8EwFqTWVXkhQxmEwO2MEm59LjNhBIAv5Bhrcq7oiiZNDptlomktrup
B2L/QYIjZ9huNP0+Op8B54D+M15wxNlSg9ubWv4QcsMFTQw5vdSER4Y4czE0/rvQnI0FLuoxTVUT
dgWGyTUbZxUg4E1TAFC7As9tsoSphJnBBw1mwyMclWzQBXtihWUcLZpTFf/xXr297kzomk8Colt9
zyDAOs/Jl5Rok81qTGBGcVNPTVhy/PPL5oaWyiH+FfzxsHX/YZvCnJD52Z6SFXJYWciOCLf0hxR4
N8VVYGt8Qfc3TDi51GP6cW88w5v85ew2jXJ+fndDqR1lWmqapkVEtYc/KXF3NKc4zNnXTNs6OuNj
4QTzEb6ZNzVzSzyE3u3MsOp2cUIuUxlna8MM4hibOsGZqhmJ32mk/t/KEgIs67yyS6C1hVhBHu4J
nonN/gt5vD6LkvnsMmI3TfUYaJQB5D9Cq9zIh917xdJiSuGc9bXwbEUTgT+yJguaUeYg8siN36Bp
uIvQO7gr0oudEbjqupZDW/EXYLFban6gwCoCHT9fsOpuq7TppgqMNR0VEJKOEOWubAt9HshZlg8Z
kWeyTpfxgDOfl1cakHJCRRdwIe7PR5ELhglcWU0v0Ml0yknXuzEh02KYJHCNo18gsHdSPO77vguz
IVyIkFaiFtF0GWW9urkxBet3zudx8jGVtlU6FSyka9q9QaDC82INgsntTDzlVq9SGzo6ElN29uni
J94PyHGH1ew7CiPnb9jcR8gyukSBT4In//J0K9yeHveg3QUCxrgOej8UvaJaP+9mzhGsn3ljYAab
RaY7gpG4vV/7c5+2TNr99Fr+C3HiRHqucxh55ESzGhaBatk46+Qs1D6ItvvI+cpwmFISBKrTeffV
0MX/JelafP+hAnNzmdV8ln/GK5rfbd4j/0U/AvQFi8un9R5uV5esdvV8IhHNCbK2oF1QHKxu8Fur
kU2YMCi9kY9vu2kGXpxpNyv3eViSzo8Iq+6D1bMIV1m5IFg5GBfBVCGkDBjdIdLLVScPqJzmd7y/
l5+lzXa6j+HqKasA/Wk72NKK78x6LSTSml/Hg1ibnK5Yq6+uqL4yhrrgMYmPjfeWTwd1t3t9WuzB
vtFZWaOZVlMHz4qPXnJIf+MNkZpxp9BVOxLBteudhRjYbbWMHlcwFR8evTC4qg2Uy3J54tvFz6Cm
Bu58BvBpiu3iAGDuVrEWsmeDyfcwqrH2jvt4CRMPwfMV+uHOc/2fn7JJDTwdvbt754xAryqhUOOW
v76d7D/D+rM7n9LJdms9VVLFCi77z8Wmu/IG0Rq6A49mH6gVTFaMxKBlY1+ZpMkcg7decNpUoyMm
j3AlC45wry1piRG1UhdKFASEagy3ju8+pH2cfuDGDLS6skXWrz3jjrXCJeQAECO0LswiMhDxjU1U
dM88yfVdIs9e6QxS2A45+WbxZ1SYx5fLai+/s87iP1D0r/1FEehOxjNsmCLIIZ3s+WeJZLcgwkxL
li9tk3UxaKBJqKer2K4KqtrQYITecU5oLsnKhLd0Frf7nAiYv3TcuZYegjlkx8OSlLAJbttQ5n7U
p/Bu9iRs8vJ4Tmyvar7WtAQP1WHS5tRzmAnfruTihWYhk5/CpGiYYSSrRBCp1+4jitlNGNDj6pna
0WAZQSKvksF1yXcpMNgcHAdDhY4WhpWPG2zqeNUuaRheNEnif8Hp5mcdFVWCixxPQGvUBoV0n0J0
KjsJtWaD+wezLnKzN2PB3jDfOe5PF694UdeyovUDAMXYHeqjRKKnIasn3xgT6CjeJobsyWCC0itI
BTqtCUDoC6ZhyI/NkOmjcFRcj56hD0XlnldvUkACFA63VyaOPgsTw7q3BShNbsBpWxxTabzzHKuD
XQV30HkhYrNAUaMdxjk2JjDCVTE0KB+u63Mp1cBTlylG6E0UP8pQSc8q5J1CepMszK1gGphfulnY
zrZe07idS1g+0rY1RSLQ8YO8pnBPBR1Wtc1g3l181Au59rcQK8cfGLjpj68slXAkxHQOjY7/Isj9
kiIYhJU8w66/367VW2weIMHambCBw6Z1SuzxeqdN8g0cPDk85pocsZC+xBMZZ897QHI4Zrm3kmE0
a1LUbV7BoDxG6cm2FiAMa2+OXvTsYtPFqS5RIUxEEXku74hhjSrenXyeDEZSBEnY8sRPXM+eaHw0
sZy0/1bp1r1JenWwOtNNZ0uTtzTwRNRuzCNU6S2lV2+CfmDXjgSQRGHqI5A+2Ncd+h3nESXbZfcn
cBqdFZ9Y+LXOs39aGBcJyc5J5dLpek8ukKwLMgFgNsDuffZpf2o7xa1BkW2WSOQPyZAjyMwWTbU6
/o+IwTHPHt011p3COSNluM5DDjs7uQeuvhsDaBfxjYMZgkAphpbbO5cBWwK6AJ5e6IX/Lt2WUh9l
EgPGitaUV+NqGX7TUtcaNusvGzUhllIrvh/ADXYbPBqvrdaFLEuVRv7ozMt7VUQcNr0H5VepSrt6
RpDMaZMd6xs76n84MbfDmb9bko1bJ6HI5RIvSbAW0bCxC1zLtaLNf+wK33+Xbc+P0habH6J9X86a
uS1GfzWujIAOd2nRl9428k9q7wsugN6MoOoyr47DG+bRvZbc9oCLQnZq8NOreoaGQbetU7QrGFIy
lb2quat2lZEtxENwiTZzSRELgRt1p9HF6FYIG8H4mHrMbHkFimvysYaeafsV/iJpThSlUu6S2yG5
8s8ZFlrWSQJqYPZMMRDbWeX+FKnewmSKHiCpJFBSpiE0paviYkefqJ6yW2I28KJFbTtWNJR8OBPe
Z8NIcYJWrRoKANK7tB0ZeQ5aHtd3YK0Wr4UHjd9OIN4GSjPpWu+P9Vqq1NuN+6QpbXWODdu1uzgk
0RBNZe9jtNx1cFFAbz6QsZU1aNzFjJsFcK0j0OrVXBvsZsFm++YFPi8tj7HMmtnmAjivcwID91m4
94kkikaOot6dTGwfIkODsYJGqogeNj1MTgsAxIFYBxFdFVG5WuJ0iFrtquSXOHXG1iP98NFp7LiO
FnUdJ9uf8Awh2wn/vF70FXQ76G5JvWZwqn5GLenxuwN4GQJ7pPbnpoedDF0BX73A2vyzzL7zPpWM
YgpYEWoxlisSxBqIQAbRVHaMDuo3nmNG4MqnSkmaSCtv7mOTp72yeVChaCKG/i2vBpre8BF10Wsu
AzUcmiqTEFGvdjSqWiQ0n8lSs1IT8r5DsSavDWkMe4nRBVuLHGUBzE0f3ijGCYGnfD6PHdOL0as+
7Qcls7N3gOhEXX8QnBXbCTkcWkip/+CqT10bgK5Aw4fMmk/WKmJztX9poN9uTR6VP2IGBuu7+wKi
kgayMU0GPVsmtV35gjnz27zgNbWOgXCuok6xHhVh0BIZf5Fb1wTiQcY4KmaKdDV4V9OmBLJgHxar
+8anLVV8PgRiMWMREvb3z7+VKngHa94HYE4OydA4hmTU7IYxLHi+oJeXWqZWHHR0XlrV6QOQ661u
EcogQwxFfEPupDPWIsjh1VDwn40Mee+giJhxKk5XUs0uzKJzTZqhACOEbx3mCewS4BI9yzXLlx0N
pJnLnMHscvIuw23yRx6fn+eyHq2D3iMYCIX4JZokLA4PfNOA/6hozvznC9IkdSKNEAlidL6tQjsC
flRFCKR8pYI1AlR57pZh5Dk/AaZhI+j4AdogWJKIimvzLL0nDJlsZXZHdpjLoIdZOigJA5had/13
yhXQ92Gtm8KeSWjK0bYuyj4JM+CiR+z3zRxkbcibf81gIBC7qSLjdsNhmlQCdE798XVnSzImM5nt
w7XzBqvygLUT7mkcUTYG/adcCldOFVZS0q77Hx0OycXpjgmNdgYqq3u1aXLk84JPn29oZ2KmqP8q
NKVdLYKNxL7W4KwnRwkOaJI8etVupd82/EXX2nxuRmb1tBkIFLfjslv9YL48/dosrQjhsL3qLof1
j/6ibFdCkeZsPGHoSdMUw8LI2CRWzX4JAZ2NeY02nlmB8Xt89gd63c8+hkR9dgZ60f9sVG7WNvwG
umbje5TTYFpxIxZlEQ0QyKC3mNpDIbNIcMVSddFVQ0TJWMDUqjErARSSj/9I3aUw+m+QVTPOrCvI
ewlpTAsJLd/2EA8H/Uic+GPO2w2nrEUE6cySiLgsSlkF2K42Sxa6hqM3s0qx58hWl2Z2AM9sY5cQ
qyRfhth9rkPFKS2ZYYF4+1IwtG0dqNipkawcDZ8Ft4LMUTiBaa8yd4wtNBeGLJsjhjJ+5delXvgP
Ldm5u4at2SJKgwUTbqj9IoHIU3dHBbHdo9+8wcW5+l1f4B8EmpH6Imcha5UMcoSPQnNRPVv6qW+h
NZVpmWVmkO9eHC6pdNvdeDnxv5mlBh0yrVpd/iCQaX9D2h7blpw3L9uCNXlM0OQmA6zms88RDZrj
QhpKLqjmGe1CbUkHq+WfLlaFi7wQtLJYAQipdj0GFyLpalafZg06VLtX5T5jX5ggmyRig5UPIauK
Rr8SGNrnZ4AbUifCydm7dZpzXuZPRnmNlJhWc95zgZ3hJQZx5jaAIGh8C/YXVhL4hFq7xbyAHK6E
0mQ6HWTnviJxYr5yinc+RnKpveVb9bODI/WuoJUYutb8mp63jEuGiqZewft63pocbnweS0qaq6GD
jWvJNAjFMGG156xwsnQ1V7bqkgnfKPfs085ggwtmrydajyUEt6r7wOjy3KJCdfn5kQnf2eLa4wwM
7BvGkuf9f3QEhyp/dWIoURaxVF8OdlY0XIGT6xgVlr81yN18w2eITF95qmdsapzg/ErgDzP0Rg2F
3UM95m2TfL8/XVx+gTckStUza4cSF0WA67IXYwWDH2nxnw6n5y4jKE0wRg6jDIdt7UwMuWC9P5Qi
9CsesH6XZekBlvFGK2305i6g39G1kBSjMNWn0hhhyXPh0t16o/IkrrtJ8vE0R2nQje8j5hQPd9sU
YdP03Qn29xhYOUCfpGDCiZGCKhdBjNTJTMh7+9o2mBNU/NnuGAbZp2KyuTzSOMrDBTicF9wr/j0R
xAU4CQXbTt38mDS0qWOEcc865uCfOcLPesgiiPnfVVvffC6UXOsIRQ2XXLHbxdkijzW/RYrZ7NlN
QNr4rqBADlufGkPjp78V1wBbONOcCChZiHWv77K1NGa+U93WWBtrJM1VkiLavHsdF30YDDWqwksz
UAoQVDIWHAe0qF+zBfRWNLZsVYj6UH27NOWqMJv3EGE0DYiD322NaSQLJwY7XItTg74/ZQE5MRwU
0EvnKfluOAUWYmae/p9Mxhb6sLKfVam+Q8Wx5ev9i0Kc5TA5ohmITQKt5fYp1yyZjtltO2BeZlFe
MaDtQsTpnBP2PRIZ9RMuUAgV1TCKfGd55Dkp1SJfagg40CYMWmiBOwW6YgMjSxIVoQzVnna6PhDK
Kb9IIzTzP2Z3uKkIXMgPklAkThb2Gu1ugVsOn3xu+6ubaXikD/EF6VIXkh4YJ4YdP55fP2952i4k
M2jTjpBl9fVzWZ15xEKicGdwu1NZfMOGTgM2vdfG588eKZVe0XJTdkdppeNbGQSqibzMPWCvrZtA
NmEXqPFB7shWLZ4fet6r9ak1srftYjg+3va7+ZLU96Wq2doI5B/HHKqJPXialu8x6ewmKst1rBfJ
AC7OcyN87r08xsCqlgO++xVhn0aJb+sTsBBqqUg9GsChIoUv4gY+N9BkW0eVbqoQhEennD2f/D0D
47AgbBJRLiauJXySZ97WkNv3Fmvg9+YZ6sV0aGLOvkSmSGN4B0KqcRpuuAgfFbqAqDIy4Zj20g0Z
a0FriA6c5g3SRLVH3VxHJZT0wLk5wPHufVDtjCBmv0ZMM9ma/X7uzh7+m15bpYOpKBcv0Ww1X5OP
9BffqKXo1eai+P+dy2CSFsgdj+Q76MWmFkQTkWbX2S2IXrA1yK9HyGv46G9wETcm1ELqpcqRGnR3
eNhGYQIba+DbwtE+xG0HNHx78ZYuPFhuimAMkvEEmm8eOLjKkbTM+W98ZqKTTZ6aLK/Ygn39KhTi
U5Fh7cTXKllD43IMyD2pQkI0HoxXGpVJSHbedlEwHuEY0FD1+pnqtub+G4aMqfpXovm0jl9LTR65
kLd0PG1RFMTlpJDnEgIV+21bojf/dz5xd4R224P+N1WWmHTVq6LciTbDrl19fvmmiVjea1mjWrjl
DSjZ+A0z3uaItkEj/z3glJ05yBXI4ZTKSc8jWfZThYJ4fQKKwpMzBXwR/MGuu2qpCqwH2qsJY81a
VikYdYm61F9TLtd04wkDO93XkX74wJ35qdHnviIVT4r4ZnO9WeD62jLC1qyg+DLbFD9rI7jFj0Ab
HEXZ/vDpExjEi+BE0zdkovxHNLrNd3TnTNYOT37jbF0B0o0ad7Kgi9Wk3RgiHc6X+z5DapGMOE71
HlUzwOdZfc0A7v1Y2dAvkjvsKurestuHch7sM+hJ4fCeXz9cDVXpiAzP8InC46sTjFdLuvgx2OnS
Ebnp3w4YqhbLh258r8LX9Is2rGBWU2rZm3kxJn96pTiMuJAslX37PhPyg/rlEj3UUkIfsh525hWI
b8AMdMfmNCtdyVtxcIXRkR2yHkHgvznjNEM1L4gHzhxHyC3lSKsP5bYwehENSEwvVVEQkhosyO6i
dZj1Al2JkvYxxdiBvnedDpgce/PLa2U3vRY5+yECjA0YE7jFxD50h7+e+Fku/XpxSB8utvzsxgqr
rZHw2Kuj2wDkbAXJDdRwZziOtjzp0af/G4erBu6RohH18ioXzNARvg4oUU/edu1Jxi6tLqQfdR8v
oKOZ3iNA7l7Cn9bD8jSloQdG4kzr7dMb0yHOj0REzylcJWzgJJYjsgp2UjIvjFZdz/Hts97+2cpn
WfV86VzebRNQWy/FA31riWwNVhhtGAtUtsEZzgsAhMvG3yT2bQs4c6AONCq67C8NasU/N38rCYwL
17gmDe62dCgC5/heghVLqexxd3WYJJNIBAzbSBfgEjziipcLK9QZm1+vTp4hJK1fNeeiuLs4wGI4
I21FbFvg159Xck/lOormpVPyLPlC8joRl1w9M7f/EpTJjKkHGVT1Bxb9gm9EO5LHUgvrTh8t9+7A
2B3lRf6+XhwJEwY4lTh8vCk4eBwh4vitOPS2ohQBicqpQV7iBYNgE1hKpdV2XoMPD6su7qgqjUF9
QpfclOtEk1YL8gnor9QJX84L/oiXpxaN5gkWuhtqBgbaSJQhnCEkqk6+LLBP4BKLe5/BI6wj4b95
tiRSN8vnnvafEKuBbZjOIBPkuO6iIK6EgyQ6k1j0CbC0bQttrFS4ioe0uobc3/ATSVc9XpCTe3+T
GlfjwOgdL9EtQsUZJcBp8B8m8BijgR/cUedI3kCznE5q8IhPR3NCcoXCAUYEGTWwFK/oQIF8F2pS
9E2/E84wuRCRUkzdU3PajBPjPoxA5S5zMkyUfA/31KaUEO7MJHIKToUe+W6mrdPT/Q/RO54+gnqc
BeVUTKnH2mATzT9FHR1OkugnL4h3nYcUW7O8pBcZG+XbGol6g6r8JGERXHdveQ4pKKnPNIzViwP4
kMHsA+lCzQ8/VSUdYlTh5RsnZjFBZZT0pBBRF5i453fMf9MzbxrhnOpv6y8ai2s0GvsHeIQpAI4k
ZyA+sNzTCIn/aVtgu4JbbkrYN/o4IpN0ieJ4sjKSUw6kU6a4kD8tMOOdzxc9PvkkuVvEb8eORnXe
BP/qxoyUGE14877ubE5XB035+pIErHvDfyaL86Nn8XCzzGp7mDycjSu3CAUNd8yeJ8iOONbNs2f+
0yRFbp6JMncHOzhH7kURr5nFmwtMI2raHx7ezTtEn8bf7plS2r65SCVf493BYNRfP2WRSloBbx+o
A7PHFLh01dTDiKmOm9f9fK+KrVLfPSB9QXqSPfGuvZ7PVLjPet1nHbjw6yYENwqLh9nulrkgTE97
Kv6FWqx6aSBkgFsBS8azIIAxQJ6H/k+QjyOaySzwhlDhCrZ1OWvPGFsndKnRfkRqrdXfiBeRtu4E
K4oHlbi5daMORSYzh3PAkxonkQ16maUNnJG5+6tU39LpePatJlKjnx0ZkxAOxjfLf137no8K9D+8
en/bbFiKH/a4Qte2Jhd1UBt4pyV5S1R7+HUWzj7QZP2Qz3Ty8TIrQjh58lJPqUnN560iygA2LrGh
oH6pXVYvwbLQwm1hM7sCBFraUITnC2q20PEEvolF4gwrNH/QB7eua30VsLRa8ZzAw4rDc4lixWux
2NMefNGYF5HUgmcd8zi46uuCdYYuDazAaACHZhmbwFnN8Y8FaGL+uYJuwMqnYdQ3O+rZnE672PCU
s8wGqScDjePf8ew6pwrwNM870BdBtfS56NIFSFPwPAWtHwZOJ0R9IyLHoFrQIo6KROMKOugEb9bJ
2dODm6fw8o+Xw+B2lxFcHLkpfp82dUX2ozBzZkwfU1ROGkhnIhJAxaUlpN0i+q9Zp7sN5Zqq3TrR
fV1pO4mxSiCyfA3uf+uEDy3nwv3BHAT05wGZHwSnjqhRqYQj96PyRAxY+Qg1jMff+Qq6ZxzVpj9q
aHIsPZE9iM2ycL1muhGhzckn4uEKiyVEvh23/U6YKB7G/1kqJZv/V3UxG08TCa9WmIqTvMV9KShL
GzMH0CuY21WFBk+cQNho9QCdptz+gdZp+Mom2/W5E3CiYNORzC+eIxBvKqfREUCn6cD/3VZ7INig
/NE0LTApn2DnPV6bJBhwe8k2G3w0hYCfZ/Cf5LXPw+Es0Fml+/e1KL0BW0SNUMcL1OCsIYkJpqkO
muT581J0LRHV65IGLVKecmSBf9vkIpGmqxprattIjMBiNNK7uJ56oNhcMMD/+rQnFWDE9AIL4A2W
a/Wpj+Y34FURtDFE1amfpguG8U1YWz+Q0eKu1an1f5C8Vp2kM1jyNIzDTxfE0R/vCbDeuy5UC7Xj
OIG9Y2UV4sL7imY28Y6WhWeZKpcZ0TxwalbpiZ/W8hZmEXli+NBaHpGQdZzYwkLSdyCb2XdvDl96
4A8LAf5GuIXp6z4bmEviOlgHzStT69X+VxVhxuSxACGGXzWNMLSa86Z4gDRXesDzSw56V9ZD7/XP
1FH6oYWd086Wq2tWFnC+cpxToAVGecVNgM0u6LmAbqrmEHyXJ1iGqwkzWtM7O1UNxbYHN9JHcTHe
sskGprL59oNwahHinpe1Es4QpsuPJ9rQzcwMStXYZhbxgD0bLbQ5/nRlVaYsh0LCwCnJkwT6m4nd
/lcjEh3w6XRSbz/qZyYWt0dVlc8GN5zFrv261A769xNyimnBfk6vjiqPRq9bV/cmI4Yo3o11ni0+
mYKHNM5KGV91hSmORyqj/JC4VaTNMw+Bpo7b6Ib2xIGbSioIV3Dap/BV+Rcdt/Ogn3i6guDUZkVh
Z9EgUs+WnGbKJgCAlMQtxl+bZuNHrg3CP6nSu6yjaaYrm7WKNLpw+uJloexyG+x7NjntC3PE/Zoh
nx6GnsUjD0gfMusnDlt+0StydejWyT+RdW8yifDMocfyhpnzX7bje/QQO87rFRxBNcB5ZeaL1Shf
f0nyTU1KNkBJEuwYheha+mnIp0AsZ+amtDh9qOv/KmUmOYjOKzj+pTiOL4FnQWiHaIZY+tg+WL4J
/yyuGeR3PX8Vz+OnMKSk7+lTyx2YIhcDPv3DjVmOfMKwmCeDn2ykWReSYMzk3QyafEc8J5G/XwOg
HrDmveZATXixM/JkxXY5+wTYz8YpNiQVYvIeCLuJdFN8nZr4b06jV++3Hxzu2zHIjCeukZ/YnVuE
x8weQd4pzitnytnx2k72nI4m1KrKQ56zSjIwQUDeS5F1L1PwPbS3fJANF7wG0o4eVlhwEp4BkgIs
HOmx3zlkrM7ifvq21xHFv0hm8VJ7AU/IJ8uau4SVb6DvmAfEUlbnPjnFH4qlVkOTtlz4WasTszn/
gq8ncq9Angvk/yG7A2dR6kMkIO1R714wcECxBRJgE3Hp7AvW2qsAon3lTh8VJzRqVAVVxBoCi1vk
W+XAlc1mePeXPbxtPm+tKgTVFkHO9L8HcZl/ABruxHPMvZGgh2mmu4kaBHJlnx8pVPAkxd3rkhGh
7MxrYE5NSDheLK37cQiOaYFCJmiVG41o9BY2wtW8afMVmek9tXMu2aRD4h5syzeqH7lI8y8+b3ez
07Leq/RPQWzt9Q2sz5xaJFu8MDhjeVxgOqjDfviDMFE+qG1+yVhFGGyhSnkf/Jyo53LSRpX2EOZC
edBn6bbyOg4i5Cfw5a822O9RIJgbwF0XK7jdJtK1e14iDiAj/RC0gobWv12zrgkHLjoSXjIWMFjf
MMyUZEdkPrzMJ5djI9s/hzSWOEX4/FJ55g5C1lA+zSwImNRkfg49uYzelgdRW4eXoYbZfXcVocAQ
Xyg6cgs39YvsEUo/8BcP+EarKwWYclEdBw8XNL2Y9i7TRUw4ucyktUHLSB6XKLAWIzSovNbuH1QK
JOz3jh/hyjrrEVsFNno8rmeqpK147ffJFjv9qtQjLZfiMm9sGX/KAfTgrpYlW1gqMEIUg3jtqyvk
aLjOBV92N8WY5KX66vrNjGoSF2lapUAObMyE+4EK0VBzqSD8h+LL1pvGobs8gCuozl3+mQlc4sUa
twTluHapA+H+p9xq8Z33fB1gj3o3yuDLAhVGlfcXlEiwmSc0ZgVAj0KBWsoZvRcHNW3/6poVDEdR
rmYDYjVZH/vfqexqn+Q5qy028bbUYX4rCpUTZPjcQT6++ptqFkX+SwFR4ssLkTfjWsIwjvUoZWuh
QMNQ/pJEExIFLVgGtClKien7ToI64INGEDoJfRO96PQeL9ZhK4QdiR95byONgiJuiKlFEi9Fkor3
LLN8xqdO0EU6hDDOS7TROdRJZMRdf/KCj5ogjJ9ALbra+CW6ZeybY/qcv5oRyVCjC6ea+JMQSVXR
DUmFPCQfWdBEV891YzZZkLko8pU3clLLCMaHy6gUd9OZKyU4Audw2HvVEP9GmsDpnYgGDJ826EKk
ooq4LeQ2epgHwm0ejEp6G4Z6fFoF3X9UNDx8eKrMwr4sd5nYiLyODsfVRBggdMf5Me/6B4t7FWKT
qyap5jS9zTRAgtr/2ZNXS4+FssuQN3iv+/01YMsPJ3VNaY7lZplIQijTSwG+Mrt2kqeDbIraO96d
bS1hYZfMbyqdiXNngcJQ6Is/aeviqrPU6B9WPqPWiW6210bv2CeL02uH2D4Qk01w3FRiRfME4zhv
gYlUoqCvcf5cPuQJx7RK099HNMl3BRZsIyemDf8kHopv0N+c9S8uEuKVAwkq6FoaLEzZYWCNZB0a
WRBclCPE3uKk23yYLDXDrik5MOk3tEb4zF86Ep04TEkCVrl1Hc+jL0UYTuEKRoyHVsNJsncr6d5E
/QPr8qtOHPvaXC2h67bOuFjYUWTiJ4qst8XI4uXj++f+SNFLYtGGoaO4z86yGSIQEyA7e/3s2dK9
RQbsklSuseMZwhIhafNGNS5aSwA3/xXqZlF5pM81EESZvqw0UtAabw3xRo/Txf0R5WNbmRGRgATA
/OmLbT0rvRrCwoEgZ0fgNQ1Vxwtao5IBdAZ1N18pbL+jku260DsjsJg9sD/OQnZO75moXnRkkB0n
8Jvff3FRJSA0DQ34r6Y7IxtBo8mBVNEtLkg9JO62E4fbubabZ0YmJGzk/ZCk60lw1UurUUsPdtev
56ZObJjyawFeeFpMx+SdSRg+K7lwGOWKE++4osUjdcQSA5wEvutVzMC5aZnEREDyRSIySuxI2zTN
vbv34bV2ni3ptcFjrmDqs8TjlL+ePWe59XwV7iYUdyLd4LoUlusvrIe1DyBINwoHwIchRmD/4tZp
C4PzFxPDBJjH56bk/cnTxqJL537QyjyCfASNAyvasyiMMWJ3Ol62knABGlwGlhgvMsnn/VJEQ6uo
MMeHK9ZnAy6w17NQ2zjxwBAeglLTB7iLL5jId7lYzEZY5JDWwhaFppBNX9Izme49OCiUK+z4xh7H
HFmIETkX0MY/qbO6w6q16CgpjqG+xZh8uXe6jLorHITnkC/KVh3ujArWM0ghLwW0ajmEBPbKd2/N
QlZ5aBj8l8iisElvNXuzb9HFpZd+YXQrHm2qVeq2rCjCL9YI0nCy7T9uqeAJ6CQO0Z81I77TdpPC
D/UFygm8JGuBLuo+h623kpmaxYVE8WQ60+Vu3uEKU3wt+Kl56+z6r6u3DEhPUEr2DE/gyhwvbvYN
pZrVtVuf64h/UJzz9Z/Wg/pq2UUXRb0fIKMRtZOG33DIT2AZxPLZ5w/L4z/91C1Gf1FlarXBJITb
TMc2VCCJmViesaAXV2Ypr1Q5p9Kf6wDnxeThKV2L5RWQEfuE7jLoEdzQoRMV7GeKxDclcXiX6nmk
ERxj2e0aKsYo9J2D7tQq3ZG2ZPCqH6TvR+NG5pIrHfsHhuo5++5kkI477wZ6BGkWnVtIaoT+/HSA
kh8l4fokvr68TY+0CI7THjQzWXDyITCbyT6SH5r29mU/mCHnk0PlPrTNfOI7babo+62uKO9Tt7q2
H/LTZawILSX093GbTeyXI1f/SB22fq/4HoFBp00p3pcUPaOes91rYjzs+tMYKIUis3Gyg7UVT90M
3jT6frwVS8uxi/neRzK6yszTPVeF9+bhSZCw+Y/lhIO4XJbPH202xIGRflGOHsbCLF1x4bDIQcfb
OHTLG907rypDgf5PByc50dojK338diZakbUad+nx67CxIJnVmmPZaffDeXL+9UJUvWmC9xRYvg7m
4f36ObzhqnT5K5OqULxZLDvDOBnZgjexeRvgCpehBiphCa7RtmPF3E7lu3MlFUdb/x02YbGjTRMG
zT+z2nLeyn1o8F7rUxp6gBYymcxnmlV6l0xzzP1akT/Zm+OpLfTdmNOGsQOT5ggLTJhjEQFs6yyg
/uRIMC/DvtcnDgciuXHPKXeKa63oxDsyW+4in9jGzZV6zXS/jndqeMg9PKw8PWrnZy0mM5nhfC0w
dlA8le4FgYO3ljTFJVTZ217yXmXWQlOkO2IjTCUNxJWVw04ybRsd/6JLSDJCoGaW/P3KuoLr2tI3
s/x4DrNkODhqTe5a/W0HadXcupUgRgSR2IDz93yI5YkGgs3gRSQriyYX1Czpoqg6Z23xJMZpoDtT
nsWAlVS9bodo+JqGdOVSgbr3IbkOygo8m28VpTT9zoVRR7ETo88ChYEzJyYCVGeuuhOxHKnG9hRt
kx68qtbG34Jl8w8gV9Y1PIXqWlft9RuokEQrRLQWd9ZbW0C39aOgRmNw2cuZ9U1Aokx4Y+xdPfz4
54LdMQZc7K+PCA9dJ+qUEeh80dbJsakP/t4TJYbNbf1Rc/mg6mamLq561Wq+seJ24HhfOZHL37jC
rQidH3Jz88GoqTVFOMWhRxddcjXCI8nIoAFUPFoO8Ct4RUii4VVFWQ5Dx+Fz7o+9MIL4w3EnB3vA
hWc9FMe+DCUpGqXBJ7BNjElSqhsIGZWoDwK2t1E4ugYPlgHv3w/dn2sOwp4do+fW0I0it/xZr2zJ
DgzseptyqfokJyTQrtzi47mNNUFCUa0Bq7S9wnE95eEVBYrthk+O/gUVTm8snzJ6Uqwyi07M0ToC
z8buIjmATQ2a3R4BAe7tFmnmivHvixEK1UnKRT+yXSgXozARMdttgcAZsJkzhoTIxS+oUkLRx3hx
OY+tg+NChfy1R3xhymnBoTL20l++4dbExtsJo3jD3BExfig3bJOSQbFRUsyTaRl7lLUn02DgiF87
r9EWXHGN1Wf6mtBrqajMqTdvSCkXKtBURaf2LOSupWyB7t3omp9aG8zsh0EK6w7F4nlIMaBbP9dp
Sw05zLhn3e28n0A0o04VmmL9JnF086W3j56Q2++sCnK8IUoLicyX5cPEcJEh0Fb2moKf1DBVbJAA
WSpr2XjjbZfxeTVF/8goaxpTVUCckwV/dfV4pZZDkx88lRH4GGJRG4g8ohqK0VaJ+Jl/920gIrm+
u7i2SWb52/bvizgZBlBkbDtw9GGPmC0mVLmYXHuRXOv6E780eeWo6bFpVn+njSwnAJWWHcHATP7r
VY1ZAQ2HV5MNNDjRe1wxKPB8du893MXtRaAGuMZOnVaXStBiqKpfw9uIIeQ5icOhK8aECQZj/PyJ
1g7jHlah4NojDtgPGdYomUZmMN5Tsam1qGmjtBC+cYzJaYd+qxlhkCezbYJ8WgMGUeLCWS/i2MXW
wjFSrcUJWMBGb2SCjpXHwMDYB4N4MwnuBHx0v/I4rK90OCP+edFCDlGnk09mFMVTAcXbLVwL3Fya
oERqeiIsIqTebrj0H7MgCPGQeWiLxN8pAY3D3o7BV3f0s/VtUvi0SurnmLzJrei60f5wMJIzOuXG
T/pPNpzoahJUq0AAAMZjIdPviBOjFdXkzcJIabI2W/KOhZQYi1vPfV0x+wqJ+1F46zsnfUxccXEP
uBq0H5OffD3VygU8mWr91ZEp6i9TLfQ2pcLx84aqvm+Uh/WId3c5UbgUtJ1K4PU0rEtEMQn1NzMH
goqPv2N0gC4iBC/lxySiz8Ikx+hWPrtKVL/bWsgWe8jBZWAeUBcNbtWJLNkKjnU7rAMNEohLKD99
NIoMvijBDCJ6tsTYYQe19MqnAc7tjvJt1iA03hvf2OqfvoagvCtgEa23En/5Ovwn+7tBMuH2KQHh
Bq7cWunbmk6/KrSDII9ylDXfDdAYWZYB7AJBfDDbuocbW22wKulo4MS84f3tL7Kgd1ZvSO4/kub2
xdLnjiVj02WvLJNA0G9u9byM4hsvDPcQcXsbgov+PWHnpLMXvRNAuH8AltaA0dpAFoknN+k7YiY5
vuRqoIHF8e+JyePqygbCvb4IREHfBxLZszZ/C2oakS2N17Xq8mrQR1pycYv1sNRhsmWnGGyJ39dy
9xInUP88mIePZxzAu1AhU9ItcReyuMriY57n48xGBFc2K3JS31bfSX6tQMeTLgmDDxtlVTDCQStf
5595nC23v/wYERMwhO+qFiHTTubypICnmYMGGUsWgI1/972/VSku/2Pm9EOiNFy3TfMC+iVWwXyw
a0xDvesqrmsoQ2iHO/GQDhSCKhfzAP2NlmEZ1iTun/i07hkMNHLQs9e9ubHaG3eU4N5g+rtkjMR8
6bvNUDCXxVAZsGktlla0gR5Lp8/lesQ67ZAEkhIfcgy/EGTixN2aS/8XOfZMCHF8kueRghft+5U7
8LhZX+3lJEBqOD/4x1c7Yi91DhgudjvaR2zln02KLWDP2NfxYwi0t3Yr3LpdyjsQPkrywn763wYI
rgeW8zmzjnXPa8pk3RXvJztzpUXARP2T6lKsgcmalVh6uDaKJwTPo/LwWo9YgcDJ6ot6snrwv2Lb
AWCGxiGsXtdAJsOOm7krIyYIAirMJMrk5uU+Hcc7sPIORAIZVKgGmuS2fQQu31PGX1EY1nxPpEYG
EkVnRijDyYTYDJm8YGJsEm77lifOuXzlkicuRW7l5mokdZSulEJ3QEuiSyr0IXoryFkXLkAKTwkv
b877BIa2LX3nt8QViCX2GDAlCghaOvezNf0Ut4lKnUmP+1l//I/w06t/noyU+VSpoIW4LJa+HZbl
dYUzr+mzm9Ren9Lsh19l2vVEUDxlbSQKDw+xGgrdusoEeyRtYijq3DyHGagkGW87Vb6xnbDmYor0
TwX3xVIHUHwVc91dLjMKrJn6vWFWLzKsunaaUeujSxVCaY1a0zxMKosC1kv0YoislQS4HScLXE1S
nIjRIjqzb7HpXtOb/XJwqg8y2Ao6/neUwGdNaYZYeyHMDCRRZm3i1ut9yFUsCbt9yXY1op2gEuiN
k2hATs4nZfKJmbibi1dSfTnRczDRkmpYYqVM01P4zUlJgNpm1m93krsrs/M97wcxJG7ps5HVWoWU
eGfnTK+2eFr4WVe+a07rvbnweKWYaJ1dwAAOg0LpotBVxtyoUmI/bQ0yv66aRWA7z4JWXVBNTgYG
rSWqHi/FxQ6enUnp0Voundr0NxuuiUuGcmoy3nsJJQmyP51oZsH83M6b6gMnO9Ac9+YpFEExLh40
8JqV+svA+YvrbLt8FUulwFJqqxCA0+/Rs3G8znRwWMPncJH20PIEpn6rHuhHXf1/E+stIU5WfJW8
X1OKRzpyWU3OT9WeLTnKVvOhZbcuYgDq0Y0zTJwEXxRS7iH5oysYCd2DBfWfrrEx8OcSnqlTNnUl
SBENGaQyEEVOn8sx+QTGnIJjZvXNHjFLv4/HbLmBLI09IciNu0PTXzkAFMTopbYIdGEYbEEQfKwq
Ue4E+L7j+TqZWyVrFJqEHoT4XdQtawAi8CzsOkEoKgkqIeQ0nTKl9u3RLQld106WTjUQprwi7WLV
0slB5kb7wV6W7Z+lQVq0sUswKtn61GVrRBtd63nH2YsvSr2YRbczHHfIjZ/S7vz3p3Isd2euoukn
kkyTTSVGvZzo3mq0DyoUj/wI006lAl2nrBluWo5hUELWq+z30t/31CdiPGYoWKw1ZBU+7YbQHRQe
/DrlAu88Sk7dgPFUSKcWZkVZQoGEJpERS1ueW38RkBQdqOuGxnTlELcv0R7UtDN+0ndq9ChrtxCp
7S1TbGL0bV5+3hqDpGLR65EYxAxq6kcOqGlvJkLjJ3lqLi34CicM46HHwFA45sw1ciQIKAuV3PbD
/Kpa+oHC7R6b5xlIh8/hJ6HPWXmcDLnD/yKzC/5sLTRo+yrl+tmD8oQYQx+Pa+mE/BRu6kXYSoh5
EDTmsJW+WKrvERMMQ3Wx4lc8l13j4i8swkqMsRVrdaBMwbAM1UriTK2RPD55ZUeWZkvShuROLOF4
IgwauWZRiXXiQLkIjoHkHmBFaIhd3J4mIV2bV7HOesxP++o+uJkAFWdhjxWAwUJZi0+6Tk+EkO7c
IBfMKpW5yizyAYHjDUZHBUxv9XmOPLPWSvDC0oCG9QNHy/29Ht0pdtlBV8PExZKXPSysZ7Y/fh2h
wXft8CQfv7h11F8W7wUUh0tm9pimHjAVKWq564jO1kNsWFlQPbbPob54goil0tl86+jT2Ket1tdG
lbU3YzaT2bnYkFXt063FEDMKShPU1hTMI2JAm/Mf3ZGFKZ6aSucS6IO3AKf6vHwxudX1dJCRtgHs
TKNEVLGucLN5ZWyMRM3ynZhC/yFCwauKHSqSNJAbkPGv8+NENXnVzbNL7rYoKMmEaYYekvHcR3q/
21CbqVXZ2Rs5H9pRsbaNt3kTxJZV/kry1Q3PcyqMxNdgeWm2DJFDSR+DQ3YDOiwfeC3PUhFGUuhq
WcQF458SqK6n6Tx6RdMu/PpZ+X5CJIdHgQjZXIfXYxgbcfV9IbZJ6uO6g3YCVSoeyRqSTWSjfsbw
6lEtiCQ18ZH1OZgh1EQlCmI2fqMpZBqYrdIlDR/EHbk8YnlDimVDRBqkIIWPMOm2WC0YEv5OzcOz
fpQSKiuEZMDgHV4xb3+4oXvV+mVAbVVhO+1CjH25c9keN7EEabSiadu//8T7h2k9EFg6nbXbOY80
xRrOzqgJfLSyawhN8L4b6vgEPyu4bDuhrSAoDJ/LGWU9B4mYkinRzYXVCTIUzKNLk3e5gCxrf71r
W/mNId7puu6ffEbcOebo+FEip7HKxfsXIG1i/AfuXRmZEF3ytnJXezt6S03Ue8fzPLlpb5LtWoUG
xlT/QJQk4PTL/2Yr71gX9qOSfn6yMcUOJoBtQknSzfonPRgls/j8n4TsaOcOnMcd/5VdbZhNafoB
aMeOyjus3+cmpuQJ5IY+KX3AsQPY2kg3McvcZC0mY3tbsPCXjMB4Vh1b7zgGnVswMsbviCRMFN7M
Nwyz0AbyoAjd5nLQLOjmoR3ihIAqBc/3J7ynPbUYYf5s72UW+oXBsq/N715IIvpYNDJt1/Slb2BJ
xsNoQApACblNWtfXQcx09hS+5Nm3P95dVkuFq8xY13eQR8fXSBo5Ef0zTDI4EjBrjKLN1bj/xXAi
U7FHw5hLaZnAyYLcQVlZ5pHqSS1KCwCWE7Ux934SPCo7I9DNqkcWW24Wb8S7vm0TNGfG5ayFBJlT
c8Fm4wSNMYma+Ix+ujv0zRubom6ttraYWDiD1a3N51Np+DqDCVzQe9ngF0JKMGz6CH5ktAqAgS80
fwQoAkh7X5VaWqtTp/I5t8Quatb80GKvCCLMsZGdwr9v2Pmaz9VTmsOSvnBHWa1vWcPej9N2jTgw
FCSpaKxH/QZaOMaeoyI9ECLuxGZ3pOfc7zxtIZEd4QUiYD+dk53WYj93WjBC80Ba515XLFef9gjW
bAiMWrRGPxGxmPdRuRx7TtybfHwmsO/8LPJWtDTQbwFLmO891eID9X5V13BGoJnZOQXTznulyxjW
n6UbJWzQTJZ73P0ykz/zenMlXHGjCXO6U6RqpfkGvAq9jvnUkthWCC+Dyym/lAojSbns0C/J0FJG
e2f2MQ+bbXV4GN0befgd/rLahY1YNxfCQON5x5hXuLkS+3DvtyoBYqoyTZvGBJ1GCoVDMuMPPoXi
vRwTLm5RwbuM5gjS2K+wvlKL8NTutN7ktT8naPfsFwhO1Xfmhl77mGx+ajdid1cF6W4ukhBtCEvi
CASqNXevn7p5TB+zMtyx7LgAedOExrvqLCWBTx90EmI/KAmfVdnpUTfjbotVxQHAYm5O5qvsiLEJ
cnrBBJArKgx2kOEzQ7gSc+i8ThC9Jv0zdvChN0dXhHPT3k2mly97QvcFN+UnOl/leUyvexqI/BES
zdkX4iuVmteW9nMpgc8VbtjwOFbDffVpWc9wjh66NHr8LbHD4MOISrMycot1f0fzot34+7ipIK4X
8bawGB5apLObmumAY66Tn4UPvx0zn3Jdo09Lx4d6n/6YOlwoRZFg2T/DE0dHKvLaKOz8lkFjG5Sa
1Tb433hIuOtxiP2m5nyD3v4oi/GZititRSNX0Ywp4wKy4nh/XeRzXaru25cUx8Cyp3oDusccZZtu
lbpfgTy/FQugEF1QcA7eDrXWiU5Ab49ArL9BnIH6SCsRt+aFNOhE0xc6QyjLsgxuGj6V09ZDMmfo
3of6JdK1ANwYzlgoexbL4jHwxDOoHRZ9Y3Rd9u/gQ6DLa7T+rJU5ZwJPNWoBSqHgIdys/jXycast
EG2ktz+/r1p3d99PXT06oP1YlJsX4hxr4yRj0YkyzWMzXzL5dB3Mx8kzhmeY+XpbkJ5oYH9RKIjN
S0lQbNFV1fc3ez9xxyL/sFcVrHojavd6LkJn7Z9OdacKtl4SSnWjpkLk6k4vO3eR200dwXCFY2EZ
nkeqy5xCXMNLbUiUv0rg6ZAvX5YUq1afYdv5zu9TLMuovikgW0t/flAJMttDBp853SIovhTCew4u
mFzCWbosAM1IP3MY4hI26bGjttgvJeHymYCmrOxakegZyP0roftyds3Ja3Dg4vzMrRjj5b93vKTy
J2yFcnbvm30+sD6DX7hoD89VYBTJ9UV55+D8pJRDvKIQUIUwx5IhHkVpm5CE1kBbHqUog1A/6vgS
Ksz7lAzLrYrvIfLEc2Q0B8Qa29zdfRbsJkEpWu9BrtE5BYPyg6Zxc8bV9wT66EHWTT4C4FhgDEi9
Hz3PrFht5v9GGrkjZjyDL/xrtA9qKbRtrKRNZ39jYfVrJRv18J6S4yH+eX1LQOiPNl6N7RvwXfUz
rFiRgQvJs+oGfq4XxcwbO1ab5NlxaH7814cdeB7JLFr5f9U+Vg8CFiwfMcq9xn9UZdAnGjVkCy7B
ex1Be+zXFTeqSgG/+JXk9pRq7kz9WqTWk9i/BIrMZeeKnkMkTeCC1njvUVWStfZzwI+tjtzQX/jC
rhCIfXTwGJYAvpPFt/vslNKVXnYX+xarUnHW0wPqa9J+wIXxYXJ8NqB0J0LlSUqgL4YK6c9ld/HK
Io8YJNm8a6xljRSwdUVCI9A6nGD2W//O1xa/epJP09kr23G3BTOnnUm8xSsEkGybKMqTeDR5uFP/
4gu4FR7u/Sk13skTecN6u6GbO492LdkBpUQ3X2T8ATvBbirxhMahhsz95IihUCOV/TWVFhsAgBUo
yMB67iUKRZu/YOS8L0Ut73D+Lzltx4JSDtywn86fQVsXgNmqQc5Bca/JjAkAV7OYpxrh6/U5ppNN
+N0Q2WiPAcvqXbZpYFTWvwLuXKoarjv2Xg781BHlmHTzzaVLjpxp5j/HWV5oL8XvCr0sZJo8oWFB
eVkjljY7txEttiodzF5lF6DgSJBjZ67YD7QDB511NPH670dGmVoLVF/FI/iY8o5zFtqZv5nRp2Sk
nt+P099wM3sEhUY01riUB/F4Voxh9ZTqb/9dA0WLZezG9hiL8VaDdTnEg9G1+S4TPYwwymZp3VL2
Y17ON37q7zUHbhl55KhG4n/K9YH4libcwQC5qo+LEZ7Uxbk6P1bXdNK38FyjjyD/724/VrqPWNdm
jvG/ecVf+TSmLXU8lkiryLoZmqAyvPBblL9WXGEUWVUU5RLP2Tdl2n7rRVdMI1AQD3mE6YYAXIO3
lk9mABx8Kz+CtnbODMrvsotWGbgPHEXbyQHFhYzZkNbzcVqf4Dvmrg6+d4Kt6X1j+sWpGyiYl8vj
0eft6jSmfgNSa2bGUehFesUEj9mxtlHLV3sAoSAxw6n+XpR4ZdcAep7Jj284GEJoxeKsBgEZH61y
TTePmy7+z/z26D0VqaAUTgCv4+i8Fmq3pV60Vdl48ID/VTy6wczA9xULTVt0/5jjmqtB5sM3u5ce
SZDnNt76NpEJg+6XYp1QEp33tLEg2CIJlXo/OVlXtiEDJ47HZaEhRiQbfIZ75UCzAKsUhW8gMCDT
GZEbkxDTngr+FbXE2D9LAGy9DGAC2RDzoSWwNnmVsplxYUBqczJbA63d3TrAM4RBiQJB32aKQYj5
1eEvxL8Y5d3SKS9PZYUA+9lrI6ZKw4+qn7JRwxqKu47min0xJkVlJOE7tWXs3BLbvrMJnToSEcMM
Hv+A2MhW9jFwDqJ34tbVZ80PncvC4oabj9DPL7qOzfqK34OQQd34pSkioZ0A0jroo41+yD9kFhNr
XezjBoCtdyEx+X0mO/Cm+1gzTfX1kixVHt5VhUfYqkHbNlcC+XtNCxz97BocL2zZT9SByaUM2rgd
z5Pyd0ryVsD4qgwIUxB9JYM1xfYL1UozP0NjyCjkKFXjRIyurs72aK2BBnPtCqUZK4UdC3Ivsgxm
HlJMFzPzDhx+a/oyeQhky67lHrCngAH7mQG3B+0t/5S1MCh+t7c1TgCDwro3XCak7T8L3bupiQIy
Bgoiwi8avF4Eu2oMuJ9gX5QkOssWOnCNgFekIaoiYs7ZqwQX7riyEL6E1ZN4DRxwY1/I8ZgpMfJn
blLEqeLkgvyMGo/5fqvp2w/LB/2HBg37HjbR79DGYgWBeUqNTgIGRPBj1tlPzipzAsyutsK+cBD/
Oa00fj1duhRzrHUVvFkk7MdZcqfp7bJSRwtME/TF8pkeyj5LZUhzpOxsI7O1caHYaLYoZM6ze2+z
Ai/IO3TltFox4KgDu+lWBq50oJA/UvkmNJFvBsCrk3CYtSJhCPSiRW/q2ubFOYn6NmEAT9G73epc
DB/U0zEfTuvKfdvvji8+d26h+rZst5Lys+Q+nqbcUkNEDMuNF03RIqpz2pay4jGt//Uxl1gmjpty
QwQQ4vhRNFV1VeP5FXmHIG4dgxzJIFqmYMauy9FzISpLnI8VI3fpPlrwHXxXCKfYPpCzUlAW46bK
DMJb8zhcB5YMg9cPnAE5G8b9j9Gj1UzIrIKuMNtofDI0Vc/6+WdNS+X5Z0ChmHleh30QYXTUrqrb
9tefZDMtm+7Xkrcd9gufTZhlSwso4qL+X6uqUV414Br4jenF5wqS57JAwyPVw2eZDL77qOb7dO2Y
M+gBK/eJOA8J5WMH0DT+GlH99kggi55BPHOA0w8gsSS6VCPm307lBfmKMHVlSnU3PLfoCNdrivAr
bthJnMND+pQTcuQJlyuRY0bH/XkVF4rh8MPeEUkb/ovEBSVPn5jg4SXvICvm1pocUOjRcW9PuXN9
zgIBvSpz7AXobd2H5J0Cb1oPlwUef73eNAACkl3bb3TdwFEcxLmJXQCtLEj+XzReLKO93zSBsLHT
M9cEd1iHMmlvUynmh3PExclAuFjn1ed5JqLRTz7ICGXNYBvviQ31WGKL6hoEPMJj+5g3Zz7W9f1B
9f+KUPFylRHa2JbCEJiBYgBL2Hs/MoXdzkbqiomizcI7P+zqUNsq9euBPB4wVgPiIgTX5V/1anGB
4i5OgL5HuvFyaxzYT767tbRfDUoqFnA+LMltvImjrjKLPsV6qE2JpL//25oMHemuSe1rG0wKkWOg
r3nw8jwApG+ZvUoNCmv0mPo2S3nSIfjO59Uzb7k3R5yI6y36+wXHDJtDyFMhWpI6TH6BTMCXE8Hg
IfSNcGIIXGtOPy/ZLjtiUo5enFIuavzIIhmFpRpXo8idSiMqFVpsea2o7boZJAJhS/sw8OXcDQgZ
db7kBeqfwtJbto3LQyGaFap+h3Pjv3xivKB77P/GH+9B7KwUgo0vrIYhQ3bl2t6dkqExNBAlFrql
aflDyvZWnIYcGw2dqaqdCA7JubvKs6BsHSoHFReFdHPaf9WcxRgYnQ8K49kObxUj5br+DHbCdVeD
aVcxp5fjkFD4TXd5iWv4AGr2CEQ2b9rz29sD5UJJrsj0uuvAhIe4yQsvifcNr6X8dfBiUSi2QHFj
TtT9OZW8O4WwY+IGrS1Q2rdp5zUzwehZa+MkvEr3LzOwYEPRlpTu6Mj5YVsL7m8mZVr1DvVfgRK5
sbbYjmRryf3mcitUAXEyX74IZme9C7gCejxkxKLyCne6y27nm4R0hCQzu3DiwPKH9grrYkmIwfNq
mLH0npG2cF7yrDWgatn8wTMKNw0/sMTtZbdDBWp9dk8bn2gYxa8gI/Q6A+rmi5WvG2f9udwWT5CG
RdhxO7UVlLRiH2/NgAU2N/Wk/kKnNvQHaT/3G1MZgaCgTdkapCT6jvetvY9ZVDny8eAZwF3TX4mZ
SzK9H2SlkFkfA5cuASXf3W8RD31PWS5UD0OY9Cl+es3TPQqWQE3zt1Dtz2Wq/IKzF/m8ncFIk9YJ
LoALCVYx03JQHVyY8Vh1ORwDuP2rujQk/ZR5wOh9TiIIW4ejfQ5wF9FI36Twcgy1aFbz+o8q/gh8
nNwVGpwOsat7v2HDfvw/Rehvo4l0dLXfmcbTHtplaxcMGeyO0dCO2n882nRQtoAFC9fII1WMLhp/
a/XNYCPO0XXGPQWBraH7FGIrnsd6VvysDtUXsO5jUsNdILtutntvtvxhBPey56+NYtSAUL/IE6Xm
sH71d9h/uFFQ1E4ANFVL6FmZSx6QPJTN+My3jFeLxp5I/sJ0/Kn7htZA6oEfU4zNLJDk45UkCPRO
2YBQaZpVo0wN3J4Hsrp+zUk+tR+Z5yqi0xmuXTCM/PwMTNceTiwWlAyXf4WB7JEXttFt5MMly9uh
dvzOaR6x1WqkMmEblrrX7MQ/+LfUTuqnxaVWR5zAHc/b5CktxD2CqyyTmg4q3apbWRh375Y1DHL4
+lfodwoZ8ZusTkLK7ViYj1IX7UItIZnZSMt5fTo26Y/nkNefIJnDnzq0VM8f5n1wyAyGC0C26oZJ
dDfkGrgr4axgueGiEDrYxAgGbuXWXi4nXXYEoF8D3aPu8UJjimCQ2p9qbV3t0APLkvkhO/Vdaaxi
nYQk0U175FqerCK+uTjt+C+jfN0hDtNeoD+NJoGmFiQeajqF+zf5sCRg2YVKQixdcPHk/MoWD/+P
k+Hu7SSdwWOVDjUhsLDWyFifiA6NqJyNo5TOXvm11dclymE6jZPnz86DBPRYAWIpgf3NjVzqe7Mt
TGiN9SGqEtWY+DzHq4GcZ3mCC4wEx35FHRbspZ+zkdqgidwZSY1NDPlHSpuz3dkfrL2qHM2zRaIP
27GIxSUzJrQlumb+EbMv/QYMQ+UTXOyFrwotXAHQ2/Ri/FRyXdtTacFQG7wSnmWbGLwaygISF284
JaJkv/YrfxntdjKqZmHAgqD9AFv0nNQXV3iMSO1mrVjV6jovg0MaAWyafcv6Gj9LsBDJCKKuh9M1
nPz15zx3DprBoZBtnxNIR1BmuPfugAQHqjKvhvaGmJoOovHACrUHWYqfh4pXXEvfvj7lT92yXdZE
VHGE/geUbcR5t/E2RmBbTwl1DJXuZlr8zafISn1EPu6BBl6z/w5RUlG96LGgbMj3ZinLlJBi1E5G
RmOFCKzkalAY+/DUWw+xpPWA5KV6hH03uMimB0X04g/zEs0xPnLt6tceWRUd20faNCPaj6gNjstN
8yv2IgAAxKGmGRILRUhCbFKAzCeVqaq8TUzXCOnkVA+FXOXYPJnKE8+9NrW6GSWKvHjJ1J6krBio
s3ZJyrwWNcwWDTsVTmmA3FpXduPgeTprz/5A4jziSwvzL2UddEfb96pN43vUeQeX0eurbbSlfEIr
Hw2qAUYuMScrV2xnCvdGATY7UoxNH9ozQzflAP4/E5FDZgraTkXnDCMMWIXz9RA0V7YNKpunPYc+
46+X3VdFO8WuT0FIVtBOXzFvH2+VwSo5IeM0Q6LaY6QpvSETXjUrsDeRbZigrIlCDw4aDHRelosa
fyHRQX3XXLY4BxMNzpDSueig8ILWJQtAPTkRTzmqwHYkncnb5qlVX+Dpz+GxTj1GpzWokIwKV8gJ
0HuufF7ar3QKTwklR3uggLAAOb4oub7IL5qiYjyAzrgPEvN+oeDEoxuDvcJC7gpd6Jzun/LCillL
mClM2n7p2E1OjEBS+TmRFCylnHIYSl9w6r4KoBd10NLs3ihR917RmkIP1fAHAyYstebWMJNIAAqW
WUmjvFNCan8M8HBAzuuE+PqRbtmK0gx1WgH0OniBfg+Jtc2xl39DzoMvNxobAT2R+sK0wUMom81O
EjOM+gKKCu5rIKMIMXRoSMs48+OyqOCdmH+W3V/tNmV1sWAI7IE4sk1ciLYihVY5K+2NLBR0EO2F
b/Ckv2KfZtqxE+Oq9MN7MfjrbPdGFjk2S0Os9pA/o6Tsw9IxeHKsr1Z5pF7JsZCYvBALcDu9L7uR
ycGSEj13nmlHS3BHWfSRJIETuLy3LzpDWgp5oCLNIuYMSgyfu/vlfcAEQZZVjbrJF598QupRZihI
Eq2ol+8jW6PgEsZUbC7GKbMp7zq/wBStkrUVIQP8XeMx5TUIo2iqy68XFS8YEhTNmgxDQJBxlif+
XYFw3Z5aw0QisFNcoQMlnmOkSfUXvjr+nRsPoYLIjDeK947EZ4p3smNcw54LGpjLgAlhLtsxjCzT
q3DDWqpkoB2V+eFROpewegxJ7pdUvKfZGqGJPWbfsfkpn3QXatDhexi4V/SuJMqhl4pyUKeDnGwP
30MSXxXK0g+JDzVRoLejFuAYvmgGDHfvTA83/TVqSA41cv8iK+uNay14lZkIb4TXNUznAjRnzLEL
LnEAVmRE19cMN7BN9Ctip6X1iZWu8MSFHCZ5GxQiAIux1AgufA7HpJu/ZIKoG39HlCsHyV669UQ/
7eOLR3HaauvorbdfORtlxEyrpAjhEGdgcR/wxf4yfl53JHjtbm79ELV2ZSlJiDnhIce9wNa5Fpag
4iuw2EvBWfbBKwuD9DfqbyUhTLHu3KI56IivbFHegYRmBbrd+5oAV0OeQrCtM9VPakn/xcaHUnDZ
4Uk+BWUYjWNXXx3X70wUWrw91U373JW49OwrTYb8SeFZIECXxu/YQgytgOe/SX5pZbbr/RhNhkzq
DVXu9GuCxRFQlCdeJ9fQhuz6rCllrwL/O1Q6ZGts7QK4BEOy6WWgQFvqVtp7GI1eeC6E9NLpoo7/
pwpmdp3eTS+Vu2J5vkfaVlVivrDkmvsVN521/IYe4rxRmotbif36e/HDsCJWV58m1Vb+u2uLRKYn
dyMqrtB5DNo8aBpTlnwwIUF0o4jtXE3qxFgSs7MZLbHkLMJgVfTlPht01B0buK0ceSsmIeXBZbzG
DuNd6cSyml0fvahh+u6k3Khs/xStdTJVDzj4Yx9yFj5h77Eh8UTMAh7g8ERbT+WQrwxHxVx12FwQ
0pZIpoRwRjp751dDbJfKqtGmkL2aS8OCCVyrbTFgOL/pTeYbdA9a2uXyNMrtn8XtZc1tQCjWnpwm
7kzuMNjQvQZkI79HFT5+66FkPvXO6mML66+Jj5EAbRPkjVn5VNwNGTMJxCMbnJw2zmRgAqdFb4ly
BpQfNnNCPy3jUm67Kpi/QTYI7T9BSNOh+RJ41eSY4LIiArDZ4G+Hw7kEZv5klrn3iCg362w5k/yQ
GU1esOQfD+J5qodVlrgsiZgjr5g2Ah3qsH21bJXr7atW7BevRQQm8RTuh5UCITbCKNCEwvmGYqkX
16UL/iTsO8ADny9GE2vwEbguSr6pPGAmIhkAKjxD8bTUD85SUkyYy6W4m/lH8q132tDlV/OdoDlJ
1KkXR2LDNF1v1fPKV2HPcOCevAUnFsSPjD8GnznR4eOo5y+2mittgCCoKBXhqSKWNOQcDD6G+0pa
H/WT8yYoHKgq2hm/r54VanaFQRiWGVyqKtIHYaj+LOfulBUjgbkYX5ggNqbcuFofsqGyYK+rSnQ8
TVG8+41avFGaA7Ygkaiwy6XHUFXyQiR02GyLYesHNBoEiu3FWV3D1578X2rf2PIPDN5CdP4g7Hpf
1T1Nwxp+jmjSRQEvTA2SPhBc7VjgStRF2awbztBhh/RIxOyKJsXkUflFz+UQke6p+BIYQjzuaarI
2iE2XmsASxvKM0wZGb9aqFR7AHhEZYQ/OL/9UUxKmbm+u2jHieuaB+LsxJvHYozQ+2WEHLS7NvPy
ffVRPRrMPZyqNO62TDmVxeAcQR/cXPEIl/L/9l1gnzKjdpLL6B4O+gW7X49/yAHrFFpcV/d0QV32
X2FEa8T4RxHTvArSCZFSROTJsp+mRStgW3ZsFQDKypEduzZO2jhOCJxAa9eBJPK5l8T6jse+oMvJ
3ReTh0o8/jUQP0j2Ol9TaihTZrXS3KBV56XTl+J+0lU6EXdQbOKlkjZBZlJSs9esaXsRTWuDQPpe
KQE+eKbn1Dy+FZVQwvU4j0482XdZ94gRgehO/zKHyi9WrbcKRoT2F6Oy0KtK89UO4AuubH4DHyR3
5TZieKq6iW3Snevx2X+BD6QmEHU8Sm6FtcuB31B38uh+MUXIQ6eHJX2ph99rjnFoBEM5/W1G/Vsz
Wi/XFuSnvx++g0Mv8NH9Yfu3FXf+X6oGHsPZTd/vvXT2tDQlpD4Hhw3D2a5+4po8QJM2fv27NPAX
Nd+XwjtxIfN/QxdYFg7qKH9IiftesBIeCj71UJvqKGkD3P6TXthBactzhAfCI2DaTDetPjQVzSUe
ceO1HAlRSim4zEMQYE26tYFUSxcLf5/PurUJ3L1icNGaeQZb/PcWEM3w+0FRSPATLNqPxQPeK9Pp
FzQBc9gmrXsskCykL6YjUGLaTosGbdHeKl+B8RFkIycvlIWJitjQ0PfHrgbyUU0I7tlygHyUZyoE
XK673dkncmrOq24JH3IrxPMNwA5KnVTd3vaJC5yghOWtFqX208Unuu3/PD2LXvCxBe7OCm3CJ7Lp
kZRvQD/JEutliBU9sGue5wMzQ1hEwFCZ6qbxiCQ3SIrTSOdPAakKZcvIXa6BAWrUz6WtjnECRfGR
VadFx/539F1IliLYx3NA2IyTd5cJ+Z+uoY231RA5oKlPTJqI573CusgVJWAqGJ5XfY185PeBilWB
Oe7anbyVekli0pa1a2OsrvwgqPkrh3BWm/292a7SpCEbzKhpFteWfsGPoh0CDph0oMv4Fwxcgjmr
JZYv+3c9TLpuA/wruxjjtO35ySEHjWFVk5qcO60JLijyjLmSbI86ZZlUxZ4d4rxuPmwDrVU0YXpf
uMtq+vlduinMehwTzM6tD5Wp8GQU5KmtTJx9EVUim+mYSt5YpRVMbJA2VOalmACS9d01ayde+PJ+
fif2MPtKfkOFyI9jLGKv1ImtYq4+v1oDcVJrQA+mhfNo+MLt9Ty6mclSMWI1AmMp4LJzAnu56Kmf
XOy/N8LbhgTE6aDr662UOw9MRyctsbAx7vOmiSbHoIAYIo1GC37mDz5G+UOx2hxA+D/UfazaFsC+
Wec8RO2+ID4yYVgXL2uHq6g3IZpTv+MXDwR+3P9bgVE1HJVo6Y8DnfpM+jhdvhM6PrxXk6vPS7gq
owZbc1Y6Iw3gtEpPw5pmrK06c9oYT65WIcU3onKs47vuuaQY2EIKG+zZhunE1MrdoJBhWrmdaA2r
8Ldpfiv7HdR+d9MbCvxk8OciopXvSIsEVjIBcKx/3xf3x+tWda/1jEZ8qhYyiZpXREc7dNr5VB+z
2XapavwMKVd4eORFNWGfOQVUo5+VVdL9JNjFv0xGg6G0+0wuEzmSH83L8UfWZAuqsa8xrBtEjxMH
K6ysOxa39WY4kPTTW+hKQ/JkqfmmMTzPcig/5iH39NOhUvm4ip6VCOauDDVbz+bYTKjKP2JVuVdd
6L7aUpf08Ny1FVMuP7wXKty7dlf5e7IZebuFwo5R0P6zy8/BHuJBAl/q9j0L95vQLdDqfTgbKQDo
4uUvMgiQIn6ubyb6E2vWsmjVd58UZlygtsNuuY1zPcrGxXDvyCzQ8ckebhMHRHX8+15WBKYVGcwe
/WGa2dMbvnv3EqU0y8EmNERQ3FdMHev/pJ0jE6rjbvwB55FyFTQ5PLqfyxHR/b18AcrykoLEgaoq
ko4rp+H+dtCV+lhyjydJoW5OxcbqJXsydt/rOfVCyOQ0fXeSBeo9Z0RKodw7vUN4/rX5I7U3ZYS9
tCZfuMgsVTEyFfyER/v8rx3dzhfH3yw1N3VLl3u8zxCIkUPao6LeRucRndVMWFtD8i9ZwP1JwHOY
m9LdT2BhT8mDy5zzoKSzQe7m3Mtz0Ebgiu9hoLYD1HNx486lmqUqdKdftjGt5v05D8VhCx/ab8in
nVv1F3f8SIZjnTLbK5Uqz0I5zDDjFvvHFevQ4s/pemaeqjj4zw0p/6otLBdAUo+eOnaPoQrEZnjm
RVCFvmNuff01UEmO9i5p2Jub4qfehZ7Dqr7f0cloK0gWlcVHgU9t/wWWk7xZA8Q5crafaTq/aeM3
aAqCthtg1EF6YvqwqwkuwnI0YJR2983+PMrC2NG8+pKnSwyhCG6tmhjnF3+RCP6bYLjXLnHj5VFg
8dn7wG4UBvMAE3l4MNgTya9VOFtP/MQiW1EzHIgZucvSXh7+Y6PgqohJpy3/kCzEZh8KGO0P678P
DflU7xSV/v1cV9mHj2q2tOQpLpGmScl1yI9wMagZM0uc7FljtUFYhC969Du5Nsu3OwzxTAZ/nIFT
MHDOLETewS3tWT88buiM0Yl6Q2lQg5ZnsyFe2JjYFJKYBPftxuWvv+XZH5+sHlcMtxIl50/zW9ur
z33GzhgioKT9YWTMKw6/8h565A85soyB0rncZ/onlTwEjzgBjZXivaHg00IpshmATgIV2gtNjwtH
cTBrrXGoxttRn9jdgyX7Ry88AffYi9veQgoe5gsPwTIh61fVaRrRnxZzevU+oIwkatl/vUVrPWSY
FkPq8lUVl7koxYc55aUEK2+S1SIeCQbVj5ci4EmMkN0imK3Nk9HwWv/4N5+0uAOcJTIHW9tGcsSG
QCPMz2kDXzbHsuQ0fcbeetY1syPKYSnJb5iqrm+dyid/lV0EAnV/xqOI9jnEoJ4G6iNB5iifuyaB
kjevIWSd3GBv80BcY1+kDir+rdKPKafy2ynimLNED6YW0Dmxp76Nf4o7hVfGI5yiAXHEc1VvFnRP
CjRQGutr6YMatgYwTbV+uvL3fBohQeE5tNYZMLZJclfQRmudupADFCjgbKw8EJ2Z83zvW88Qa/v5
YDZ9plYMc4pcmAsahVW89gtxs6n0VtDVMdKytk1brQPDPwcdH3jHARnvSMxGY4pQPWZ2Y4qaQHEb
qnzqpIoFvsEybUZ23jozHdd5Osjuus97K4T7w9fQ6nX9HSBYw0ncQuMdNlzuLpwkKghJScF6eMqx
mXkYnjTOn9n+jn3l31uYbybJdyU8lGIFOGtjk8TjDk7lY2xMTG/2xJly6TgkrS+IA91CGTGVX9ol
s0EVvwF001wEFt1Wj76XWWL5GSLsiXtUXJjxFPWVDfGZwZSy+3ssGk28pgWe/LKOIbUu+1ZGW9hJ
FQ4IkMJi42xsI7MFB5rp1XzKCaPJECaFd8JO/U+o9T60+J4CVl620mON63zqQgxa46dyoPGnTC+I
jzuxj1hW9EBqJfM8PIsUPFmdz/VAEqOQYB9hEIWVE1IP9W1NGYLaylG4XZJhf9R8yTlXGFR1IePr
uSQ+pzxxG4rhKn2S+zIvVRZgZsHPLva7CO3sBivl9WFOV5qM6+SBiOqm+JK9OoohlvLQfEekuCxk
OWxites97h63WTaVxl+WNjLoynv7GMeO3MRIeV9cIBT5e37HvIjRFBgzXO1EpOMQY57cst/9i8xl
cxv//QZaEyZAYGn1mXljqts/f5VCFwReMkxrHZJ3sgMfVzaTHSLxF6+Mk1M92UrsiVomBEhQiyag
7ZaKFeMLW9FCr1dBqGfYg5IpjbUfBk0q24VXjOA9pmJ8pf0+gOeO47KJ3Tb+QaNb3tK3V18l5iYS
IE50DtgaIahu93gqBunsHgec8o+iypXcsXyAL+yCM/bnYVfwA/K30TyFK+UdYqo3UAiBPMNQFdm/
f52GkVZ6nyLvLbQs6EaQuNtpTncIh508v66f4eFDWjFzsMbypovPDjetHiso0goFqysppUjetfkA
ghOtk+ed+MrN1mNT0MxW54xzZ9N1Nxpi/70pB1GKCQW248m6ztOwNpEkK9fOJ40QBPCpP/XYpRXl
btAoGz/2QZLjMxCvNzh+PrMny7k/CaAUcsNXHo8VHLM2vESzQAMIllVg5VELZAq/9rh1dnL0L6aJ
DeIa9yln5Rdt81sz427/TKpqIB5/9WX/CRUDlVdmvSVDBTc/CFROvHnmQiij8Dd4EkjZkTw1Otvv
FY5ji94dYlpWiQUQCWhCgVmM5HrOiih8VjhcbXw+b6YZMle8cDpio0uYUFSMT3AhmY/is5MurYfo
vgsHxaCkng8wr8y9FDMkgvEvrK3Yd0gJjz4vA2uoyguFN0PhDHgbzILUHlnzEdpFrXAFWBrC5M9g
7sorcrl89w9J6s7NuWwqaXBP752kGwHwCQX8t3oXN7YOUjvBjxBZHeFuBNlZTT4Ro3ZOXLGFPWgF
kjwsHJtXTS9y+HirsQbW7F/ARUgnO61IHImtDX1EDXDTEpMqBnDGiU4s7GR3YHT0ZKC/HZCbjT55
qqRP5CzHb1vqLp31Ied91yJbnhUJLn5OdYjwb3SGAQV+9OMSdKVuk3E8u9S7zvl3Enah3PKoGE6+
A5tDYqltQv+980J8aAbNnyP3JzoKNl8FzX1MfW2YtLP6Fp5vNAyhSyfYyZ13+3015DGL28mwNs1e
hY0T4odUx8ukhMkOTt1ItQ1AZBIqErLwWwbUdnox5rEbfPx1fkm2L3+6W26i7uLl/jIhqTTYSGeh
vMWqZzKn4WgrGJB/ipxc1R1KoIa1uwhdLv+yz15rDUWdON3N+uY+pIg8gEQZSYWOupmUFWrLbJPN
gxP3u7QfI1dEiHDwKZQM4hctvOP6igWO3A7IN6KPZ5Fjz2pZA300737vVxww0zt83NG9UoIyooF5
pGiMEFJA81GZXExGIXGyDaCGTu5RRv4733s41A7stsZ588GCk5A+nWTW8d3KRSD33mLA6T9pohMX
+CR3LgvcrM0jVHf0exR7AIhR/NlbytyCHIojYV6WnHrkzYxeppj/oplvq1FHbYOzPNOJIoVSH5Ss
ILR54MbXCoSUjgYtIbTZegSOwVgKlGchgZIEBVrqksyOmHIbCpYwv/25pi9/UglSqJiXE6UwZT5h
HsFHxaMpC1CgHMqOCR6YTUDB8iJw/NO/1klnJK71ougCAm5lLh+aZqW8IFtsD0Za85kf1d6oUhKH
a3m5Hg9yCxXe0XtpOy2D+cI2uq0MZaQyhA7XeSVlLslQKy8/ouZMWEQkipYJ5ArFZResXUqDpPRQ
pRqJQzvwEwK+0cbdZyXFfkclmzcsCo9+6DKPVrrGfnw38YH8T6326Ndwd7x1TsOIBpsTT6Md9Dch
vowm3UYdnbxj1G7ssqPBl2CQK/FMI1o5Ahmsv08M8Q+o8BBCqcA8yQNcOGNuhXjyRmeYxky8JiI5
JLXnuqLFCgliJh5I7uubJnGD4XnVAoBG7892LsU00neowbM2ogc5pmTG2g1gjGpYmTqZUsXilT2x
9G1sSg5tq1zTSd3h8IQBBAhWsmAQ+2fsSz+NbWRAn8MqylEm8rjlII5IE3AzwWc76XFiTMHgNFR6
mPxB+/CF2pff+wE4JRz+HEqQf6nHNBSmIsrWnL//pWm6bVgQByR+cI58tcFxU4NSKGDEUwTT2pgk
aaNHIPdyNQ+pIZHrwL+jXVUjKyW1M8IcqEKaroC8e05M3YqvRDfn7YvgkAavbf6IX6g0xFpntZeq
aB/jECRZAO2/wtZje8IT1QTOMsihFEl3DDy9DnBOYOYffFW45yJKQxdTxCd6i5l7DhoZZweAt07t
EcRCi9WjhRG4/jn/VK/zTG6ovRk9DFW3fBe1461v0hEWaHuQJRfX7tNxavBHhNW+07MH/7yBr9Ig
YjT0s70HWXM5Lza75FrLHK/QJVv3QYjLFb2QG49CkGFuFfJ3rucLirclz1+H1NvyPRYggwGsutdF
jC0PkjOndf04D6MrFTPpA7zWgVJE/MI2N8uO8vrEagu079Tv103mgTjibo+Sv/HLQZUt8ifZAHJe
4jRSmCU83LiI7N9OOuemxvnr9pi5baF6ALX8ut9skOk3fR0pTWME7zQXVZ0HO5bGOGLIEYwfRVrI
U72fGsKHYl//iKRNh3auKQX3pq2BzZToWmZLu240Hg4pAe5AMLKpiiaqXe7zPO2s9W+yyCu4os4l
CLzOfRoKqqgFrYFHqm17GxhjE4a8IYzo4LbVxL0tNNRJ4UMA8pO3ybrecJl1HfwtwI9npP8xrCiK
DTpJ7Uit04BXewH+OVZaYb54cdTHV6LZShl747r6w+VIC9cYMx2NKIXQ/w/Oy+Kp+qZ8l4VUBgZU
wdNIsc0R93/wdOR68z8peuJ3jkOyU3U+gT2bDbs+90YWpLKB0m1X8BxsU8C4TItAppDasgaUWt+A
Gn6oL3ygeWTXTEHbGs0Jr/PMi/9xXk+7D8RjZX6MUmCd1X1jKSJejQFVa+LZiOacHJdVI2Pzz3yh
fnDhQ59W2gXtHXjuhpKVcHxFt7mhwagj1INq8wZcq0BW5nn2admT2l6eH/gOkCubvKxIIm+dY1Vn
jCQQAkJSAkoQ/G/j8Vp28w1iqzbMf6mAGIbvbUWLtih/1iVRccrCPQv4nUVA4KHinX1UbEdNg40G
vGoboMZ9CSIFVz6IW4cnskb3x8+SGwx/G2khZO8WYBMkEAIO1hCU2Cyc+Jwwj3ywB2Wylr1MJFPl
+mZaY2TrLUWEI46VY0Qh6DeDv9B3rdyqd9SijF4YYEexlWG2i5Oi0Gy8wO8EWdQSplb2J7bRKB26
jD+rpmVYlV+kw27UDri4nJYYQ6hniTNwGaGkAqUt/9jtJt0HiNBNBAujMYZ2VFj+/LH8UGyhFQ3Y
77BL1cnCForaA8uaFlncZ9xX4ij5D4iTkUCraXaTXi2mAixSjwU1jqKjH/jeujjBifaupPQzXvsP
+EImkOc6iTE+C6ljLQG+BPglzigoF32Q3JgBGiJceHUbxkgsNgKbU0u0bjMXd5WIw/NKTukTB4zb
oqtEIv286202LqV1AbYU4RrhACaH5nuJtHxwhqtpxYPoU9usQtryXWaWZvkySzlbg4F/XAWsZVeg
CPcRQNZfCUrAAeTK3z9s0z8caPUfxggueL7V6zGW0jzB8hasonHzk/pf2nwUU5b9cQDqLuZNqJmo
7WUD59XahdX4W4STVgg1n9MQfTykSkPQOg1BHcbfcjHQn5dTDL/y57T+umnEfuNJwViG+agxXp5v
remsD+VMM5w2V3mdmecKZ/Wf9Y97qO2lxgony2WhLPk2ePGO3Y2KpU1hCx1ihS91/KeQ/HmnmAMI
3r4j82eO5yWeC0+8YFl0nuA79Radr9LfdWZIYiqpj4g/LSJ1i20xZV0REj2S2UCWgqafFugWpxma
DdCS2vhEUmw5Twq1dKxxTffA8Tk/+v0KUbBdPjqCsmUxRatfk2q66lMCfI8Ejhcew1GjLDZB1ckL
QvNIpEaOOWNbhvoiEbIh1iDudgC+gelLP7FJV4gOpRKipReRC3ppbxrBiu/AzYKazCKVj7dZYZqR
hUbOA74D2mkY/fhXQ01fCoMt72sYIcGjOAMLelBsOYi9RbIejA6yrf03Vr/fGo34l5eKoF+Q0qwd
mlWB5+0T3xoJYXhZyoqg2goFtK1ZphN4nlwrLip/u/CuxiYPUR+qCjDPhZr22uj4coAOCJf3pEyQ
JVXlUqincnCPZAP/3o/2uIi4Vc3ct1GyS5Ao5OqDXA885lC4dPg8L1tiXJ6IEJWoiRDbuLWPWANb
Vkd0x4X5h40F9EcXFBsXY2N39B6Txtu5KyA2hP+F0mn119R53O9QkgZTSRGApvriUum10hnJ70ti
NkTtjaD6X45oNqGmtFXDIe56ypzpKerrs2IEm7eY0NjfZ3uC/AOL/NnWvL15Lsxj6NAyGLjCND//
28G2BSnvtynQ/8LhwKaX8rwyNdSvs0nnf1umt1fPJ2i2DRIhbywrNZCcgBwgmnsCLBia6gt7Wznm
AAD8ijXy8aAX+qXroUiQdcgHVA6I8os/fzM+MPnhCPf5+Cz9PEGY6TIBf0LVpXUVDDg7GOX5B3h/
0cHyYyK4pn0sVipMyPE3mf7fXEeOZNVMC3hxk8aJoc4hXUwfUOl7FqJ94jhjSmuMO+CJhv1J62KE
9sovL0YVYwICx4VaKcNyupy5+Z06LbbglPOmMV9cLD3xhjm3MvD3dAQPH8nYlzt7Dsji7mqowMyn
tWVNI5ispEKgtPxVQK8arKYLz4jqQVRFZl9VJfbx5Pi7VzMqfDXXjcqA93OCji0IaWVCNhV8xBi8
s/GdEe9oHjGE3eQnmcfcSTTyZuNXvA5ikThbocDyv1if1cPfI5BTSTTTjybxQFpN1gaBd8PVNUOM
24/N1yQmaUTAYmE+wWdTpTs+HDGG+O9DuEcGsj3kaD8oedHwRVmRcXfp7c/vqmhQTTzCd9n+K91e
s1sro2qCMXNTMWqOK4vbmTGkcAyqftdJbdGOSt2IO6IbknwEHeh9pjo2N263Sv4t1eI+lHgzEe5K
jzGI5Nd/QKjP5wX/EBe3/diYiy5MCRZRDMXj5Pos6OGZ5glyN1MOQXdZRmm9CkELT4k1ocbTmOgo
2uTJCYOVH+YXmA9wkMPb1hScAcu5BjCp3R5+4rLnBoSYOfVVw6AbHDgGPJDEGy5ViACdCCH70H4z
xqlge+AvyRFy1UcXBCuAyDQ54PKqxQvQTpnA0KP4k88Vh2tErOgOKOdKZxIeWsUYDMYPMYCFFGBW
NwLK5zoL+yHoQKMVbvaFHZNjN2m57INT/ofYjN1+podvF5o65cVzR+gFgZgdi4t+ibx5NrJ2oz5C
fh6m4b1nIK5TroWxR6ovBsFqOqQPDDwJnrLf2gidxdAMPIQs0MoCQ23EYo4IlOW8wwMQdc2Sf7pe
9asTs8EWNP/z2r/o1lP6Xi54FfUKpRw2FWQliQ+TB0+HbV+5tCljSKxHjEfyN9f+tlRpocu6PtuV
eRtP/9N2IEq7rxxoNB3Aqzlzb99k3mKPqYOVTj52YBLCUCxQQALSAIoIfwJPa85ujAd3bCdmyINf
9QrjwRYCqvsaRR3/bboP0g289MvZlfgbPAH97v1qwVPA5AiM69Eph2zIY0s0WkCY/dw+0xVnjnGX
MI2b3FzsfTHMqch/tLQBAr/dUTt6xzoeFX8CwLQWxJNNyNGln31MP2CcOLk7jAikAN81CUY85Ld9
7xVFDadU/nPxvTE4ouYIw59OJ/dVr17klhGjjOvUCpP5dY7rcBM/qdeL0YYEAndxv78gZ4z13E15
F1T3mYqrHqEWpxyP25X26Whq1azXM7nQUQS6JE1jSBnLYMNfrftvFkkXb2JTtKCf9HadZajEgY9p
mvfrfCXhR3DJAFYDuJ7J1qXCM1c2XWiENTqwTIPY2uQPcHAoauDtN88q2s7FdLwoZfD+i1nbZVAS
WI5YbY95o54JkqFmUhNAtIgXSQepHPRpVXJKHR4jBcG7oDmpLbuzjTwkXg2bN1eom2u0xUQT7Rrz
BP+zWqaMPJ83DfF2j3vd/bx6ACGDtqS4YIQiV2QS9iekemb+govurnz4p/fSNk5RiqBvA0zjCO9X
gPST7EW+r5n5Sx86MmCGDrINvToUZF+1OCAwfQhwz6RHbffUtXl+NFtwOgBblDJCwOz+nciFIAKd
s3EeoESXFVogPwJwfHuTu/ruj+VwZH1nB6o7/lnA/AKuBbDWNDa8pqoy2mfl962E9VV/NjqmjZuE
qJ65qFV6TnBamfTyJt1F7ilVo83CzKxVcXCr++7frhwm9s97aChAWZE7Ay70xf45Tiht1YC92UgB
HTrR4e8aF7wdlLfL1VnWoBahJLt/gMc4pajK2KVHSOsiMyW0T6HVAivb7nSTaemYilUT0Xo4b3Yc
gAnLRAatVoSDDW+dmsAFvZzLqgMbHmlFORthkDKkQ4d8D0WsKHNItqfIXk2hVJHPXhHiISC2zvE3
XdL4EQYf+X0+0GNIqVapykDc3DMYwSf/YjCwCwmDcisyGGLMVhqwyyNEHAzfIn/Gn9y77jm06mPb
+17fPaxI3N6OR1oMqkqBJw9hEdoCmL8/avSVnoHL2oQZZr/mZ1yS5LKMbSkZRVpibC7jX64ZjXuM
fI7xPDBLHF62FPlmIF2pwCVLiV5OLWybWz5v+Az0vryP5t0EEIIwu9H3NznCkGjpM2Y61d7c1mn1
roSVbB4liJonfSFKGUai9FkedjkGuK3a2aq7VMwM+9rjBZoWbQf1PNP7LhrVztb4yjqMusQITM1a
ByODCcu9Z/NMBNf3yiev7kmjKmR1UauGUZ5lAumVHIsU+pR2bLpvu/V/++lTKSUV7DzTg6Gr+9/0
HPqiJbKmydtci1iLNp1H+jGJ2qaOwdMCs5bYdM9LkluVAbbKqlaP28r8pLsWMKxoinT5nVZayKPt
h6+O5F97T/KjxZzYzWpTEZu1Ydzpvvq2aR2xP/RxsXSEggM8TEJ2/tPBQLOSCDRqDyTMya51eATn
NI+pooeX64WrV5ahO2YTgremCWyrnX3DwBDdtdWayXkOcPHjDOl9tL4IMDCJyMrpy6P0cJssX0Ph
6BIFNqWs0unTOVULeeKKG9eXhqPuVOfjLi+lY7cBOM91Z3aMt0NIvPI9MDpYQZjUrvEKwEXO7jva
K36s0LDYfNh4li/xMUTSjlHIc+1tZgPJqlhgGtsumBW/qNyAuEG1ccUzrBU6aAt6gy5CaQCgPdk3
7En6X8zIct3/amLmHTS6LOCEysFaEJzxejoHN9rf7lYKy/QBn4hSl0D1wrdcE67UROtlRIECipTt
mFEv3eILo/b86BRorDkXcuBuNPL7Mx9//TXPAezc/u3C7pfS+facRSlNMfGKByp2+/eaFy1krSys
wpDTFXIODiDvc7s6lXOagyxmbvkh90NkgXGXkPCNADuRUwVQdlLKRKVrPCRqzlQkUeXaYe41FyGn
PkGy66Y1fbvrd6i5FtNy/jK4MpIkgqmtSHLoq2dDZ08Vq+3YGA6/DFElaO3bjzwbGX+0CbAd4Iwb
od725K/tOPASp8Pn4FPEgxeBcikA+IbQw7BKaj21ekUSljbP6dYstmSEyQgabzxr/jnfc23CvwQC
7hMMEuWgwBluor/ovXl4xAcSik47oyQwcbDJ0Na/mGlkTa9vBY1Cx0TG3ngKrBL/TkrXvpGGUI7t
+MzEUUtm2AaFBRMJPXeEIRxFBB89wOnH3SxCNP3Am/ePolrJr2hCXU/BIzpXzfSUojpOtMxXm5gP
+EwMdkgZh/rBb6Q4nCMVj/eMu94ExlrYxrDuIDPDBAPgyfhgLuADNHEe5tkqPXIyKQkaicrqAvh8
PbZAqomoxnTG+N6cTQUxgCWsIn4q3Wil+LZ5T9rvm3I5DBsqQgrfaG/f6rNosWH9E0VR4mYgJDp7
ma0bjxE/+yd4OfXXzqYMBi5lZD+LPEqHoRQeeE5wluRFm8ulZ0AMe07rfL5P2MZ9JQyCFzprPFwp
ydaiZY9L9Rj0I555D1tPuUUj9/Ca4dJkCgLoj6uA+O/QYaCT9ojNEikiUANlQRxxEVIOYoQQZ5iP
OvZzPCCIXu+OTBCMt7MEKWcrRfglWfnuwCCUAl6nzphHOW8TVrk9+rJ+BH2rgqh1cdD1OHV3/7BK
P17Uk7g9OaJFFc7wFhuzMOKsESh7qkgeNzDuuD7NbiLuQTRozqL5W/JkAO1MJ872reZME7bYMCBb
NHW+aVoHJxxoYgojlqC3uRXKgAkX5+dspYm/LCVP9QeNmAyOblOl8glxh/vjQgmihE0ox56WNoX2
0egiQsWL2nkrqr3+Y+HXt+ToO+1brnoJNJTOZcXYsipLIPIIS2CnR1EqthuwRYZUgp531LR9kazA
1K+hTGcEMVIRBWLpDdk1+v23Nq+TB1eAznR+3/3iLPuDWC8e+h0zf25O+lmCvyLlV/bBkauK9H95
LGc3ZRiQaELWgtVzkJ37F2tCY+4hRnYxO2KkRKIfQuysO48aTQVcvTGU4jheKtNfQ1OzArogcr4f
FBP64vZF/YD7mo8M79GRDM+e7iYgOnZyVjvcw2uhQW4pjhQS7RJ0vS4o+XDyeVCeisQlMb/jMo0K
xL8DZiK16HhX+T2A7aUq8zH4FCQQvJKucL7G97OEN+dWgDX+NnGBb356uijeulmhIiiAPl7F5q+O
SO4woRFWr4Bc4+imyjPO+Nm2Wh5awtrKWoT8/Nsvq+6Dee4qgqGExsMx7LJw01YSYumXe8AnoRkR
1EfmaMZavfeEkIFa8DzVzIfW2A1JS88AdP/zs15l955kYRbjXNstrqmABPVmechpENR8/mQguE9m
2EFg6V1zP/P9aGlq6d/fmpU1Nha7TygqLwz6TIqJIqh9HgUuXC9L1/5tz8hjRTJeWj/YGT0JbeSX
KevOSClst4331N/OUL4G2zJkiVfzJAkrxfNgRyW865IitcgIrqJ/VzjL5KAc/wSpg8UnsyPysOfJ
lk/hTbWO9dj+bNoawI2FFgyRf9EVh3R4ibJSMufa1Lc3LSigKlphnsC03fglmeF7INl+Fr8HzyGl
3IEW2PEnyL7ibP0Thl8xrkpO9y1miF4u87eQ58gCs34DTFeMsLGwZu51vdAYhTysFYfiueEEhJrE
zBgUOrQzu7r1Ho//QayGGEB+ljCwWyXnqYkDTQjiwfyzmc58/CfqEXgcEB9oQyb6azzMbBoeZiD0
hakjNbefxF4AyBScSj4Wq7vmZTetY83alG4VUa40L0IrcSZjNUpIMTp+47bun6prD7KJaMLX+Ukc
xHUWJJ5o2L8CywBru/cEnb4Ft0iaV2bS1lTMpWwyHAl8kjDqgDCNhZQgDfOm2knzvpn832ES2EWV
qVEwOFoakC1hwA8gvbMnWiDqPvIFyY3ZIVWRcp2pw8Lqbl6zrmU7dNyzsZAR4nmZj+WT2mewz6Os
EkcDzosCc68kPU+l9ZmDykPYt01fsX44DLhR+tTTNZWyA8xzuUpXLZ3Z4VsTt7zTdVT+Z5KNc6MT
ISozwqZjIEs6n7RTp6uaH5D+L4cmbXDaXBzM1oqs6Ek7yMtSQSHWxlLNdae7PVhw5odbbd0xl1HG
0g1auXIW8LcS41np26oh6yV1N/1V11NKygdIYhrqzbTa7cXLR3yDVcYU6pc8y4gRr2nehf7BtzZT
wPtxycFrQnS6VAKkb9wdtF9C8F7j65qZ26QCikt69H5wPhua8ZdwYmKft872u+xr5MFz5F8fF0GX
+qsKAr293W36NQZZNiPJQRFmBC2nP6i/Qeqaeu1OdiU+I8sSo/OIct3wmufRDDRBLF1mAIxwZshG
aLPGYyjlbT31DdwR1vmfjEvIheQPwOJSkiIqWW3UfLCSixl/e4MzCfqTu3+7dP9fKB2Yamw+9h0p
ZNfhXGf6h7gMY6ABudMFC9AMcPPsaA7F+mLRiLxun7+yBVedPXkAO4oMZ2pwZyWbuC+o/o8tUTWN
YyjTKXIVbhHDRAHcrL3AMbRYlidgfBNj/KDi2sA+pzKe+9G6zf2zfvRjfGRhsZz7aFkHo3cj54J3
YOG1V+Vm77VmzwlbvOvmQNKM12en4y2noRSqolh0EN08i7lcAA8AbHwU4lsjllr8rHpLYikShC26
GyhTDmmmVzZLnmUJrnlLp8EYKqS/cyFsxybxSgajiloAGoxrLxl3FX4tyHad8XBLGYoUoaoTZtjw
8/rI8EMgCwEqtGIGnk8KO+SzvXVPQQRUF932e/HrIOKVubhgIRZ4KNGxffHPCN1tVUe8PVJ/s1i4
LeXhg165MoiOLuP0zk//fQ/1gtV5IaYoFYKLCU8SkpNJYuNZTGguY6+SqWFkVk1gm7SPPZBHoznz
OZ9H84k1Fv5LeRGptPF/jURJgkFFQiBFZBAq9b92grMacjNb9P+YBE3MVqtw7OqahjcJhnUlnOQ0
IoE120CX/Kw/BXb6EQvc5RH2/4VELRjj2QMSbLurGFpFQ/+Bp2Go/31yDJCqGlNNgXrGGUzMZ4UU
IOanqCtu12liBcsYEiEUVCPg2mAbRbChQy6EivNkdcq/r//TUUvxmAWma36WQo+IQc3DWDIJEkDP
RMFI1Ua4FOoJe2T7IjceI5iuPwdy6qxNC2f0J+WcJmP+bUwhhjXv3qMh93aq4Sol5ekXDluWgPpt
SNqbzYes8rIybVc/DW9my03n/r+VCOmD1ALVrNdwbQpPKFX+Rd4ccmNkm1aEkAAyWTgU7eK40DRg
DszmLIBy3TvmSoc6JoUeRqkX2xWwapxlEvuemFi01CAAePJ9rweLbhm6xCgGDF93uKy1Bt3+a5fo
EkPqRqm8Y8yv+kGnHXO7dBFuqjcIF6Bun/cIJsyaQx1wPgFniOLQv5tD8XgFujZwhusq24+odL43
lHJp//4q9ByKB/EElyTqxnoGpoi8U0fkuyiQkdwrrhqSdLCJYFQO/MhCg/ZPpWUKtQRX52RKxCE2
Pg9aohTa1YNYW/Z56FOXymibr1Yh6Jmjjc9KHIjWidVDCQmvb+Zp6HCzX1Xn4EnjFX3emAD8XE5y
jcsUDfVIQFVBOLViaJY/noC4vX4HBxNuy0NM3v4YpyIfSrrYk5zVir4TgnRJnPiCvt8jP8NNPHDw
aKks9N0QxWihQXTyoq1FwrIXnttj7jvu4d4Ooj6tIBt74daVxU4ZUGkrhn56zaWv1YjHzpto2wtd
D/OA3ZS8sB9oEW11IrnM5EvMBuyXoe1fdlMy8Rr6TcKISNgzSnHJo2zudV7YggNnB9Iad2o03mHA
XPDg3IfTqYaw4r5Li+461jup4+VCKQBctrzrjOQNSV0YvmnQzqAhavOCDqaVemmveVTVQZpcMmHy
AdhSq4bZEnD8GsCL/HMMTkdQv1vJWIiZgu4gERVLMX/yXtoKHWrhBSczRmmRvRJCl6GcTFQuVeqb
Bt4NwPpJKkHkT4mr+6Fqd9xkhzMMZqRixPs0L/mdemw4a4GtiO/gF0CwnctR7fNtEwM2Zwi83gjg
VI4IJE/FtcrNLP6QkFgIgqsx2xhK9DNcBu2fUx7foobgTYdRBGQ48dBQztgQhhCOMqs70hc5Hqpk
z0H6y8UC3PP50GM2878n6jUcsI0QEVHHhCZsIfqB4md2JNrHW5U2Cm3SP4Rd9oDL01xBSEWBVkqi
46ID+uVKmoCuV2uvEQsRpDzFPwxfgOEJJeNl7DdFMxeaRv3oza+R73mEAz7zL4TFrg3VJ4049npi
FUKMYQSXdMVavEEXdJe4/T/T6+vBs1c7Sa8tF2IZnFD2PmYRRH9uUQWGYgZU9r6gUecHqgLxu4nL
HzfB0CjicmCK3SvVaYaq7CIhx8oW9QN6/htXdj8fLwB7t7TlpqbbyavFQ35Q/BymVMCZhpovXv/S
hJYmndPzwTQfjlJzNBc/3rUHKs3tlmLGNUuSO29uDlPyD99fRV8aCl7eZ8tMN2PJtfsy21hLXiBk
AInm4gncSqZC8ByLQeTvuQrdygiIPl386qiGXjsN8ouCBkuaKwbrj264V9Q/MRmpKK7LzSA8ThxJ
r/xe3yylBdDUrss84T0SndHfI4IWVrSf5wKdNnzA4j/tUutjlaVJouRRoekJinnJIkOqcqS/Zpgu
IH6m51alhy1HB83gVqwaVIEsYdZBINBITQqnoG9WYbPigE7O9N541xalwsHOxLYrsUuYRoTF95Pg
285a6osDpN9iG7Btvd3+1VVBloDiEV1iqOb/+ZRcRNREtqgiQ0v3hqI+ac92hy2yTxVddw/ELYPQ
zMR1/ejTC0jjELetQenMT2G5HevCumX4+Txp/PT254zjjeQV/4rQ8Kn8RiWKlpuT5mfhWNHW3rp3
cZH1AFsFUg2YWvu/HkYH720cqbdXED1wYZefLvrhyjVxevEiPH/7Eewa1CJhjXIaoSBtlXNuJYMG
MQo7UO/xHtr8MLb0cWD2ENAJM4DwRtIVNqtWudmVMMp+XNKPzb7dCdw3iDM5mleT3U5FiToZ9b1N
6HvRWzSTX6ajsQIIgxIu70JL4LqYA/IjIkGeZ5guLqHgH+SFMSiBggIOhjHDabBxdoug00ZArXp/
LePCy4X9jm45HY3331NG8nNnCUJceO9NljrDmvQDEYyM8QF41LpJcBk+nG7POsePzRYiNIdQ749t
ykidaWDNiU1GwLjPFD1dYpB/Z5ktCwy2UgxiB6jY705q/tNQTjMOJm1Tht8CtDT75TJArIcd2DAs
vt/P3RX9JZ11WchV7ib6dHO1DJfPFn2LCicq4ZqkE4XpkKyQAc+Ldwd8g4IXRmKtPUmQkqsQ03k1
Dw0hVGDGudITrXIGtvbcklCST2E0+asbWyWSHg3C+ZoATpCW+6OMZrpSSv1ze0hSYvxwpUIn9Gbu
2jKoPeh8xqJ0K+pwvHfa1ydEnXe9ZG6ePkXevxCwbiRGnXEhQs5Me85NaWlRXBNbOG570sfSoOKU
8tuP9V2kq2m+5u55VHM86nBxiwF0ilzL9A+vI3N7tWIi+0p7bCUYoXvutnkPtra1uNammRnr1Qv+
SUPVFj/SVfmpE2vj4j9ESOxVE3+kbEA4PYpLAY54MvRLeswFn586OlWhVJn4HRE7A7V9OBElGc59
FOMD0Y0wPmaJzR5T19WtfjWQB82YgtVp07FaEWYrlwldDr3Z6buy0ZMgrRlb0FlzEcqofmSxno9I
klfSCyg/h7WDiSMTZVhLdFkdJeqknPipKWAQD24kaIuy1wP+Pf7Ikj2o9rjbqxtGvTVfjNBjCcmR
Ri7ggqV5vHckvA4hbgctbtBik1U6QhOggHnpn4L7dNChbTyOId0mh7mrf18sQUlQpPFqWr6cSaAC
QIzJuSUtsziBFHjiIS5gHWYcOWqEwD1V5znCnadRHiV3L2OtfzbE1kT67nkdxgKe55yaBWiO+ptf
LnpsJTlesTZDTLtgwpVUPp8fERWMn8TUwHfYioclUS9MVYORKjCSLDlDg+T1jlzE4prT0uLVcFeE
WPTqFvow5y6BaLi+wvDQtm7HutFy8suBi0/nCCvs8Zd8acFED2elcOwAKB1tBl4Nk74egUDjdEYr
8MLT9MlZgwY78l75+qlVHTl/HpKHwkaxrOeXk3iSdz+x9I2vTVuGb39EdqrMyD9JgO/YZ2TEgC3O
vCj1uMMzoTKetot0ldTku6Z4LmjBzxvY3MBmQZZaX/zq/P0OsBgPeU8vXwtyoDT1HO664FDHhG1r
5YBA40fEwfU3Sg88TbkXJCIvxSGAPrsjH2IoT/0/ESy5AJNIiUohFDRZeRp5qsuVzijezVf5iTua
97kySgX30OIlDSEqMaV74TEoANLAqS6tAp2Rftoj+p4CNV2vpYjgrV6Iz8M1vWhJ2ywC7xwSvarA
xPwIghXu1lnlbNr9OqUupE06iySF7tQRHbUi/H72UhfEEvZWiaBzFpsP9UlO8jlRQRjNQaY6Twdb
nYO3+yCTaKK9hzOhLQRwydbKZa3+AXuPMatKx5XP5JcV7CnYD/xAnid1wYD1t6LYQJ7N0dgdNMUy
479G4Fuomcd8c047zRkrHnCOKZa51oaGsvjM/EPYsYH2th05Uy0p4wZ/WpVp7h5kH97yVp+FdGI3
sCJ0H5RcFzoXxGonko57xFARlIpj3IWJUmK/nQVpegCLTcfRdE331hetQpMKjpH0B/nnh6eCaPvi
F9Vd0SFTruT+HKAYTfR9GYmxVlYcHnotSRhce7PiI3jlWgi1zl6OMsGE8i+jqqGEUnif+soxvaq+
JeJXIcIAngFBvKV/a5QQHcaMz7utUcbAPn9+eKZbFlZUxYqqCwAkTIcHZkzJsDJn1bTCQ3xMUEQ2
5LSYEdL4ZchTdUx3n7gHLvPP+K6RawJN9D03zPZNgkcTf1qG//0D9iAhDCpnCtTc7J0uOHyPRJVh
03XkPS4XBBzq1+HaauyoP1pBLSsg1Kuz+SmPkkuZQ/TFkxYj8HwuiaQui04abWwIjKmW8djYF9qO
6ANVGNpE/LazW4K0j7EifNcpaJVO1KVF012FJqA1fYIMH7a4Dmx5ve+2xPIX1OGFP+4VbTUhUpEj
4+3m8du7QnHpKKyXCCbT4+q+4R3rkVyYkEJvaKsv+cIBZ+LJqdeA46cQ94nzQr1nFboYCqydVbp3
4eeLxtRPrKbCkK7kskwxOGYhpSPfWhx/Dx7lSM6pvoI9IKspfgddDSa1Cj/ALGpZ2lcTsOnosoaV
ZhZsT7YzWZZAvKgtGWEmTNfBBNIM0udnxX9snQC8CMpjYT3Z558CimYcZR+wG3bLvOHRZPnaNmTI
7D7n/3pZk6kmkgFPP8O/1Tka4mzixRHb7w8msYxPcCDhUTDuhjX8XEisUmIp8lgIasFAMlUWmMOv
NqtpkaXbZa/0Zim37xzgHsuC8JDz6WGUoZX3Vpj1Ua8v+mS/flQaVDcvYJom8B+pyht+wz6fo0uv
KGHf3MWJk0hv4MKio6Vf2d3y3y+dBhOhVuk07xBjfmCK0eog2KubFyMrtmpE78w3e9HiCm31HIFI
7RVzcOrsDl2tX7SuU9EwFCmFNX8o/jIPcoCLE/bhwwQ4kLHSEhe8vVs8YoM/L6Oax9u4ujM8wdYz
/qku80RGVwaboXXBUpdwBuSCAox+Su7BiS8dw/hZJilyq1lX3j54au+OH+SxOexBmzmshoAPKBez
+V8fRbCdsSrfKkEcmII78Ti6VpMfZy2SmNz2Uv/69+ACdqlSuTBz1PlRYvv1VK41WmA90SSmS07m
pv7meyQsOZG4LlS6QZXYau2afmZGEVGxBYnYYUZJqOxjjef8KZyldSdHlDdtVFIOrQOLirBETF4Y
onye3XH8XMKKnLXoA43APTFpknSH43puJFHFUhnYtARE1BbXt+VerAg2m7EGFsIeJiQGNNHOtpI1
33UGu05QPQ2DrVE1uv7YLa00B7IBxkBsvS8pMcqSZ1IMylW17HvX8yGaxjp8pd2/KAHnItEKCmKh
Vjuhuy3iV+eb1d8IVDB5N9L7V7f5/JuMhapTbg5sL0AjM/GOjrq1GiImnZIZpupqlKlja/E463BO
eNltrtuxKkfkZJX2s6CBceLzmQ4sKqS1TExrugrR6AyJOA+PDLKOrWlrCfqguvCW0K68jpeBfURh
MP10ylTJWMwO1DNwXG4qpXjR5m+HTV3krbUAD6gFdY7ZVSuR+S/kleUS0p2ik+/Xdf2gnkwWQzlW
d7lyHAOtY9TexwTIToqV/YpzBtlSf+TJs2+/9qBSuSdl3n98iDmZkNozwtayTgNEgtpZs3bMkzwk
oHg0GTMSALE6hbRFoFj3y+xpKPOA9bqgRyAAqScEksDqvT2LW7EXTUQ1dQ1q8a1w2QMqM3y5de5Z
eVuzF/KnlhQ5ZxvWDQ86ltQNZEW+e83VQktpwrw26uFsazDl05bl5ZRaQEP/QgkeBkWFKf2ffCrX
t+TGcWsgY52zqjX8yO3SKfSwhg32730qKpYoxdrK4Mm6XXEXLFk1U0USFUMrlq9dk9rwsFIQ13yA
v5aaugC5qRJV3KtnUsnkI8u0fKajCJqeKuXPYKv8dXzy96ovkhDHR2o6QmCK3Be+gFiOgDAVlfxq
sq4KaZiniZsv74pyKFp6y55H+/J2vsRuBhdW7FY/d7bOsVkyQQDhK879tqSAj7yCwR7E/GgtqPDC
y7c76I+bs9azKj+FDhrC1x1Z52cFaNvyODiQSY9tWyT6wqQBsQDYre7dHOHxl1SofzySqcZ2TcCA
CwaeLKeu0Bi2GnHCvBWUCHeXFBcaeU8Zs3RMtp5S5+vojzP1hp9iQQ7dtOE1jqE8FtmwUxUkvOHn
neaqZ+lpz3tSeBPxJkfaWxn10pfodXasHzYRBpUCm+Fxs6OXuPyD0btxuDyRlxC7092uBhBgljpo
nX+OaWK+BDuIy0GQRs8FornBYfkgJx6irIMvM8f17M22n7vpu3EmpaEV6QJybLTIwFjhjuAb08ty
5nl2q2/QmYtuvLNDsfnMl6ibAbDdWTxpQ42FpzlmDJ8ujIAYhJxrQ+3H06sJ3BKmUkZJl1QhC++d
M5iRO3ApuRVYf6fcEJj9W39bj96g6Qyp08vmHnS6kiePXeeA40b1zYKkymOykOGD7/qld8PFdROE
sxw+pY6iqdWCza374pORD8N/XG2bxNmhkHYQWipT4hKOxG35T+gPR42XJoAuKRvmnFWFZD98Ct1H
C6RpBG2TC8BiNtw0ox25ikNLl7DW7J5wL+eye+fI+dnBmSkHb+9tmWuQU8HGeJ0XJ+kwZTiGh/+w
nOJZC8hZfn6lODMncjoMK/uN1Hm9ZycZmGn/Ji3w9L/hYMyCFmyV9DPEN0Qvc2DF23SvUlV0wdWu
iwbBO+Y4o7/GOdGk1O5X50LOYL3epCn02AkP/TdPApN3Yr/XqxBY/zYqlW3xBPaRwpzT2LcpUu3O
6JhI/e9fn9M4ch447ItAg1Fnsw6YN2ZFx+RyjNMajdCtr4Uly2kOkuryfvUS0mN1Bw0kculXjGpr
vQ6/ys6j7HnBWBtVZBHqgkqvHfDdosZG06x4yGeb6zFWB8/2hNbe8W5eW8V1DOreXD/jEESv04uP
9sozzp7Z77WY3TSa/hymxmCAH/7jXdq3RmrPCXh0KgSQSHpA+TXGrMBB5H7YrUSpYVtDWIHjZeK6
sok3D34tija4SCn2EaYC7F/3l9hKuSllSaXgfKULMtJ76Co3jIuiaZ4A3QaaTZ5eCeUuwKFCnnup
/WQ8ScQzzIb+2jgsVD60Wood7idscrT+zfiXQgUYwJwITl/Ldoo01b1o+IxVLlT9Kx+QucKikjhz
gVIiYrMQKulTXC+skhEg7H16L0qiWT8mh5ybgTACquYdOfCZMPViHwqLwy+ibsdVlp9sFMc1nHPR
JzodHO6kUfkQgJ46Koxl5f5JSb/j/1DOFr5GaJckTGy4M4zcNJY6d11s8Y1w9i+v5C3xIovCn/SE
Lu7phZF+SRV0F7ob6XdrERw0cmTnKShqjYSc5mNMlQD5aVj2jaWtgmie3X76QXuAmevHgAla5xtE
rUeZr3ihgwUukcc4FlpustOSh6z/tUr6emyZT7gEm2/YHwJeqQWU12X5aNv5O81Vx0TvtIpmOqbt
fN+jcBeaqkMuyLMbMy4AM9nz4vNySa2txKrb/zmYTLQG5IaS78kbaGgREON55V038FkJCcCgmW7f
eM/W9YrMASH9clauSJ6vH5qvdmIDgo2QawgEdMPwhB3gnNBDyHJ3JTcTKRoDKAE1R6qWlUhNbR6E
9FsU+JE4NUd7+SB86ep96AoRmQc2i7phhcGGDrYs4G/5eRKCFySgISmQ6igcHzJueCfcMfxsnZZl
a4uvIYv/1bRRYp7IwPCojvPMMLfExe98dd/txdJtj9KArAs7Pasizgk9gLYvWM1OYwavDk02XmaZ
63AptkvNCE9pCjhXTZWZ4eoXopttOi5/OCQwfyfU+K3n4IjL6Vl04nrcrpXsVaoB5+Rc/EWTllkB
3NELQ2dSYyYAh4LHhz2rVhaGJrPB9fgMD3kmAxbMHUYjNcnLh0PzHninK97acqvOSMhsUa4P0YHX
ZclakL/qQeGTGe+IxYUf0vP50uR0Zlu8ydBIQsBT0Udx3+qzH69mmbOD9qqGuaYKZPl0BQG+o7DF
csjqNHt8Zhc5/UVWzTzTD6jO+FwUFsZBX6uYGTnaBOq7rC0/qPRsOs2qMzmKgVRRYmdU/VdXFm63
sGHAQk+Yt+S5QuK8FWxzD3oeUiK46nKbYLkI+LhExt1Ix962AFZHa/2cleStyc2UWDtu+RrOhq9i
WkeH2iFkLTdo1Xu2QWVhE3e1GXR8rov8Uu6sqcbg3VEwzIK8VCgrfB5p4kVdfTjmV6hX3o7E5M0j
Ocni9OLSWwxn6bgk2wyl2zaEZHHkQXi1o4li1nlp5mUmiJ0fBx+hc0KMgc30xlcnNmk78SmGt3jv
KdtfZK6YGUaSpFe7EkXVJjZ68p3+qtxcY6Gfzh/Tk206Fq3sN4J7p6kv6hmk7UQeAYbSWVkappP/
FfS5fXFN0DlaIpvniAt49BMWNHMzJs0lFnj4FRctA1xdOjs6pAdTaIKRFfw0OMmoOCTyGqAB+spY
ru8au8iaiftKqSYDhcTHMGNmiLtTwvCXt44SeEmohXnfQOw9p5ZNWhvtOBhJ+9rX2miP2cRUs4G3
xzUrU5rhwKkyqJ7S2JUCjabskPuJ3gYGDDu0zMPSCEEkKISd5dZj+aYtAF3/er9XhA7iRJGHYGtr
gqui0np5RgSRsK1lASlfY5YRRVlp5d//Wa6Er4Q0XM1Y7m3PeXWwGjnHyP02KxjxHC3xQkfgSSFq
cscZUlltaQkoVAUBNYIDnQ7/aD5EDl9S3lTFKB5TV24110lSjAt/gMFc09Kfk9j5uspHRfUz4XeG
RXUbisI7wxGGk8aoajTjMSBt9YU+T0GlNK9OOjZD/Vi8SkGQ+f3tpQEmXePojLvGPITSaC0ezWPT
Fd1ly0jDLhYV2J+OjVPBgXKtAH3R6O3EEm23KmjN2nFpR90HWCeC6mYme318tnI44umCIG+s4TcB
wv7WDfcCUlUeSMW1Wv4UmkK7ktQ2dlsnaFo9pkSvtVTnoric7314YhlXe1as1j/6BegP/Tv1Dg2N
W4Pt8+glkhVgGC4YEmt2HkgPLKrjTsmuVXPAEEShPNzHJVJgB0J0o29NYywnQLQjWsvHXvRjV5uH
ORdftKgudo+alcIc/Q8ICo37aRGaL1z5IIUOrYm+289kXw0sXvFljF7D6S+MLWiUapk83oqOE1ui
FM5NtQ6e99st3JMICmif80iZ6Uugj11k/EMz+zDf2S7D7lZVHW9bEfPyeK2EwUUz0NNAKhPqpeEP
jW24F7roMvV4vD2NedBHTmYBF6vY/rnxiqoovubMlGLyx/KCc7zp2si7Q24x52m0lgg5h4iNm47s
yo1MW4fFL9gk6bnCI6Np+ciFSdEgFoCA9JKnwKETulT/n43LiqcaMpsArEtx9YpJne+Kdp5NAGw6
EeB0PwVU74tYJnYYTCl50fXop/gQ9s/BZtB2OiLzzFKkSeMhDyXpStSIWH8k7NH91FIyiZftEQg2
xSr/uiDBBac/4l7gRVFj7mOp36fpualXu49CeyUWiPuN8VpDoFh1okmJsrO1EZTN06Ayyz1CHYvu
SSO4BUWbTZxKU+dEeThTa1TN8Ym8cCL1QUS0cakSLUBr5vJIHSBh1aKh/CDz99XXsFI1sZEthYve
2XBC67qy3SQ1pyJ5b536Q2DBe2oGDe7EbROQeGqfyMTiS2PuD0zf4o0MnqUm6WkBNQRWwesGtKWB
CLAoRwYVTE3awhdcHcV1JmXX2hMsLW6Et7FBaRk0KHyHWa7JkDa2tm2j5p3uwEXln0CFRt+UAjUf
WW/iu5NrU/auhvtXvJLNzuPpj9A/LqePM1KjPB3gSamlz0Fr5iGT+Ftmdps2JT2rec66RQJfq6tI
oFFN4yw+Pm/EtlV5Dg0b20rpjuKp/CxC6gH99YtywzryFZfUdUZ4PMDalRurQkfCS2kPHL6F1uke
G8wK/q0zp6bT1/BlHSNtB0LtpmJrzFC0h09MDFWnpNXHIMRHfzOg9vRQPkLyhECVGYfwTJu8NeFh
G40+jnzZow9fDnG8LA/3ww8Ip0QujAkf37JftXj3LoGEcHgEVXyF+6TBt7OWfhNgdrqvgSODpD+7
9Al4TNsNVLJrRtJWNHzLRo+LAomYyES8F0VYneTkEaxBo2GHq1ennghO3fAYzkvgI2SzM4vCmdV4
9cUhZ8eDFMNY4YMmyM8ipM+MRDDv9r6EGnB8+wzLCOghTn+tDiWm6i9HyYOL2uvT7JvJERoFJ3pV
vkjxqyxhIico9uf9URcTKjdOLDOeLzZl5znlbta33lYH3sBvFD+Ma32SzExP6PI1HzSbNZJM5WLg
evGgeF02CIBXDape5pmpPzliJykibFkVoXv5dKdXmiNfLtQDxLBCOqbUFEokpPcajkuU9rYQNZea
tsQZzki1hQhb46axtJXOZJO6G3npBqPSpm89z14IwJdowAjpPLF/QJFW3bMuFS+8+jIsLJ1iSeYh
3Q5OXICBg6uhupnrp8OSi06T2sY5IRqSmqHu+Kmw4nGK6zhsU+Xb9XFgjRzMt6+SpjPXRuy4IBX3
+D3JDPMeMC5DtUmXwZmwms0mPa5RtD8MFXkz6OZEpVjHNa4uiTe7yc2Q3hYujPGp9Gsi/efeK0Zd
YzdOryfmJyBytE9065bYpydx1ztVM4Nm38oZ4lZ8XoKGfDXEQRg+wAxosRB1L6Vwd7UQbdMIOb2Q
2dSeq81Iw2DBS8egophikDz5QiUkoVVSIjafhKCHBMnZIWSIhZjjvS70fVxC7XqI/VlXClU2mmGL
sLHCew1oxMekmKCQWszjVon5IjRUwLnWDh66RctiUqhdk4zdAuFrJk4BK0fj0xZBNp+4llfFGASv
edM+yISLs0mcWuwSsJzVVaAlhixkbY+VM/VoWJjLoGAQY0JqcNu5ABjzF6GEdWB0oxecVJpXL4TI
kv/THfEp1MHV7WrtUetya1BvScx9i2vWcui/lTeIH8DJfcgU0Q1nSJyhnI7RZpWP+gOBEScF0eZI
KDr7JEJBPKfpR8Bck6eIzFao1VbzE9o+g3t/K+uIUdEfHLuYFLPDkEGDoNcw01w9hHqNwgkASVYw
+4gYAMHUqgLcmdsmvQgGoBltVtCVMsBmyn+u6IJJgfnKZoCD6NC8qehFQVP7b57r5Uz/QzIL13gP
SKcaqbHSHsxrx/xopHAp+ihxOT/9KhckxAFeV1Ju2qiiK1BTg/cD7CyZTp5Mo5GnuHsEkj/vZIKU
LYtiqYyVeYd8X2dyXt8hUGb+CkLsZoZTV1g4cIyOw4J36NZUer07XnXoVxaortoy6/Ozfa906z0O
HOJNYoGbawCm9qqXijtHwQvcCzY4PhGUmAtY0UQMXlNS8KBQ+TrNb2NWE2Gn7Tv1gCW2H3BIxffJ
vl4zytpMu1z/5hwz44zOK88Xm2G8Lu7QRc4SFeo9Ff4BtWmntgTeNzL1ZtVHTerhcSUqRQ0JLLPA
VV+7Lld9NHPxc8ZawTigEnMJWHk7JY9l5DWcP2M9bLcwtWvdJoy1LCVLAV+fsfe9e6c0Ms8fo1nL
wa3SYir5PmnW1SceuumtVLIbB3/YZDT/BUgSK3+uncdm5JCbk2wNdWO/XRAeViQqgK0B7aQp+xZE
quYD5vOplbyVEg7COTzxGIXwTIvqLHSOfLjxLpt1jPMjS6nywk7MvnXZIG16su875iIhZay4Qy+5
YIx1ovCWh9/iiI5ORkzKoWczHBLavvPFsbpnErZebNHTX8VwEyKVhIoR/QSkliKARE3qb9MQNCLu
dubdDDHYqwNvM6Lpv7+PTAsflLb3xo5b1g3E/SgxRuqn0kCnX9ZEy4RYrVAv4ZPwU86/EGOBTSaL
CGC3SblC9JJA+9wUaBxBUsvZogKDdK9oY6MbB5uaeRwtrJDMgc1buYfJwbxC0QFfAefGMkVHRU39
dDTjUecYUSgNmkIaf2o4lEaFqfl9mcuUrkVAzuZXJYOQMK/5in5Nv8Bqoi+9yBvb2ggVTtmXH4nv
+qCRdXwShqt0EECyqCNLmFCU+kmMlXfFxw4NxrWDGfJPk9t+HH0FAGFpB908+G+Xzx4tp1Rq9IAH
IfppnyuEaIdi4O266Fymwk9GiYhbrtzXodCbvwr3yCEimZp1cJ8NJ8LaHbjbpN7MKl5SH+59YdXh
1AF10OTRGaIkifNtttAPp7hC//q7xf1/DUkoqxkgOA1uF7CJeaL8DSCaJvzrHikent5kf1+TlNvE
VcGE+a0XAhuMlAn2WThHpeicnHQV3PyBAuX4tlKvx021wRt40dEt60yQN9AZ4E7fImcJsB8o6lvJ
cONCJu2FcCj7ElhVbZDLozMemjSXPJnvymv8xN/6KHHDMiSbWo7G8vJDOQ111FDmwdVAkj+J6uC6
mAJD1QGbvx05SocCG0TJb2knSBExmVtSk8Fj4hxQp2s2Lf1nMBN10wlipeKrGI/GPhCp/rHeLp9J
DjmaMHRZR4AzMq7KMApi8pJVfbn3COA1Hnzc15F67bwgShp4QtkAG8MV8I9nhttWBdHlfXHj8PWe
j/j5iZohPIVaDh37o4bWJVshQ6+EZQWEjk9R8SljtJv4nWGjLukPaA/3AjZcpcPRnE2qmvTDu3I6
KKfloRtRmuORg5Di4KBAQ1TpFrSytwgG2qkZ07/HSUp5rkxtaa3cb8suS3sf2eAXvvXIXLYNxuhS
X1aBLniEdwk70slX0KtfoKYRhZZ2GAzLJFlgKdJvYIP0a59gECYxHQndi4CLUAgWF2Vl4IcTfTYV
08ToJSy+cC5Z25gXuexcdVvFFwOZLsRLV/PWVHOjiNvkga6RbsaHjlNA4F6DT4TcGQrCzl/IJsvg
lgPbpGDlvmjmM7YKQ4EQDn4h6GKxeAaju2SkmFw4w5KY/ZE1SxXlmwlXaDNwkXEztp2dp9aFVsV/
cdJEEFRJb0WNf5JT6gtUVxlJQ8VxICMI+1cGj8CkV/9pdYmhZTVhqVkpTltwrnomxaX8kCc6Z0Wv
bLxWcVFvS5IF0bmSRz4I0SLrynkRLXq+KsPA+mCwBE+POP2mUzqvNYhZNNJRyJP6SQTiZrt2s4yy
lo+z0xN7g9LGGwlffBt5tQUSR+dLfjPRFAmyHgs/fr3g4u1z4iUVlwyR3k7hLrncAJ2Y4MbRwz0D
SH97hsvuPoaq3tOcOZ2dJllAnuB8L9Al18ynT+DkSengkQ1sGT/q97PP4+c4D+xb60tNe+S2L1SR
mK9XzBlfC5sRO3+1v9DD2nlH4o5a++ySL81a4qPXRRP/Eo1GcP8SyhHIzWgNDAY8wS8DN/K3XNOj
049U6PfQb3NDyIysmFt6AFoq9K6xhBVnKHMrF8J7BOKN5yUYBGPCa5OVKcCnjwwG2HGjHIY49zLH
P3xxlBmdBsnplA+5bR2CCImZMNhyTG5Df4Y3QXCAfv28IzgIHbGB3zCsrull29OySvIYkIfcYRa6
zkpQufaaq08xhDp7ESRBgCBcvqgaUECDxjAQM31BPx16rGO3pv4YbheNkTRoYzs2BaIglf5IrNLT
fks/ulHtgf/EaiKiFAiv/nAGZ5Tiu+TA+erex1q3IMnDAhkWyf4Lc0lGUZSBhSn7yJlTARfElVep
oEsjJM3Eq/4+tvAR+80H/WpJVFp7dZkDLE2isb+rAWSep9uHVPPpCDNpVDv3Stp0F8yrWiX1IUOR
lws74Qps6/TfEGUBYP+0TLn3/SMxC2Ina3SKuauJZNqa/GCfRAtKap/vO9hv3FmLFCJ1mycXeElJ
MuySimtyKc/BlkZLIPuepusFk3qZhJ+No3sFCDVkAlk6KwM86XitPgM8NUyPomcnU86jP+uS2z2g
eN9bKOSoOEWtnP6ze5njyTut2HE6duQ2FTUq8F6nDKGvCmzMMfuEJczYOkFNwn3IKXYa53ntSwwb
57GPDFwcBB5fpYtHW1qmpOGy0sspm7IHZ2jpxRu8Q2HNZS9GwZqj1m/96vuou+SEICbK7+gjtJF4
nUPmhVYiLQybiFnROymdeYqd8tGmx0jpGs9uC432m/uGqFub+20RDF3Bv4GAiYeTXywPJXVKaxGM
+PyJYhlWqlsR/QSwFaKFEser+4M3G3s14T8cyQpY/oTDWAdJv3OPjuPZw7NOytne+pLA+5agu2lb
oq+2vxLXZW1O2tWwjo1StoubTLJ2Xi6E2AvUQzhGQ+vLPQsWlAg8oChWtF0TCsN6sMTmcZAHka9R
6+Ckm9F1IxycwIeUCH74P8FLTb0+fXYwribj+awgFz+Fwix07lJryyYhhenovUvNfacR7pMh5EBW
nUACpYth2vMWr1N3uJj5Lg5aKiSnnh4j9IIBEePCWaIy/0BPS1klaBLKoPDyoNzBZKU2tj1jZoM4
iZ8xDSt8fl4GoRAuBgwLKWFNVqaZqg4ay0saZKXeP90uy0dVPVWkPb7jCyQoopyhxewqu9ooMyVV
+xNosME/DHATD1ezGsj6qGYlSV0/nmEfGHv+uw3thQQPovLcUYp5JeX4yUdecDo2dkkPLt+zlLp1
spckLhqQJTfUqpeaZSuBPdtKHbACUB1iAWUgVzH7LyDyfe2zgFmA4PdWM8SFk4RqzYL+Bh6Nwucw
djPpT/zDVm3EoMkB0klsW3M6Bx6D39hGXVIZH37qm0/GVHv9Ifn600LjMD3jOPnuwHu8Ug0Ykc5q
1wVVieJv9pnrmlIx5anP5d3uVHAa741+I4XBHnUSPIp+P9cMP0d1Q/G41SJI9NVNlj1e21kftosX
R/tu6wM0vnWtvwrUWnsbeCkCF/gFlfi5PWYcRrFaq2b2KLdNB5Ueoy8rgv7w2WAhSyPgxsB1pbQC
6TKVparizxGV04jEwxwPkv8NyvgEQT3lcntTXy12DOmD08/hdKLJes+9PCpWLMaQ4hY4NCJ8U44Q
eTEXjgqEJKvjeYKA6xmO1zTm5LBn5Q0QVwQED7+FOgJLmR8770lGHS7yzciCQxiTC+umVaWHt5kS
cByhzCQ3sralQxrgb0TjylZi+CeLjdueq2cf0b9VRS8BNOm2lLQAyMcEk8nkYTtI4PR7cllcYgUG
ryC/8cqcXDYPCXhFWvjH3XWYhMtYfp2Alrm3/32xorEN/ECT6l0MIs2ax702vPZEHK1U8qWsti7M
RNXmd5UFFhs0Jl8NzchZZ0lH7YYUxlphqhQZ/y5ORYempDHAJM3t/JZcZOk9KDKX+p0CcCYgwI6d
4pBgFsm6hvGZx1KhZN6HJxEQC3WhoSiiTOkTRGZVI2GBKYm/TMe6MbNk1gA9zed+fgdNH3dSYheZ
gT9v7uAB55yqHCIyfceCFv6fHN0KxmZNkajsiK5QRq1PiwCojyVuH+N4N/+PWUfj+KQsF8PnJ7UP
qCl3IbQNO0Y/l7zj/4EfybFyM0hjIT78XXWxIU5L+cxQ2Yv7zR3L9xbNoN0R7i8NvKc5V9XNv4Ki
khrBq+ILnOSvD7Y3roVqWNETvDklEl1J3Mtrym0eXrGX9yIZVo1lXEwMPyCTLKNtx3nnBMcV6sJ5
6EP0OS+zVJ4bXvkJO0aj/hYcRZRB3JuCls6cpNfYfhy5kL0oQkbj39cZ7V45u1zDIJN3inQmtUZ2
5+G/RnwnrhendyPXeOWQ3PYVrbCqebWvCKYfBPAfOMidWwrR5h6ZGy7P2MvfK9kiVDLi1z08xUi2
LNbb6lG8OsAakba+Dgh5xdc93NvrrN6XebDIwHeCx0ecXS5Xzp0hX7bRLPy3ytwXg0Rd2GN2im+Z
P7NU86c6RkM/cAoToawMGTAWSc/wqQp47G6FMjNxZ3vFWh+G4j9LlHpjlOt17gyUfOd3EJ/1IL46
3tSZlPu6nvF3bOBoGzoyBxFIreCk3NubzgvNVWKqnORYWt1T/jnKpjDGe5HftFKqwvPuwMI+cWGO
9AM4iVz/EBQMMs2uqIAG2cKRjUMB7P4evOVwm/JzkuuyB+ApO5Xo+f5Qn2968UKvox4PxGD/D2N4
WkPfZYyWCK4gmiElmQ/VUo6gxBdB8gTUR72IoBH0a9tyCm16bKrtmPz3pshz5Iji507Zo7RtqNIP
n2Xv++VZT7a8c9cohACk2sSBvK7k0vPBqkv0+G7N0fmFoRSQhzb7Bi49M0EeIonuvMWcfNdKtsdI
1PEd8/kIEOP6sO1FcVBKh0YlW6hHkhopoTQjXaSG5iIAcgQHxNTv3ySL7jvr8c3naC5s6LcuV2kc
tMPaY8mWIO6c+L/0Wn4mhOxyDxGoX6mmIL0JVTluB40Y//PagwuwoXJL79xITkhSB75S7D4tByI3
UcUObEvAqDEtVhuCggqkpcgbZB2gE36NU3ctFy7QSJgXbWjkZ4pAdklc1EAo55w+16bYfdv274Tz
D4J3yb9WCVPSonJT34PiWG5bDfk42k7hUfVzd+HiHcVPCdk/oUqj8VHfTreMVTEjjdVvL/Co4JyM
0D3TctkUCrftiRi+e2RX8V2TzyrY0s0CZVfEoOrJaF3B21EgqSSg0uTKxbx4/CWwLDZJyIcCzjl7
htpTQxiIvbsW02KMrHNe1J2zzMBfKq/4+FepRGQeZrqxHTQERG5vZVVkl5sLnXWNkRv/Bw40XOR1
CLxtttb1zvhdepreTMvbzzhvJFbvSc13q/n4PL6oA6WXFqQw+nXw0pR0VMyGQm3WY8mNN5juhFqd
ofscVtsKOSkMcENrBGgKInopap010bHpGRasGMrinZCERPYGkXt8r8F3crMchEt7xNOcj+WZm9mZ
0VaaAdyrUkPRc9Q6aitPbJowXmoQS0j357wHM6htr3veBNKdxSlxpVrEdFSPT9qQJAxfg77fa7IO
q8B7tBBN5rGK0wfccFMh4U8dXlzJOKkY2OXCUbJZ7snysep/qKMEnTflCeVYikh0c+7EhXKU1C3V
WP9HNabklwqeqxbD+xAAtWWcXL6VClAdNPj5GXFz20JyN6uONFIBTnNJ8Ub8MUO61YdfiVEOl8hC
ADnXtoRFNo64lztmBTyZn2afQycCwWSdNyt6uJVeSPGjh04M6io+yzYYw7VCnH5rYOtBwwRzYTwp
6X+8huMAgt8+7/hyXmW4LjDHjpo1bt0Ul3Sbc73QWpX1tmnJVKKdFP6HTBEQIo4jAzMEa1k7N1CZ
OFH/nrBqDvliki+BmMYnDF3p85keLIe7bkZBIzbVqqK6Rk1wmXRumKajJyf3qzu7nKZLNJa1XbaZ
75H4R1j8niBMUvjPPcCKhzsq5cEGQW89eQ9eqnFheg+cXPuu2PwWwIjWs4mu288ukS14fS1OmfUW
lldXNPQpsP/Hi1nf/tCE8qzWW9vHTqTXjh0T1Ayr5hRYkdcAeOM4+qO4RFy/L2GW8KJO1NYPvLu4
7MibgqGYvHMBiZNoxxV/ANc/o6RnLCqdW9n96sBOQ/tusMViM1JYdf+hDFjDtImMOf4gPlmGBZRf
4g3iMc5RRvy7XLfd+p48jid7EoogT2zAmr0k4bZlgxD9AhnqKMNoLoZfIsDQhyNoRGLZxFnkqCNH
//1KFRlgrK1Ie9IHv56zo5ia5B3V2gVmeYYivadiCrtekuzjp/30qso+ucZUqXb+NA8kUQKFXkHq
muv1xGN8NSgAw16Opto4/g4f/uOsmJsDzh7yS5eov++Nthlt0pd1CD18Pu4u0lOcrFB7aqpkbfNa
ygtHlh7CY/cy/d4l0/6QKmGdgSoVJj8roSmBGVzn6QXLR5PcMkS+BLuDRnLjelUW2PVOtUYP+9/H
9dpujm6kMVDmiJh5aLZ5lUOXYMZQg19v+DyBmfl5LTEI6XqDQkfaOIznEzXUrg6qtPTAFIy/GCvr
J9JEVdeHUhpuJkhwu7E12SxNUBmM20VbSuThjkK9UfsebFthyOR3dzQiNELGPv8eSzNkXuGBB9in
JOIxYNpXpHQHbz1qE0dv43sExT6nS/w8BIdxdJ41+lWNaH/NeZ+YHrMGMI1qFOZBv5ArK5aXZVk9
Y58DbMqnvx1lNfDjxdEOYeqxgequAGf0581hp8HANv+Z7nhwp3ACkcYc3HrZpaQ/odX7qYOHkLQy
U2antSnRkoYzWe+JqzI1Ulcv87amOXGfTSCMocz7m5iYRFQ4EOgMi3kfhlb0GVYiN+EL//v6sFUK
onKkH//0Et68qjMvoErnSosd7AFNdTTjDGb8wiwJv+aQ2AE5AOP7KAqAUK094JymlCG8tYva0Dbq
DbvM5tUhL9ckVH4MjeoFglXhTRYgaYR7s38L/86jtcsqu8l7aDSCS+H0QT/n6ysx+8lghJKybsPd
wtSF4GyYmpp9ccnNSIrYgZHdzT8LB2mxrABG1x9i5zWymLAsnQ9VNw3EE6AjvxFO9tVCfI9IZh17
UNDsexe0vNsne9I4/x6uEcK0v66sbbjiIXovCPX0Y+aBRBdHxx1IT6nqQvXsQvYnUXhOXgXOt26Y
aqdkHBQtyTpUC5mmSSQeaGU8Q5TrIVxWG99LOq7/d4btRGD9tLoKfJmGexLj0+gHhLMjSDXJgCxI
cz6C+f0SbqfgfdxVNl2XQ66tu5BqE6d3BHrrVRV6ZSTdu5A6upBWdfPUZSlBpdCYknShTwXdxXN7
zyvTsio+VPl1oBJYQqEbsACarEPexhmicwzDtr+xffL8GsNZ35kMl1bla5r0YBqP9JTkHyUoJ7I4
GY5US4wNzi4wtDPuVCRh2VRCo/FssF9U1ACeeu7jmZsuFO+wS5gF2KD26QAt1I86wpK7m+sjn/Xz
bC980JpuwQBFtV1qI3XBTWdR2o1nV3ML2pYlLq1Pz4DavXN3Vv0BJGM9dwoz2qq5P9Dya5gW+Pmv
Y7OKR6/xpSZUkwCAoeK5X1wPPeTKgwcEmtcOh5yCvOs1VfX3STbXUgQIyHYm6TU2BczEgmnCkvLh
xp1SGDBvJlLcNSxcyXl4Uu+VGUFrldob6mtpTK1jVmTgBVaBf+b6dDVVJflhFGrU03K4fUjbhsgQ
0mY4rNccpHflYY6uwDRDqSPQ40RtQiaPs5NZ9InRLbNdFl7RUgwzC7D+lXluhWkR+XipZK0cHMnw
3pue6MRGTuBzrWgMgcDuURaAoLreDNwUL74F8FFNXECZucBE1Xj1hS940bgMr6Bn5Oe1onx8qj/7
e8RFK/mmpH+lLgHSAyTNE22oqYRTdH68zQKXH7fxtAGLv9EkNvvGv3x8F87rRlH1nIgUiKA+RhW6
1I9KVfEx/m/BtkcplDpOGOH/Y2eRvR3SSxsClN1bHQ/gAqDY4Bs7IBf/IvVZihv6sg3f8zMww5J4
tJtUucrJTxDBa84wlZNLnC8B63lgdvXCpiHzL9kn7l9thcPE2YWpkZE5k2kivOjk9MH6QbCSaTN2
obWW4aq56f1X/ju1d5i+FyEp37yTS3C41vZzjpxM2oxVpUQtUKF3lIE5+0Vx70ApZGzcDtK9VLOO
mDqC0nSmwk75eenTciaJ1ds4FJE7Ke54OrazugSB2Wkp8POZZXvtvZjD4GKFCJlQ7chpo27eTHbd
fc63zl1a5mNd/qR8rwOpU5mgvZo3IkgR1eMm6sVWptKJjoa9X1iqU+W+vUIOL5VeygKekwJRukv0
lUruki4oYB5e36ZkrN8wW3xdQgSLXSsdWX4iCnYq4bC0+kn71nhsygFbLxFjLbd3xO+mzANutiLn
zrtSr6rNn/tvMka3UkM5g7Yc2eiRMVTNV7sVjWVFkejkKuNxD9C4luRqCkWsCxnKqKvm3s4J8hNw
MffS0MjcrAtS9v9607hmLpRQ0iWb1bjaKGje9+r7LvWyIlJ9nkRy8ni8M2k9xAxqENfO0E0zdJyY
equ0cZcsixMyRC9+aF26ysbCOfsCIiZdgRktaX8U+gIpfJYR9gdsYaMj1X5nMWIySZMSiHqwafXv
FfYgvZchIWZRMpV9O2XaojKle3Skm7UCFHqPBE7dgX0mC6oVGREWyqmbqqudnmZF+/R1nO7Ew321
1E0WxgZ0s6XE9RKvBpmtd74nCZW7VfOaaJOzvymuQYVdyCQlb5jnebBvCq0qigOSafFduGrBlooD
W3/psFu9GrVFomS8GAPdk2jQXC9jSWzWoPU8eH9UazHz5rI2l77OUlMmUdf8g4u3+YHXV/9Lo/M7
CNkrFFwjOBLZw8JakHi4INk8flO7+0qwgkMKsP3qNfBTjwXlPhI6O47uHYkqluWOQvjRG1+xvJJ5
HgsZvtsNDxPhQoiHU1xqRfS+c1XmPBnAXYxzmcog73kVlwoLxUfYX4AqETOauUOpZJfkJyr2aeU/
t6y6pVjtYDZvjyZiNGQfkO6KOta3lc+8VhSmM2MDnbM4hMuPv/ngjH19azD9a4njm+a2Zf453dmv
U5soLyWh0H6vE9+/w16LjSqJb2WJdy5nah7QGOZmjc/3bGvVmnpW9YuaDp7l+6l4wVO7wdTPbrU+
l6wIYteI86tB00B9tI0G5isyOyljzoL20lT4ee1T8evNXD8ywZ73fFj3j6ZD4aNSsGdnfk1JVBrg
S693uT23qegN31v+6iSEQnwg0GdO/vA0w0tVyAGtOm+AvMSjK7WR3UezpB742s/uz5P3AEmP4R6n
wuVafOMEvvmBiiyyiCvy7cMLM8/9VP2EFj9ditz5Bjp1litoQgC8QI+9mdGdieKIWIRd1lZMg0y2
2+zewjRvmlkQwWdehLiVakIGWCxcMskrfjRQIMZJdZkEc5gzj2eCMw0cG2jRGUFScIFhUGiPYkNp
L4dBaQgLnBFXjp8BNGaO+pj09/KHCkXLvgCJZx3D3JV9G4YvNvjco9dGA0KA0Hj/jNK6xIY7Gpjh
ARcIc3wi1dbGfnCCaqJBov+xHs2rid5SDMvkJz/dY2eso9xxJkIWMHDZ2SsWqzP6KaMMw6SbD/Pk
i+sYU9gRZEy2AlE9kWRDrg8mUms+2VMKlZPqRvOmscO68VHMKno9OL2y5f56juqFKi6JYxAtgSt6
py/qdS9WQ6uovnuHKYOrHOaEKZ5rhkUFjJa+n5ZUHA/VRitPkv5X/6eGFmaqR6KBziWqI7ViVYI4
AwfqthtyoPjqE5chE+INDg5PpHtc85rECo4Gb+fpE+AxGFqwbRlTOIrhTY1bw2ZeXs6xejPZi4tO
SBzQbuzFLJIW7e0buWEN5T8AYjO+d/YYj21pKjy5UFqjvGv1RUv/kg/YyGTbn2pCQ5UiRSiWBZVR
1zspxRvV5BtJJfpr8GuX43iBrWE2ujL4iHjDueeFoHP3mGXoRMYbaNxBXsn7Ks9Z+eHvk+3gl6us
TPJ6vLEaKaSAwRF6x5Y1PtjxvAHjjGaMsj5jBLZ4xLFNjBaqyBVt4tWKt83TvCPCCKuoZ/5tZU5d
q6FD/1RsCsLBbqR5nZe+6VUhveAM1VECXhr23WgIe2nB3Y+EGaD6qPWhfknOHrRAIYn/q+PC5fHp
hnX0JwfWVMs688Mhck/5+zRdirVCLw0rgG9eH19WMmx98gz5OCAbVmFmQF+2vCFQVJUygxwb4bvk
S77Jlo/DULkUgwBxqF+H+5G7i93ovzPah9GQxed7QoS7Vc8X04XlmR3ll5s839tb/FYuVFbWh+XD
+l0SA4QvzlrABnP+f6gZCUclVrQZzhfHIDuj/0b6FciWqmVdW84u9YfCUHjlNloPiH+9oEuH3A8m
Su5BzpoyEKbHS3Nlam9Lfbmf99xpDN1o4xosDvQWYl+vKy/ftrN2TMitAMuAKmmXbF3cWkYNRx0z
Wt1drp/wAQhkm0Bc2hmaRMVprLmxc2HMCrnY3UPSfcWHiBGROCoQa6U7OvkVRc/q4n4rr0ieVvhQ
LN7SxJHjRlx8jsXCUoJtwezomJuwT552nBwxiV3qveXxnO5KY02dlXUxuI+ndE3y58hCs7HTq7In
S7RFJTnQo8RmTTj0rC1m0o5k/dYMK7/H0mK+P5oI2PxAf2+eGJ0M/4AMqHwTj4zls91jTzONb1yv
QIjmioITrxuooB+beG9xWnuJJESJtwH+ItEloaaPIn8VZLCmdXAw1qoev0YBnvqrydKvfssjjRJc
YUUNvPrphCWt5h3lLyaPUmk5QuurtzNrncOIRS1he9rLSP034ygCdE0xRIPhuFnAWX52Ci8UeOW4
pW/ANE4ULfft8/YQ/U/ZvigntjcWzYrYCj79Y1z3Dv8Yu03fY527krGnsCfFkaetodRXhQcHnC6C
R/IwbA44t3VKrk41REBXZRl2o5hLDSWwBP8UWxuyp9SNxZ6uuycIIHj6ddDkswlE5mYz7EnWylr2
hXRzMhfB0ayP5YVk795SRm1tNvi00A0/xaqc9bYLGgU/epllwltucyN2SHArRrjlP1IqUa9FGw/y
eFxmtb2pki2f/OCO5wrE6II2qTbhdn0y0y/CdYZ+BIsfMEf//tz938l5m9zMzce3Fs9NDsploSym
ebIIB6/fYhAu918nbgNVY8pCyM6PpNXrVMFmM1fz0GyWW44WTjRByB8kfA8Ahg7N7s7C+DRVHdsP
m+hmEhM9DV+yQkxgMxI5ylnHpmXJg/Tk/6dLvXe6Hcuw8pVzw/KMUpb7xzTV0NtoOmS53dmpvR3s
pYDMmoOfYK7GK12UMOQEty01QOeCzfSglzKYYyVgRuw9vHHaFxxP5cmfcD1FJ/eTx35EADHwrQbY
3lA0wMLIVflgCbJPwUBAuXAgPNoZbBDFei48g6ouiuPTsKbqNoL6/jBGoxLLOU26MJpCeVIGGMgQ
mO31POajOCRPNTlTBQNYj4DahhgwMH7i+Drjj2ylzYmQb2Ik1tECx2eYzwgj1upBG5WaKMplEp4B
LxW537DDJhEzaFHZfocQ6bCJ6M6/E6jlkeN7swPOMRaztjcAj4ympre60ni8JXN+3pEr2Hv+D021
bHu5pfwXrWEpFOSkDn1GKj3OqCFix0FFJiqthRuuhxPZxQM42BCy5v8QxheF8G6iT5fqaWJTlBSL
UA77wEib98YfmTaDtyUwI8Ju2vVPfkTnxfOK1+FU8DhYMAKfINunADo2sP8/7kFpRg0tMZmgILUH
oNQSYASKRQ7vpm8Sryz5UuX3bI4GMeLjiGEJ79MkwlyuDBFvPn4SsBliQGFUROH/UCHie+sMZvks
PEtuK/hvTI3eEqi7bJ5xa7NQkdWIHoPtbzr/90779LX8/ipnV7zeze51AIJ0PqG+TNVvBc6hAoab
6XpC/kw9kZn+lAy6HyJwABrhzNHyBmECWVzeP+9RhTQVrVoJ472G90WwaUgMok5XFV1Dw0vuvrYi
/ELF0AbJ5buINkdkM9onTL4lpmTE4VFhUe+mqZVqx6RARIn9Ljt7z55NZuYode8xBibUfCQyHYPu
bUCDpIsFtiS2IPCrN9kJjdSchnFh8HZ8g2q70Pevd7KLen7Th5/EjkHBqRfkuN1bnCln5Pu+261x
lB5dOdCWxXm42NBm9cVdU/OkY+iGjmVX/H0t89/pKLJJswBBTEAHbH+zx8S9slVcwye39oGjI8MV
MApc5eNrtvXL7UiQ0u1C8RfiKrfObXh8pheMmLH0CsU87s0qapFecdr/Safqrx6arIES3OOVStN2
SqkcgVkrXTCYphJSDU1BmrIBv/ZrkOx/HOSTwquWwKF0QkKc34MYpuMhld1tRvzxh2yvPj4fQV1n
RM/vaH6AwCGyXYOj0Z94Bj1jj3W+jkfOd8oyu++73JCaGXM/S/C6uUWJc1VF9RKs50yedDv1FPFI
wOsfupBfz7LCnGkTB0RMZbI71OSswGlfC4Ad1EcIxFR6QJtpbaQQfhXxMU8vVcIUWHMUHr87bH8G
cU4wqfRZAl87asvJV9nUtSQuaXbdz2lMS8IEzp+eoMzFUzyKvVdDOuVevDTjHl7LF8jH9xk0wGQ6
+Si4oS2k4osAfv0Vj097JFKL9o9v/XcQq5NWYfO4XfY9hQ5zyq9ZlnDzSKvwf4nLeAhtU7k/1roJ
7o7Lq6fWqFnYYIYoyS4CmCuwUIPjHzuKjZy/lfOii2N0zLZTeyiFQPz5W6j8nYr3PGetmgY+pQrk
gHbK07465kXk1RX5AsdkJ5fNmtIAd2qyD2DmN+vqDki6uQJG3Wc3NyH67XYEKWP2pZru0Ei075RD
b4LSt7FzcYCjCR44+JTkEIL6goHOrEyVLDTCh25R0TmHC/V7Z94B3gdbz2pwhG+O9kCJ04Pss65+
LRxJvAeAf/ubXu8sXu+sJd+KW1ivGwzgxzXCTUohlKw0p4ZsV61KHoDZYHZhyfXT1L1UR3OCYdKj
pPrpGHOhFu6GnNcJSM74MH3njvw6VfeIpBrDmfnRnKDSSXbHnWwk/VNt7QgTyVqC1q4d8xxf4Shp
kUUWmeY37aV6QwAl+D+KcBnIC3Iv3kKraxxjRb597ySaBkGZbSAKnVXyqq/FRWzMS9quz7Y5APax
C4TbbAvLzSDhmB2AUD1PKMxBWCb/BlZSLQY/BClo2zB1Od5i+yzW+QLzFUnPq38ualw4WG3IxATc
EgnyY+8FQ/4oc6AN85DX/njkW6dPZQRX4Bt8Q2ksPwxqMdSyB9Bp8WKBl9XH5/zXqy/oEheBFl27
ax6RGaNoXVxe6D37tosCk+G4dGSbOLVeaXGC09YQOEwXvl2poneEN3UQ5Fu9YZQXrQMUhxvYY46c
Zm5N5ekFfSLl8VVAzPvz9svMyUi9pjLhUGjjY9aSMvCZCtxKMPT1PPPCJ1Hn/jlnjosmaZqJZPf8
zldAeKJiiRFc/1PiZyRe5rWS6JGCKumWgNPUifZfPuLE+/90mzJRL8kMy4d02Uu7kykQlfq0PgWX
vMBBfjx+6TAxrTUsAQTuzZWVi0l3sjE2FeVGaZf6tM9+rxk2zXEp/OX83Nin5GuSJbldXTub2aoK
ORXsm1ySICYyBmaLcb4Dj7TVVjtj3iy6W6SyM/GM1KhU+Rjrg2kcD2waJcZ2+G5dtsmeL9IIgwoe
3hWLYW0WgLddZgSMiUDx8IvQlN1cmSe9PgEPFf9Qx7ZHVQl5/FiZtrymUr/MmMg3QP4W3Fe5dY+K
IDchLskJAMySw8JTVkKvgsbkYp8wLYr+/sQVOG54GUma4xVsD68iOR8Z09fT2IMkkpRLKrLgmiz0
ATYQ/rO48XAJst8NqKM9T6B4U/c3kUJVvs9X6gYinysw7B953yKlKu+87LZ9PVINDGpSy9nMnjyY
WsGWqdYzRyY0e1v1ggnI/XEj7VLfrWFSOl82WtzMkfFNil62+sZI+F87Fvsond9PWAcPeeRlNFxv
Szu23DEb/nDrWaugGbaPAMp9u0lNsxRJ1Oa8chPpmKxOW5nEmaCxs0rPdC5W6f1A23dmmPyrctwY
ZtUQM9nJ/yHA72BVHEwrJ8AESxYM0FtVYjQAd/XAj/pFiA3oxMiwtgSdczEXMxR5O5Xt385SyHnm
QDQJn2j6UJAwoSalOfZ7A1EJqeXCK48x92gIWXkbq6Qmmio0IHtFIRkhFXSLbpDA1iB74ifDJy23
qm1A5kJGtpdDRydmpQE+wJVCi0OqwJrggTbpLQ8bHcqQ/WJB5BhbyQk0yDACy6GS3TWvmEqE53KI
hxjmIBlg4MeIfBlbrZTE8Wn11/PcR/d/C4sa4ImSlUjuCvqEf3qZV60w1G9Aopu6CdDpkTONegxl
B0fn35rn1Pi0/DNhCiJHqdHqTjWIzv+RQUqnaHnJ0A3MfG1J1CIBQ3XWiIfwTQGnyQK2H7A6+WSr
FMc960maBcadXQp9LJq4fx5Gm8krO8AGDP13pTrTeQpYVQfoDf/mlbrJY5bRO+8hp4T3lu1s7IUJ
XU8WOUAkzAQ6deljyg1g5dDkw139IrYAsOEKbvqRgOwknBeh7qyCdqPnBxLgG7/eyOyMsiptWaTu
AXlJgSqeNVnWyHbG3cyi01YVaFDnk0n/LZFm62dX+TTynFG9keQIv5ce39CQgV+eXgqJ5nlUeLQU
8FTRS1ch8h65kSGQFlzZSWRCjpYLlOqTWvfnbJr/F088cWhzIoJ5FJZyUrfQ6HDj4Lu5z2jC45N0
bbUWPdMwaHaTFTQSez3OsyS7HHVHt1OOX+rV8g/CjPQdA/V3+RkLT95PLAvlD4q216S/Q9vazlI5
mw5KCNTz7meMCpOlfqLMPkVn8wqb63QIPADz2MjFy9jwDnyRKB///Ik1hhbwZv1SboZy+46NVzU5
Fl7e3U8dBIGDw7d178SG+Imd0K62bYnoATCeznQ4A32fu3kuQfWISzdYCrs5XxsPp7L735Vzn5tL
L5PLUuabjj9AI9tJxsqPyS9qFaIkZ5Qa1quvMpHYxdeBDmBNWHIAEUynW8cBXGPMvN5cbUWiZj3v
YLmta31KNZ8I3bWtlt2wY/ao1WBPBk4Rb3p2Q1b4ylXRoW2Xfzi0Ob35U7bpIdSBUEJyTdSvLfMq
WNs7Wc1KxV6t5ez8yyWWfXoTn+WbJ8z4Sm0eVNFXOD7RqL0P+bqySCMQ8b6KbuvIQb6UPUw0RyV/
lSxYrpdDOhX9Nnff72xvEBUlLEOMLI9VupP8hS7F8LVeqIIY6b9qfOZ4dE1S5RTiSOEFvW7lBhmT
dHsQGSlEylbG2w0FmIb69Jd0oMkXOLhYY9krLpDB00IOsHx/oTUqyIFvxjQbBu5TgPytny4WXeJ5
lAq+NbLa7GwLsQQkJsLN7gWKG9SNwFpl9RyY2vt6NmSoMbfrpy6WYnlyGhr3FdPV8Ge/QEJyqSXE
Jct+BShPefu/aWuZ9Rxu7/WM3+CsgPDoT6fTjDwNitQ82cwp06AZJDrR4dXoW9PmQS3dimL0HrGy
PC8LFziSy1U3G5ogSYzzX3Qa5f8XE+Kcu+BHiSEy/xiebsv9W3zb7z1yKZfLVvWT/ubFPoM6FKzc
Ql5PQ+k4igAuROqCAGUbVvIupMAR3Ffb98y8Vs1sa3uQc28w8qcZBbXLaQB2hWeLppTzKFjRsNM4
Wu2dGFhX7M8sZXG0INDhuE7I/IdL4kqZVQ6gdosu3BBaS0wiIegEeCq4LUxrYwKKCa19DfO6A63m
dE6HG2+TI/Fx5s04Ly6+hT6UYc4xR9fi8xNdqATBU6ojTRVlYQhsngbDzMhj1cnZ7gTkNCaonyru
+UQl/JTfLZ2pQRn/BolY65ETFnsoQulg2SnQzvU/YsTtSjEqfmYRt9gSQN5Sz27qJ+wOPJBZLi6g
qPVGD8XfOufvuFuVFQgZgXM4ibMVdonP0mAelGG+/NBxZY/iZ1MOyH608R5IUMmjnvRImK2iajXg
iuZm9RaR5XwpGDbXozQUuWprEiwX0dKouvEbaiFQft4BEnbN9ExnIC4MeguHLmBDKAfHeNXVmHRE
3TCUcUVPyly2uIoX2imNPQrssZbQnKDKG6Nejvh2wWbInPfyBNLW8LuFKK6GKwBipIZv43lOgX4t
1qcjJ8AXztbZWr0BIAtpMTZXqF4XDxqvzDWRWU52SBG0R7n4Wap6To8coLXnL2pbqb+KaHreHTu8
fi30PEcdBfG6xwqlCDZIR0ZjTp5wMlz+Z1eJRAwSJg0zphvU1O+4giKOiriJs0ZL7sfyGNGg1467
z9QQJws7+yfpTX4LnjI2sULfKdCUarxSEkjBFWtP8ZH3q6QrvntQUHWvR4wS2kAoxODpTXuyjbdN
aKKPSr60q68jwhja00FpIN6vELJXWK4mon2BewtfqRWfsaFnA1pDQYeF4l/yrU1XXFrTwPUrkQPI
BLVTyfug3OwY/uzf2gQZr/c7RYAT9TMLsuAx+7kQ0z0Fiuh6JSd21g/Ydhvf3ELr/6U93fmK+0s6
LOcYr4J+ZS20Iotd3fX1EDQjUnFQJPF8b7tVsft0r9urvP9hN/Q8Mw5zUiuB42l1nNRHdBqmKWZd
eNkSHdJCSRlgWOCV1UfC9gFUHe7kSVKL1eeSpoRYaCrZ5ipZmsNMkgQp7bqhT/MPcPbrNdj78jY6
QZmipbOsaia4gyx55M+wQXRhNE4vmXXRM9Ol/NZrSfQgp/6J5bRTzYFdP+8AvNoNDfrcDHC+VhmC
TrCfUu99j06oWPSLu+BU6ds3DQ6CcvE8wNL2dyL1KmHvN3P66rtWx0nSgO6a+u8ysyG513tLdgnB
ze/OQ79Xf19pL9ZqeNfV+3Je6oyp5L+bg9rwUdx8U5Ul9PFLn+k3oMhI+d/ZvIP3T+uYIJAFlFgA
k+stOGkeb3Dkmbs15d46i6p9uU5jE0MMqv/eFxcE2gGIhfn76GVzdrlXOx2kitpQPMEZuzxBjBIK
csBErff8d1ZSOcdKIfeTWvI6QMgO19SlDdTy9DdO7WyW9ojXnCAHHksMPlYrRcQpXidZCLHTXLdq
xzrZualMJBGaoEtCB2u+NI1EfBXX5NytsschEsZBnk+6Bi8KqvJubm/n0CYiOJ7sOXkY9eTM1xg9
wCSAq6FLVfKVMsrNZE4raKIbjmKL8sxSwnyUQh3WIxhYO6/k6gUQGmqs3welc+ObypIfVqX4nRAQ
gdklIgux+ryfzDxdruL6G45XTCRL3RRqw+oPN1FtGZLai4iR0uO8S0q7ydCCYv+2ev8vajPdciJX
/k0zkptltxItyEYnO8E+NPpsskH9HGxFX5oLzNEYSX7SXQ8+ESFTWeMQfKTa3DV39NwqiNt93BR5
fSMmphV1G/B11uFbRj7FT+yjTHQXHZ76K8R7RXR0wv2q57JHnFtUuuQ3PlCAlWKRDZX4GfMEkgpR
qWKNX7AYTF2K1qUyBN3JyuYw6ZvevGKlEe+vcJlbFLz1v3zHkfz9nxPVRVOFq7Y9TOCHZVcSCC0R
MlkvML1iKoYq2Y02fdbfYqBAlFAuwn29kGje54YU9bga1ctG+Mlt6Jar0BwSIrAeHdJn7rdk/pg7
MypYxBPcA4yZRTY6fdhsXGiH1OYyM572Q2huqy67cvnINP5bYcxOQfOolZKpX3GIQCrKx0oUQAx1
dFmJPA8l5jPIp2lEBZptxMy8CMY/SmBdPORrMjQgcm/2wOlfju6OX2uPuwxjigsZvH5kX6MG8tZE
ainyJqgddxHw0xE6P4TFYY5fWwsoDXsXuqlJheTLnd+YhXiwTS6X1z5laEK1XfwJtnC2I7pV8GXM
OP0QJQZNoyqW2CoCpHNP1WF2w667gQ7GnYm2fMEBQL48DVPG44NO6h56ZanFUZYg+Xyt2bp7nwys
kFIpDDEyLKtx1BVU72aBgiC5QWbp13VGZt9FxUZIc3YPeeGDDmXBFaSfBYUdhPfFoxsZSEBD44Ee
n4apZsr72DZ3XA0uJ36cKeDUSH3MNDOO50jBoipogTuQiR/3UA9M9ug5uxjKSXOVAQudyKLnYNID
XjU1Jeclf2v2HqgQocOC9vt/nVmcugXgqPd+Awp73WpOakjq0x3ZoI1yrSdzF/46PyrQaxfGUWaU
+S3SiWHNL8pR+M9y0LO9mODnhZBOodPBe+7ky21zrB/qf9P2OHxbuQrdnROllYiRhQZfPKRA7O40
j+erF3Pc/kt960b+q2dFm0KW2bgeaeuOWxeODEEg1u5vpHb5lgUXwwPhwUkJtoZvVDUTV19XPllb
6Kj5yiyyfMmKZ7kD5gH/la+g6RxpxPLluWkfgQyn0f+nTHMCHXpSyDSCoyH2GOyhh1DJalkkxCpq
IwBNW4KDvBr6KkbUbhKB/vRrc8Q0F/mq4H0SiLWiF48CTRf6bddOXjWTd39gcCFrxs/pDyhHDIod
+EiNbrKI7baGzmTDndnv2706bmEjmUdQfmS5yC/xEmj/phbguxxylPlGTRFY2xGVekzSia3Hgoi6
I7fFZw6yWqfJXBuHdyPCrtYiK7DTFPU/ErEPw5Ap5VkA0QWOxFUJlR32ApJEjzyUDY17qYVt13RB
i7/YGyht9QDWDViAJQyscDjGJAJN9F6hMns0GL/7uuavIpWNjGc6S37xKoLRIRpPPQ4FHIsVlCGN
/Jkesw2z7GyWB7EYtXTm1k45ZrXiBKr1ErkHg5hdpneVsnLhFgVrXVXD0UrSmWB9uEHitgIrBqc9
RCLL1V4Elq5KzKgAxQHt+4zDKcR0jcuau6L8ftw5zoOr01vkACCP5Svjs9aU8geLbB1z/uNqLTie
uWi4A57Hr0v9tdyLCK+toy5CP9UerL94cYry7opTJgXv5/y6h2U47KuXrbr6JeN6sUfp0o+MWkQ/
dySoo5uZpMcX1E05WgjyHojrYMQ1OjHhSj68Gg2pphzhkX54q82/h1wg2U0Hmz/+0fdZxUbo1exA
U8U4UOteYhRKLJcOeN/2tCLDYPqzMgXu/tioqzOxKo0gnnNarmkbt3IO15dW1HG2r25Wb2p9MHxq
Mh8SJtz5BdF437ZkKpzl6U7kjbh2qSNQ/KpqKIwTLWSWyljzE8vmdrwvko4Z/gax3pFph4DCv1HD
t7frccMSPmGb5mVMgl1JL869+BQV7Qb2qeuLGxSxwOgeWbZhCNAWvb7DwXytQZWfv49ycN2FF0F5
thZKkHSFy6NGhWRkMMeurKntZYHp2eTUKXCC/bBTfWmRRDdE8n2ck4yGqIaDVnyKSyizJ6o+tTuQ
jRV9Dvern3Hmqb/PY8VU9dQywPuIRsU5XSqfJEm04R1HajEOLEjxtH1Pm6M+QXxpq24mn+cdA1iU
8jYoT8Jc0NrQsefmUimQKEUBu/p/vXQJ6509Qf8b1JpGGa+dBYhOtsHiYMdvQjXecUkCcl6+xV2p
LoU7cLdyQh5Qo+Ij/CYABMWkypF7zsZEQJtCCbJdrsmIBWQ9qD8dIYVb6OymflChqfeyU5dafnzJ
Cnm2WH8vXPYDdRQoiyYjzJhojJA21zn4iYsxL5ipa3EAZN9bYfRS3v8AeD7swchl9WiHocxYji0y
v+S1rESlmd8Ti5hYDcp7Z1qekAwTSXWFZqx3vfKdKA5uPfNRUyaKuXCUzg4CM2GIcRjFlr4fPdR5
ruY41lSh1pQHvx2Mwo47Q/CIWk9Sj4xKUAE5QBjsciza9GytYhj67/oWGyjGqj67aVTWJinV3ZFs
zdkRMp3UmUr0UvDUOo4YfIka+uwCUa2jTIxK1H3xYA8ZniMHBO9TWCVgSzj7pT8xmWzi7wuUP+J9
fIGOZyEU4aprrhmPYZBCW2Ohz967tys/UpZCq03SBPp5quVm0ub/9asaUNmseqrCTTy1Azl/mTsu
ZGgRZDEjdnfvzx40GkbuCttn2ciszA59zqs06oaMWXc1UaYFQrUibXjhhgZMRvuI1/zBNl83B7b5
JwlMwJRbK4+aLz97PV2KlLFmQtMf1ZP6iVsihHXdKvzM3AVlvqewC1zn8aHONIUt1B/42+jUxi5b
15Ztqnc5q/1guku8DAHerEXRp5A62PNCebqUTZVVWqKo5AvI581YG88lss1Um6lpPNDIsWEMnNy2
jM+hoDzGLpqqPWy8UCjA7k6/L/tI+ISZkDJbHzwCjs1jaNzk9a4WBnXUOmUw1PQEYZyIDVgH5wYz
IbbGUxFVp6QK0lm20ISkZIJDITbYfjbx8z8TtN2+zUPrltwJEOiOG+RmaV5wJXBLkC+prVqHwAZr
kKNFGKDzU+c38Q/cTkeD8DhrRewCJ6xo3KFAWTeIW9ek0lMQ/VgdS5y93e+L6NI7I9UThsLIqaeU
oXYPRb8DJHK03XonR1U3+yYKjcNuODbF1YcSpNUpA+Re+wo8gVSmWvCFUamdoHI10pWlm+xb2qQf
49qvI3ejX2w1H6vy6DhKp0Ba8bAc8Xwb0CK2VFic9SFFmwzteo55I2+l7qdgjANzYjjh7xLmUUFj
YyKTaMvosB5Xz/vRrjmCVJ7zo0dCukNGWo9IhLl4DYP6OSHGysLEMWewNj95sLDXq2DjrHfrFKKz
v0L2qZ25oCFHNtNPA0CnhT7hIfHymTUb8GIUCy0f1Fk5wGxqYRmpg0fv3AERY/Sp1S11M3j0nFUr
89qh11W6z2zHUlunWaY9sqLH7RKt5vT31eP3X5z7eFIykFoWl6TQr4ZHqdBE9/0jBaRT3qdvQO5i
DFzjz97BNpcefmtDXkeH1Z/ywULTLRuwvQT2V0CGv8gLvbPvVDf0K8pe6JZ00sG+6fPIhBNprdfn
xG7JXweONiHTIMMJKVmslaOa14hwdsnkcx9VgQGOSyun4S0S37p6VBSziPAeXC/cAYYlQ68GFb8O
4wAROLutuNtfR3D3SztlBK7cHKsL9UB7+vcuNnnoIMXVBFEOCj/2MP5u3/fGy+39crYDgj06uLBY
WoPqBxXsbchTalOwWSLeF1LyC+B0skK/4doXL6pUth0VivOMDNeZlTKHkSt8eCUqn/Bo3rupKvnZ
Tb7xBrgIzo/SkwVHW1LRezLWrrUaUZaPSROyhKbLzNBHFPcCj597va3CrJwWstJ2OQfIs9mYDE5t
ponTCuum+PP0BbBipj1fbTUMvIaFVB8mI2FsJDllOXsHijPtr0HcP2wxsQLhtgVoMCwHfMLBEps5
yXO4ygczTP69LuZzjdoyqacjp2QzrirF/wUUYbcCLh3CNkxLxpkt9gFHh5x/bCytzYxA7Gz6VQCa
rEclwjafH2cU7gFSFlKODMnQVXSP3939FFc2BSu1mTK7zaS3+Z2gKatuWxbxexqBuF9cy59ctT58
mDWdXpGx2LPW8OBtJCJrHD/lsWFSE8fGtVV+jB3qPThmAqI+uZ0N/eBe6HUWdpTU27ZfaIkunh69
Z3+B43H0Uo4yJ0NgaYhn7BMsJ05WZ2lwr3s9/gIbOMuDYiNj+KYOa6m89w2tC4Bfk5r79HSTv8mt
29QQqHhm3/SPzSEXY24H9ajEPzQO/7Bwq4EJm+kPSN1CZqJFeyK56bZgPN4rJ4dcQQg9nIGh02gK
T2sC15+0aPAOpv5G9K0bZHN/gQl8zakegaTDE3pw+ima8jIo2+eAAe080sUDhPWDlsvgE0/NrgNO
JEgA+lokE68nIAF0BvseHGKOXK5eaz+lmGzsJZWX/z73T9hgtjMRxSeeK6XXJrnbSyCe28+ZG7i1
LpjZnfGK4THGnzrBOzK8+pl5l46nGSNuXVd3oy1iF2BU7jzxMJ51rdgwqSppK3OEOeIqCFI8dz4h
sKEIuwcOQAbMmT2prQcS0nGd/TtmYPA0lAye7lFMXaA1BL9XrgtKI66scuLIQul13AMckpBkaCpK
60F2OrbBDM+qhoo5Gs6Ij8Le9NlGo23Gdc5JFuF2NFPOHLIVqR2tiHGF4D9E9EYPfxoac3glyfIn
uTP6d+4wPMGRlbOH7ohYRniDQjVMaihq62lEtdoeHctBkwAW2KvGgV08baj7DrtcZMmJBicmfV95
PeOyIE/r+xWlO0g0bPAK8UeHH6fjgk5GNWSCBbpjudDtM0SVPMjvmPriD/yXfuA8YMXAXyYwLFuN
KI1V3Mhaskl0doo0dpPPvSNtSs60Nitmg08iIy94xYsSkY3sGLL5qrd/6ojzSVnfbVVa2LlogziG
IhAgKKRiw9+qg41tuKErCObcq+m8ppU/5JxGoap5UrhNrQJ6f5NCmQk47lKXS6mlvNS/R+w0Nii6
3UxdT1pmUNewvNaxW7L7rOvzr5qx5GXGdtwRJAHjdh39xo+fE4aGm6OSMKn+wamPYDXhYCGf/Ig2
TCK/cqxECFnKxk2qmmxwZFc7U8W/3FDIW4IbD3lT2mtbWLQIPVdxaGmaV3fWxzlck5jqqDeXjFAY
xBTo4JLaYhwe/wzgygTZ3k5V5oxz7UKPmcr7n3fOBYEpzOHs93DtlmCtCeySFTe06llcJeKOuu+r
8ktXCvaWHDEwEZvniGmhhoKlyZbD6wzQhDnVBbclEMyT/hsOHDyY5JrmXRjTz6ANZJQRikWduDMu
ruB3ga3fdS/kuuwQdZ1rr4vHOYYiRh1I+oVt0PcT5D6r9uMQ+tznjBeWv9WTbB2LfCGkD2tRKw2G
MyJD+oTDMzVeeDMxT9gC910txrFlgF8FxSRfbeZrH0lbp2OnUupDKNr4dlvRkXT5LqllQ9ODdkko
ZFMhetCaMeHT63Z2qTYO7WC6l2LSvcjfR69R7MrMss9I1v575VaPrQmfKQtI+sWUkYlh/3XPfkHB
lUD6Pub2d6l+f9CYfLZB3v5StRn+mFaEOcvTc/7eh2lwMSVeSdBvJKh5FU76QaW3IYEcMFfMU/k3
8n5Md5h3PrmXAeYNNVdp9azNUf/tDP0n+Azk/P0eQBLSZgPs4u/7klsiqW+13RIt+SZJ9WKwc6MN
lFDb3KahL0ke9XkPfz/YokUUSw0KfQONc+2sI7i1b+s8nXAxpjxgmMTuM5EwTue/d2uSz75mKWZn
iyBErkmkvlHuUuamFjfeeuqyEu0jJiEMzrAtn1M7SsMP6baqI8E1srIVLvFyFDS+6Ap44x+fuV9c
+UxkNIuzLug/rTggUuTUUew9JmaycA92U/Tt3I5+/RC38kG2q81jJkKInR+mkNFOP1sTr48WHkAt
WFdMqAmu1IfwEDZCAt1QCGfUB3UxP2rSBKbgQA0CFFLt5wVMGTFxTa+UoHmwiY2GIo4PJi3S4KDO
Ws7sngQypJzdYImIXFoDTmnGgJNl/t2mKNXb8yxZylzTbEo7/rZ15MD93c8EFM/aOrxAN4hVDUc6
GLuMY/ApLVe9RCJnIinZBYKa3MSe9E0gdbQcWKAJUqy7vie/gwr44EIAfSZeQtlFs+2RPsy0rM66
grNmKf7v8j8aTCdQEj763LmuVJovtj8gfU4jbHBjbYyQHTH8BQtP531U8o+6faWeEVuO92McMuFx
ARqngyo1QnhhMqEu+EaovveBo5JMXC0T3ym6Bv2WwL2YqcMzFYo19mGxXq+0pdKxthdE+BGpW8od
jBZo71yzp+N23lE+JhpEnjLLB8Ll/eX9gGjCvH95VzfOG7QXeoGWXqYWAX8urwaGiLJuuSwinvAL
C+rT4ubt/Ub1H4K7ZTQDXYii3eGRxTvh1Ox2LKSCLzmEHWghczN/Qoc9dnJMPyMpIkuOwicHOIXX
iODLRfj3qyGCcv+siiFahBmWyzVH76HclJi2ZRqBMnIkV/7JEmC/anMmUM4JZhslRePtBhk+AfnN
ql32cgqr2kKaWEJ7X+JV6Mond5yLF8pgEiJckSw85wRJGaSFT2ZZW9ujrHso0cLIPOPOCcawzK2i
A0DGjke/I3ji10mRHVOa6+liUMb1iLDqyNpbpAe5B8vcsWrHRECcLYXeJLbxAG+gk8yeO6Zf+qwU
/L6U9YUhoAMe+PdLnaPTmfbkuyJ+z+2Q8ZS9TCcDTsxRusRGkJOuN+JLtBrJSWbYoS3alxvLzNf+
oplDPAkBX6KxtL5LXKZzG7Ihs+0lRborIOhBtBgHpao=
`protect end_protected
