-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Vx1P/Os3LPZB3vCBKX61d2UxRAUmEK8WDWecioYQ7KXsiBzBe28NxrKgFW81tXpnoNt+9KDQcmoy
UVBxBgeGmxgTjxiMD6/ehg1ioAmOnKB4KICfLiiWccjXNVRGJwBrTAOcj+GRHABohlU+HZzBj/Xr
FVlxwTMdo7QSWoiCNUHpX4zSufnBK3PaSjcL3/vFrFe4IL/KJZJAmHuRChfuj4tB+FkiW8mQEyGX
TzF11GVtXlqMoysYEM4LQqYY8nd3gpj5PCOwRv+nb3WUHQgi+iFRzp6iAawKXJgzzr16L4NULd1U
yXOpp5nX5ZeqHhGWCq+9pAMW97XQR1nfiw25Lg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
/ZIVsvsu6kqN5xXQbLRj2OeidGzJWcx5b51/UlmHglcS7sQeWIHEGskUD56+E9uMAmHepLhnMVB3
QffrXSLohV2Wy51H/nz68FQFgM+NoKeXhwCz+wDBb6qw+EzjT5f9ogv08Uru+Eq66OWOIQl1nNtV
f6OQmwNr3BOZszrmvfc9O8LqoMB+c0WWYT5OMxxIDCRDBe1zTf7l8a0FDi82skHM4IRqWB2EPfrW
simYEqcSnclWRWO/tyQosrgoHYiObwT2xXr4wqfjiyX1H3is75qkk+KXyMWf0x7dGebqUs643agS
6I2yOqAetzk6Rc2C60kqZRZWQfPAYYQqI90WV7yzEcdaSwY+jI6fqj431SCeIggNgdOu+2KEaY2I
6PFXRGdWzywyLMPReIvsk3sqp9poSW82aSq2XcwhZRghK9meuzcJlJ9ydSzxqGFgQbYVWHMMa1tV
PyFXlp0eyIi1PMyWBb/tht07Z7EFKOnZgJHiRq8v9l9jSdhmugzShV6Zh6G2ATG5FMS0NwPa5K3F
N239+RoL9e77LtNpqZUSEo2xQi+ytwKI/SSvcLkzrvSMoX37KULfz2crdYC66vai2BF1NyFxrr2P
6q0oH5Jz93rvMlLRRjw4snm6rYWeTsGLHl9LFRq1GT71CxgasGxGBbh7qICdFtYwb84Q5TILq8Oe
rXPiv1rRUDiSa7GLx0LLBLShfPurFqVk8GYxYRZqPOkhxjU79qC8TvO1kiTz1a3Vq3XGJtV8yF4A
YRUDdAmXmRNE4iT3y0airnpiQj4rN9G8BNYAR9V/J6X22v59YV7gpBeaWnlIEpalEWci7C2o0NgD
VHQ7yXdpP4DBx4CXqSPgAX2R0tYJxsA2hvLY5I45v2Edrs2wrUYOrovFYnSU+0U79s02gOQ08IEO
adGfhCrFFOaAK0HKMmk9QlTxipeI6vjhWaMTSmqYPOWPKw05WVtFCccarskhElYBFplKhyN+PH9P
K06LQvn2VjE86tPtPD6YYKts9DElQKFNsePxAwg25onG1XOo8AQdhuqCpPTxDAquw5YW6ykvqlEQ
zt06ODtTqkd1LKs+iFgF9ljFo+aaq9NTdBpnaVsk/Pzse7jzhuAHDZmQhvAU6tlZDUCkUhk0gj/y
6KBtWpr3jN607ldvvYchODffeQPMjewN0bP4QV/gcea/8j2FpW0VFwXvuzlmJPlXUG31PtVz6Pdo
chGl1CIbNsY2NcApFJRDKOuMvp5Z3rq3B9+VkrqVpY/8+iCIAIRBkqT6EU2pIzyorZA3bKqTU17O
hfghOrpWFDjRfw/ULESwOb5KatfQbErqodpiaa4kOxZmc8pqXr/OzR1aGwfyy2epae0HFWp9oRFs
YGKxBlGatChye9LglzOI3mXAxX0sWcpJIqtkOojrfuHS4J6gKPIM1qnJB/lDtBRCth/LvsR9WDs4
b5NZ0clJ1ip+nvYxpF0m43YMI72s2aoUANCJ0aAPw5U4F+TJI6XWdT5sov4sVsdxHI5edjbdKnEz
mCkINaNxqA5Tun6CXgBiaVc6szP1ofbrnb+HFaIgkflDOg9N2jGdMLv7GJHW9EECoogkbqk0NPri
GCPPa7hbPHh2/87nAl5il/5CoJiTpITycFZ/if38AjhcygWlEf0PnqmwAaZ7sWDe+QArXeFHLtoU
O1QuRQ4Gvpfi1d8reKWd7YXCiBLyOyTdAskEbsS7vf5gNBOe0/AvL1EmnxZhuzDCwuCjtMFbN8WP
S3GIbMOOd6KmYjXKDCCtKrrM+WSLUSn/7zvARYN0BGWcaQ41NVX2Gc7m5g4sp7dpaqirptH8jnYa
vF/zetwziREf431C6LUWKPCcgrs49KqvNawwVOouk5ChDjUG8Y0CIMUyx9RDllfsHmFI+xXrh5OW
E4OLfGrUtAZP3PvS9QPw22sB2wuWSkvSdpj5hOHdkOrNu3ZK3gL+ukfF6X8KIhoUR9HaSMU7Wle2
aVjXo/NvJv9AVa1IRk9r6qRPNK9MsQeKCAuACV+jLLh8whA1F++18+VB43K1lxZyCoKFsgFDbdB1
ISb7g1tbi2jMNtaFnL3CzxT/42LI5MDs+5CMV2stUmSXWc8ll2Hw8W/8WFA1ehhkwyn0gF4q4ooH
M3qE/DryHYN8KgZIoD0IUmc5inNO7vpIBnLonhl7wuHk8SS7HKpaRzy+7D50UYhwUR700GkQbfHf
mdNojZ+8g7XrzIn4ldFKKsbzf3NrB8SUuDbXhV4JWUE8fOh7rKLEQDmMKqnHyrzVW469BHdHUamu
m6lYYcVAxPAwudKvN7hkk8qQ6t6uDWvRjzF+v+egpACv4qjYLq70D1ghtt0T3AAj2gw4HlhHoTUe
ZmnQ6r6wmXlO4nPT0dsK0wK/J8P/7Iv0ufuP1v4Hyg1C4e7CxKiRVMmsGGatnZLx6EwVb4nNY/mu
s/gBQ5Qe4aAMg+U85xyjPv7BVNI4LX+c0fqsoQtULxdH2kSWY54RP3hOlWHmQWZNLeYEIr2qiOkJ
Sj9DRMWFyTitslV2K/6t0q2fiEnMRvbgQuL562ItQFDVciYnnOBwEAWuflX7JCraKoa7HcXJqBWz
OJckqCBqBxBD8gnCdvboerWYgr6iFifyP/vS1dJ/Zf7yTzS8qUgxBiU5/+ULMl+kntRx0HHIWpV8
6/OMyw5lzIHGj5ZMQghPWKuPKe9P0zGiG+57QBbsOH/2Ptxo5Rxd3/Rq5aA4eWrrYPInWvwadqd2
wXON7q+BxxzcCZhfXmf4LwZn5WTUOyVfYGwBq0+BiwnBhIusUokILCavVPP+e2PfH8jYrC5RSo3B
JzQPOUw4S6KfN7f3gD4JUDDsvHAVygUB3nUap9D/VvTuabWZZme6D1QaFzL82mTor7rdVy42tthj
O1/zKqVBd6HQYCMvxjWQX3yGcyd4b21wzJdnDPlNRtc60lmOpC0nWicicIwbMaP2ItEWpLqnX1nW
435AzYY4KBK1ZdNZNsrzOw0N1UjLG5yoLACyHe8yVfeayt3AHLlGPlxzG4iBsL224GR86FWVE8dt
uCoQOJby0pvXQ73OshevaDHPtZ7XIXTgW7Azl1eDABP/AzXxXb/WwtSYVtWJGojZjRYWUnQq0gY+
L/BU7ShVJvNRRRcO2OcBiArnTolMa2esWQGBYIVTQXQXwNADq1TtqidPS1rgBhxRCyHfT8xEcTy5
0Rq77O/Qa7VGJ7r/28ELVez04BNvc+VRcE4WXj50CQal96QzSeOAWxEqZH6Avl7Scy5fCIcIM9ol
uxQyDEZiX4kRk3cjyXLgah7tQBYDy4i+HIbRN1t0KP7SDoqAilGUq2/6c6PoA4jF5P0wpvalqrjP
J3dstmD8PqarWLyfu762NY9NsnYuIRLg+Y6N41asr06TLrp7UKUVRlfYV3r286hIEbBFcU8HbVOq
M7DnXDGeLm7Iqa0VBicnjxhH2p17pc+mVNK7lXITHcslrj5ffi2Djglim0xcYEMNDlAzmW02mhHq
9aG5iJKGKmFDy7Ybs9/J59aQSXCN+y7mlZeSHfp8vTtZs87i2c+6Uc0MJdiKv3kSVvKs8CjbjCjv
Qj5UgpJW/ybdFFs9Q6qU/MVRSdpObuTvDCUfpYZrnvT7temYjRGHCB89MQ8bwlwiVEhbQNFG5FnO
N9vfrFYG/w6okWKwnxtlUgY1E99Je2225FsX46nnZn7fnx4GcBEartnMt6b2HKGNCUMuHIf2ZrhT
Qe4OYparA3UChGTcY9MTqgmvKBfO7o9Jg9GALkZm3ZdSHxB5N5l8hYi9QPcaiBOCRiUqGMYoZcrZ
rcWb9M1YKrdz/Ww2u6+K7Cq7kwgwR6x77r5VAIO+g/dmqvH6wKwtqRJdRtAzGCZ7uC7D4/ikmE0D
Y7MgaM4tqrisdMOR7aGF0VlLcIt6WOv22LY3Qnb3EPfEzSnmiIjgY92lXO+G4/Z5G50u2fW7aBWq
se6ms5wv41H36b2phC6IsbPaUUrYH94KKpXa1ljBJTx9toYvgnp6RIUUUhvTVB8Hvl8rS0NxMrM9
Cr234BMhNCNltvKssV0cttyE4Hah8TpslwoRy6NTqBCR1aACLg9XVp3oloxj5Bc7e77whJ6bpydr
cPG3itWqvZGKWkhd0hINAoLEe2DsbktYfkPCXODCwjjjkQBXas1MC6UR9ZM2X0WN3m8nkA/VQUc6
pt7YVFDvnMMTFJvpG858A5fKe5zVVo9MhWlE4JXOpKV9So5d46U+rRVuCPXDFwTnr8cdlAUBXLJX
23wwxtJGSZ8yJ32fDNMjmvUMbbuVnWExmRgvVyXtAXmeiW+gvojzG83ce3kCy09GPiPSShAmwumf
ZGrcrwrvsDJmxiK0oUud8jhaDkhmwbWoVugxIdMIYBm+u10wXZ5D/pfoPHbpTaUKgnMFolHScZcL
HseCdSRHGgmIAXHeywz2L3gsYryOcX1xeKBbsoDQSQtkDthzHUPGw90G0Xa11/Nj2uzYsn3FMVRt
Gr5gP5DbPEg6Z2g65+iZs5VHn2Xy43N47VX2XhFdZNruOeR5Qb2lSvSbmp4Q90CoIXvQ2CsdBihV
c5hZtySvdDuGPDtGS57NZOEvguV0VcRAz0uK/6SPylaqIeE7URG5pj9Wr/mgi9fpr3mnebhCq8gP
f+T+5ddc4newrf1cVnhNqnbtOZr3O6XHKKV15lRtPfm1Em8qpFRKUdPUfVh1x9QSgYXm1NsF+FVD
rWsO5aygKGCMOzvyYBcX4spMn09FzeakWdmg98nQthCvcDoTvf4EJQFWkYy6KU+p5Ix5KfPO5pnV
62TGVTI8TYfogipuHwJDPozlAyCRPpcWoqmvBm/RDP5CA2bsuES6Rrb8SGkCxaTGBnqrTBh/CP4E
erI1wbtubnsLALMnmT6kW9Yj2BlW3IxLv/gokaY+zp8zXbESNVvbO61PJ9IqOOc1/JSfZF/mfSBu
ePaE7CDy3fliBGXmeZNIkywnmA2AGQCreLbpLmCF4JKXyhwBnBVx1o6WhmR61e87B6jpXCv8Dg4c
TDghSIu8hDTKioM8jTKForWr+LchbeYGlIiapz0RU1CrNHHn0o08aj5qBbdljQ9dL4URzTZ8UzQ7
S9fjS8AkA8XAA+ja2tUKH96sph2hbv+xMCghgRNd6usxjE/dGA9rbSZ8dTkSDLxC/Opzo107bgHU
J/QR0SZPYBWC6J6EW7sHdpayADr9cYbT2hgVgHDqraYNKx5VwGEoZwTOr0hHYLRMceF0afEjM/ea
577KgSeI61rj7/+KIyfWELzEpZePRVOb5pajjplHZY/60P+084w+6O3FPdphxzVmlaYc4WWn2zC9
xO58hTqszpGn0kAU0D9ZYmdFu9HIwkGnjTsdYp09GSsrg1Dgi2TI0spdWFDQljhfwcw1xEuQFya7
EqguCb5ehIt+wq8hddCJcuCxSVvQvnCVvYsduB5M49io/vrpnia8rfKqIoKW/aS+Gbx189RfPUxL
wMwKJcFCPi5bkIFnvmpPNokC5lt8kJqmDcK137Q1RtoecjgF2CqjYZTURMCIywNX/q69IJ5JE8qd
4peQh/LzvMDqT+EC13VgK9D5WMVcmB0RelohOlTvWO1HDal+TklXLIMgIAorflPDhuuZxNA2tV6r
TxNYAbsRmUn3sMQD8Cwks9HAZtP83SJ5kN8IcC0xHTvI+c+5JW5RpdsLGO0OkjwXpQLeex4wb/S2
4qwO+m36j+xIhg3xQZNT4VA/yUfXXP9Ch2L69tOIZJ/pgN6mRAyAllaUWzHld7X/72/etJphdDsz
XYiJL/q4yj7hEH+itVMeUs2SCBP/4injIEc1BVpvY55/W99BP1DW2T91/0gNljpmoPoxITyN4kXm
46mjUrB+1ZoalxiUohkH6aF9CFkkwNehLa97rrzwG7GV/1YbSDFbZkHLNk3XYNcw0VGcbkQeQMOw
rygTqL8Ro5c6L+J7cfooJ0eeK06mtGhZVVhGNbzvODa+ibb22CYHIKciDCxrnkPNXQp7K886sf+f
xKxRduyNcJuFXRmJAaAy0keMoZ64le1ByaigDdpqjlol1x2/7g7aAsSSQLXKzdQUgk2wJ1wH2P2b
j3UzSLL/O5ek9Q0KR7pRLlL8OyEWzMAPCtDXzLSCXvN3GZ/KG04b6OJVp181PGJaYf2RIWp9DRFw
c/llYZkMAlJNj7U+S0aTOYG0VAWWNIt0F1wSg2nFVjDVTQTkc+uY/8PhEHBBk0HgA8SMFV0DDyrk
pi56TLnmrtcooKtakutQqLFkrCq8JN0Jb6/BN3RpMIHDZcqkWWWroZw1jbqj/LYaYknh98zRwS73
vSC5cbG+dYy8iQ4Hs3Z8/y65STwW9syrv1E58yWrhSrwmlAI6m5TRb2lUn6cLXRKe1Yn8adAeBbB
Pv7jai62a+5eUO9duVqMNjiSweJ2/z5CUXIU3kDXWKvszuoWvxVI+UpeGi8ypuO9EqKIvE1CYr8E
IJCYpkrWs5G99moG4WtGERN55FS+OHA45ACVGXyUIdOSQmCTsPOdaPH81r7XF5VxXQ/cEd38KNT/
qIEYiAp24xP2w9YvLONwqq7tLMHocbf/+n799/Mlqh35tIOiYa9X5YTa5lhO/kmq81X83T7nl0wr
3myaUMCiJ0esGe9VH03e5V4dht2Fugs18+vkfPJchVCy0sQBAN8TxNva5wq6GQTcCIxmLca57PFn
OsJbFM798eJKCcksfEzz6vk+s8FPJB8B2e7InKgld43la50p9T/kdeT7Tyi+vVVYgv5yRHA9QyQo
cBp8y2KsgCNdkpxMkj4umxrxC1IqNnz4Kl7giSY3IsL0pRUIafhSm3UcoIh71l/Rb5G3sWI2DV7y
1fMdpotHLCK9aQepyXo1uaQoEW62Ar3fwPycw5ZsPcCNbKDr29BdEEqVF6LpOlFcYar33N26rE6x
/xkwD1OAjWzj47RaaY3Bw5YAFdlB3ERZqvooC0xbthA9WIVjsdWUZ4fE6iOHcUMIdRUy0fpi520v
hSZNd/GY03hR0b+SWnGBF2g8kjQY9eQ70h/zn/+Zaf626raLufzIUuXl11nJGWU/TgqmuqhGcQec
wBRUolEyC1sfADgJh3YGnRc9KIrM9WmZ9jHcwlK1kBGFlhdaWGO9eBTp0wOqKGIlg+NsQCnekPZN
a0DZUS7gmMxsftex38kW7Z8YNyxnwYr/HJ5KBH+UI6idUegKX3AOF2UDlH6g6HpyaUMMyPb9KKHh
i5TkE2jAH4+DmvjffhbsQbEBP7fuC+rFWrw9F+omfMJFfy2czlsPTViFMnBo78NOpo4N43RQ65XT
FJXGAOSJ2KHZ9q1FBolHZMjXh88+XkDL4FJScxUsXcOUahmJaT5tqekmHJTN/f9XLSaZMkD+8I4X
kxCuVGypYbbbYhCHS53cvv396tRHXQCpUYMe7XGfYgomveP+FW/PSdIZplcpcc0+oKnODrytTXCJ
cgyk5qUvvfJCXDn7Qbp4g/Ocb+7w0/aILWIOSeZjgJNJOiPJtPJ4ZD0vck2aDcJTlLt+7TDF5Vvu
ZLXyJGpbqFHc5+zNha1OS629JniDAjCab12N/CCp53Uc2V/rD/2tcCRH2/dFF5kJocEoUfBUtbrz
nEJfTOgO010XDjThRDdewhWOpvlsQABHoxEC+SiuNt4okXWuGus8y5pMlH6I7K2OIdE/p0ZZCerm
pRRUSNBSMj71MdO5WqxA8NKVEoYNbJRRBZoG3iZUtOISHL19MrvARXxBVMy1FbcXKsLlzCbJdsb1
V8WvUjo6IKvQTv4vLKjlVlBPApuVe2+GElDb4iDvhVHxA1wE69FcC54ssHGiYSCo84PgeTUCu5h9
DJYSlcCrO28wok0qyVC46hpDTuA6R4MhcjMXSXdUkJnLGepN01lKudez7kLv/+BTyeCeR/oPWnTK
Uz32g/5jVLrnrcrlCDb5kkB3SHdIa5tBbr5pZgErhLaz7gPXPHsaEMhODVMBp1imOvryTe8oqd5z
cMymB7CiRkC9AwDdshPRL3VQarjAmcsLERTXBNSN0gJDd9dpH9/XrsjEcEU9BIMIEWz52XVcKwSI
7sYJ0vJlBrEF0uFrmzpALFIvx6Meb1lYD0yrPYIkDqEn4GeWTCyjga/wLoaFiT7NBHXPvkR4OEyu
4Mf6q6aphwmOZXwQt2KcTf98gChfuNVYJevY00KFbmUvEEJ2jOTbo2l11+N0PGOTrWrgWV0zqZHf
4GmV65H0GKD7kpsBNFV4pO/4HPJvK3IHLSxkT0kMYqQrnXX1CRxChXpbpcbTSdBSbLOY5+JX3gL1
ztZqt/9B5IxGHFipSd+GXMvlDkoFd7+Fbn4qFWrmwbJ2MiAwvodHXeWQgcprIxFboIUkdXqkJsTz
3ebk0jNRxqpHmAOR+82OJDjKYcTX1gH+0xR4qd/CCSwUjjpnQQbZUKamXMW4FMPJqXW5R75f960A
BOyF1RwggHHOtAEg/OXWAXArT9q0f99zoTNVuJEJvmSCtnqJ3NF9P0fK3KDjDHvG7BA0lTTnJSGD
GO7FAYXgg6t3BPGXKSdIA6OghGfUF4hwe2hHK+To7pAqrAL0jAnDpq36ID9h6U9Bf4rz+ljM0bYO
NV5WVbkwE5H1F9VLCMuZ8qq1m2SadpbWkBjZ0szngQb/wFFOqyEz2LgO/NxQdwmRLHlcu8uFMXwA
J6Tid6V1vOb7xg29/HXZXxQTYa2OOOtRK97pjy5l5HQ7yvPJA/exWDpBwHedxen4lKRlq09sgu9Q
lRdINtS9ya/6oV/KnuoKYZbIITFRdNazOeV2wPnCPak5FC2QzogUn5izOs74LiFq+N3j6Ep6lt2u
mkkK+QbhQABZvO8hVq3TBhCxoC25lRHu+CGj4Oy1hEb4aIXKB6w6iyLpt1iWQxdmAGoYo2mf7cue
gfaSlLpePR0Q3SgTg53gYvvTA9ua8bHvfbhJwutaAQnyGP5Yr+pOpLxpswQqogZnCxqaJ5FjWsrA
evwD7xHeuxY7t8pJQBDBo/wYUC4Kr2fJNR+v4rUKDk8HZ58TuaFOERIo6oy1ufz14AINapJrIsx/
nQeq72BNe9Op3jfGd3EzpvaoV4g11LrRuGM3ftHVJGToxsma6AeIXNduT4AWgf9pJUM+JhPupXSE
SynssO4Hr4kQY9fkMEO7/TqcEV0/pLjXEixZyT4+SUYRVcGjCJrbNLBtZyvGQjD/c/iH34OlY2Pc
/wM43eolvmh/e/gJ+b7tQfd/5iV8AYYYo2KT2t9N7DtrN2M+kkyvvN0iGGNyaMOuH2y2rcN8Cf01
6iWvtniKjKb79jWkbwN+sOOKLeb484732R10ZUtxqPK/xN3hToKgmzxNy9gIAuRwTmI0OoctYHSI
HEOsznKnUa1iQD2Nq17wcGt7/qEfWmglB7i7ZkHPfG4gJ1Fir+tgZKmbUXifpVpaumap28D0HD8r
Jq1o9m0S6WqmUgke7SlP9KRlRJfugSANyxwgp1Uw0EsgnNlklyl3Ggnau8h+q4C3loZp1Z8zHkUa
3zPCAhSyWpGwXb3zmL3wMFXd2Jk5x2JF3mQb09R7UR6iXOUoF6CNjn51gocCmZhtYlWTa5S9pZN/
2Y5tFmca5MdXfn9V36E43SxE/eEHXtVdH0Sip/04McIuVKdN+XaWX8xYHHJhiMZo9O2YFCUX3F0O
ukyT9cQlvlLgr+gRGzRgJTvDWyHzQbaUJv3maGWjd7OaI39fs7Ea6WO/jrYk0P3KASz0zRvYQyXj
315OUsoQYhpc2wsikT5u3mg+YB0y87zm0ymirdbf9owjyEDFd3Z77YoEx2MPA9NuYegbU96DziMF
PIrTFc/YWJK4g8DWHvas8xKs4GGgcsIEzYqMW6B2C7bwLcsjKfblEjesUniLEkp+apycUsyYLrRT
pyRZjxph3mrGVfAknCrtOxaIUC818wTattN5m5Xr8XCZ9yN6uoPIlCteXoqSMpbtAjt0J0b9jYlA
n0vlVcwhC9NojvR17eOHgzeoiGeCne6I/K6WAgbtFSXB63P13CXpQ6UEcRnr92vjVuJLb1okiryU
SxFLQiNh8WnPZSbGKDNNa59MHpcVljzv7xuqQKb6EsXaVedxcXciypSjSKuHYS0j5Iz7WKXkmpew
XzvGOQ+Fg0/PphHf+zh7/hHgf7OoVoMY6EN8Vyc/0kkk75IFegdd29PVhU9euMASrTfqBJOi0XyQ
oJOiKY3Qy/1YNTowlF2l6f3lfpi8cfocOmkmWbbcPh8hSbUP7hbpDWQaAoz+1kCtp0EhT981e3SR
okhaBh9va4qkmGxTKFIq2OOVpINuUlVkbp0MCUz0FOqFOmpd2S/ID84bLJZmiQaKmtEq4Tj0Xsvb
cbb7+c8vrLPL1YQiFmVCVTRWeZ/v0cordTiQyafMvPE09q60zq0z0Qacx94QGUBXnKEweCKaDqku
ku4v0QPmomvtGMNE8CHZTV/aqCKoMbHS4VEYtEAv082cFXaEZ++GLsCidUDImnGFZ6u2rv7uNrz+
tt5ZggWu6pFLphXecvmutZxurHrHpKh7fuxyBLGSE5qeV5UcXZqvtuhY9lNjIaFdW3eGDUgOFMGv
lKJR5+a4buxOANvOGcvgNAmjYI5PzG4CCX9OgxHQlkxGaMSNz2IN/bkrCPjfFvMZSvXvrHBk+aXm
BfN3qO1WdFPBS2Ceb3/l3wTMa+sk31aV2OiClazYRjkU78Ss06gFF4/720GeNpDg/RyBa1RSuxo8
/1x/XHyLKFrkr/dSwVQgo9oNTZx8Yl5v388v8ee5WDgwL048ufLz5d09fzHwjXw4ZDlmm8hJWZay
6ubXGiR5G8GBx9m2EeS4Ye9VDf99BTCzL/XUChUJbz5tCwjGJueO0C1+Ex6DVoeIWtclz9t7VRy9
2sRRR3NzQENpX6T/QNAXxkjbVXkDVuxfCYuamllyPI2MEKiNFz7Lm1gVoc/ZrwNnt1Zl0Wad/+Y9
ecgm1iDcqQdtrb/qlLKTO+lNUCg0JpTLU1t2ESMvNjzasTk+jD4/R0oP/y3NH0G+2M/DC7igA/mZ
Qn2DxWLNgSY0I8rnw+TZDUg3yVys8oy8DM2UFEAMES7xpjnrDZlc3DUyn16e0RS1elQKQwU34/5y
jT5fPsrsG/+UZIfgYzaeitnrfyaLuxXQuZDlyRi0fydRIAYmQJ2ePSktxg3uIMokc7Ekr6+aIkMH
hmBBQwAVOZOHZYn05xUmvzJxjevuKWCFVeOa63jO79X6eQKL/uiXSCFQm9HABQJ207tbI+kARoMJ
Hqz0m8F9B12b6u1P1cLX0nrT89fyoZVbQtubK55tl9B+z1IgAYhOk0IUlM0z/U+i8FwF0Im+FKZS
YrFiMyjB+p9+vsD8QgA3KsC6VuF0UT2Kzy3EDvSo0fECqzLIuIo/QNcKjpuK+TnyetVCcSvHEbjj
BdGkVxCtiEFOSGYFghOkbTg8LxLtENupYDC6dlt/5aXUzLuc6kbeOlZ1Hi/Uz8cP26KNlP/ZFGw0
TrDBMD22+QSuEgNuTQAAMBOBH+wo3Equv2x8+fZBommOo/+gaHbuM49gXbF9dPa323FMUFLcy4lq
BLCcAhd8OECPwnYF3gtMMFDLK5Yw2sOBGB1BSb1JQ5TkwTnb15Q0Yvc99R6VFsLETrJ3i0TIwV0V
rd+InkloUSwKyKdNxuaIbT1paocw/aGf6uP8xZkOVzZBu2whsV4t8REhXBruFJeOllKLZ2QEQ8w+
B0hvNUEGqPkn+mmj0q3oS8w2+uvLTRuwXTe5fv6mkuiNnLbteWOZKgB1dEuz7OA3xfaS+hM+MgKL
oEBPzC8SC6Jr58DYBZosaHc4SYS8sPpetcvyEEka/mlvl0BPcJ/V+DpCeAXi8/vhjqtminRODykv
74HyHkzzoMYqLmBV5gRic8iHTt4RdWabuLFAUDUDyR3ylZ0xoUogArDXKmxWBII6cS4L7X4VmRUD
KZPtQUwIebnx6aaqJ/83bjzyOvt3KsGerb9wYMNoaVDpzbD4fkim/DQMUHqrc880QFN/j08dpRFH
0+SKsMAAV7IC0Bsr9Mbt/zD5ED8aBKrNpS+nv1KL4A/H368Ct0a14elznL0sCN5yjujeOWMaKFdR
eo4QFfQXpEQxzmiwUZTczjnG1S9If27UYB7hglatSKh9b341OarCsj/xUHYQ9UOr5qvLsKJOyKTg
D6GpHNWPDF5mY8WM/44ZB7tlmfAVTlSbptaMEXpsbvgQklAaBpUlwT8MCek5hBLTQPAVGjuU7ldV
txSJ9bhFjsV/9U5TDMSsgumif1WXB6lv/ErK4PKsUK7vAgzDdPxOMMUZPGveoA0h3058E67S/365
HJcqyERn93YEuFnz1fPr5gzOAVY7w3NNPUnAHc0uJs/cVAStlGGUfMA68gwKyVp0+Cm3g+yHePm5
SuvV/JgZn00qnUMIOr3dyAtpr+ubTT1pdmmvxU5esO+cljIRCxvEpIboqJ9DuqYpTEapfQMilKWb
gqUn9lFQz9Mk9D5ru0Ba4wuwUWLhDsKmMvq9LCiBfO26VMS9uGahiAVa8RHoIDQhOkburSUbWbwD
yrP05zJN10nUY/gx73ndLLqhyoyPjta7BrPOEn3hWjNNYGF2iU3SJhHtFtYHW9N2sj0wZyQsDHoN
imG8PWSMnvvvr+U4HG8dsEZpzuESc5LkcFqG/pkzc0jv677qKFitRO5tYxhDQDBeq22RhyfroXdz
6bFb5wbGBH9htfF23b17VufUoTWts/hw4kAeqPczXncTGzdeiVuzoHwJ9FsWL8ubB4I3m9wIou+A
9yt101CJm+WknkGdkyBNgEj6VlQk6wvR7HkY9tm09mObThawqewuNmvfEkWj/DRJN8sDs5B1QhSV
U7KPUBNBhoE3Ksp8ZHj+MGRTeMC6c+0Ei++g1ZSu92ASQzFQBPK//vkQ1CPkdA8tRrmqPDjDIWBJ
MUFZqnKc58P8a/7QIcrosJ9UzMYhibhpZkorHjr+GyJUy1Abn86OYEY8ifCBMjzVFvJj3o+ReCwA
Pi0t5/6u9uRYNH3ibxYP+A5KeehgBr3oyDeOsoaHDJcd/aPjy2SjjuQzXbgVlA2cjFAuv4TD/7D5
Q9wUflugZ8+L8rPQ253xYnRc1SABw8dx7Lf2HLZMlTdeX83Mm+t9aq5MqqpT92MyVgTmRctTeG7c
iVK//AFVMuosM8LI5VUw0sxnY6/3AEAQ3gmrQmp/SNasbejpANJ26BTQbB0565jExGi1rLfY1N9y
im3H+bMjCFt4CWb2SW47p2mbPTZeOTQm9LSh54Qpu3xececgLm+HgvTjw3MKEGZLMAD1dEqGw7g+
GZZhkEarEbBfPaULNrz5OwRAVo2cj/qpzhE+KpYnAQqrjEm7mObSrodXRKvjP3sqx92fBEMqOx3S
Xlf3jyNFPe1jtdCEPj1Iw0HtKCPoE3QWOn27I0bJ0zgPClv0ahz5mvzKrBTjSXjN8OesWfQ3+cpn
3b1MAYpVTq9SoP3DhkfK+o2LBG8ei0bUQS+gvag6WnvLUoWC25EVQq7XtXIZitFLQLMcXulQrwQE
JLLYhwWETW9mvQVShflL0PaRVDP37s1bpgvDurDAAcWBmKpqzzdOrT9EknPU5f6+lOuSH5dcMCYz
maDNX02Hi98lvXOhatipOR7Ij800PZnnuQf2/+JkBNxMgLHOV/m1REUFrpee1FybV8QPYSyjIx3H
FesjwnpZWI6nunKsiEEPawFpDSzEqRKA9s7keRd96fcl8eCyFIyOBdNDbPlCWDNwTvVQF786uhal
AdahsSjMJOmO7ewztFW1zXQ+b8EfrjANK0BULxvptVMA2HUG3REsq2BgTGZrNJWeW2AILTxB9/Dz
W31Ub4sGlAUWg9U6JyTUFIRG3JhqPT8/z0WY/qArbP9WLDVy4FJxENCcJUAKcN7yZBWe/SUFo76l
qzzVdW+lfWh2F3VR6uBsVCyhtWSHMG8nPTGxX51RUCYyTXgn4pUsymucvEpM+8CcaLEUdUOZGeyn
yhnlGor30kKb8yCUWHv2yW56TYUGEsUIM/AU5/qyQS2rsYso/as0TGcED2GYQaGCmacyGSIRsBlq
PzVxDIrF12zRXQaakrDaMBEKZAl0HU1mVZJndBdhpw1cmWjup2KO8VYOAHocNe4vH/twZtSoqf7c
h3IywEG9xjHoWRhaw4Mwdiwpm2/qS52O2dYlmyl+Mru7ey3CTDtFR8YyJ0tOcVYllQy9ZIiBbJ3s
+/+4xlPSdNtEVQLVlFoNiXVybrExX/8VPbdyS/a71mLS72BhYBsAGkG262X0lqXXe8DTwcORmEve
KtC1yaqWnmIxIIuUDKRu0NjcLU3Ab9UzUBBGWqq5Zw1wTTw5Axbu/zoHEYFCoXnQe4NKt8jpl3yL
d8MVrK3UQ143NjUXGJAMp1tuetEtUFypqtE3A+hAXDYH/yZYLDM6TQvQPTBiWJrR9tETl43TUWWF
13+lawjdj4j3lDCxUEkQvRbx2YqSDSCpg6d0QTKClDVL1ALFeRMK5nEfR0Vkg2Bwjt1Qd//6oaBf
N1u8BEAcGTkSfYhwfzPptNNV4sgKZlWiW88K6x35JjWsnMtAnJQhirqE1OCWnZac3jCfBWtZNAOf
w6/3y16dq8P9K94d2rUgnFuT1xUmwr7herl0+nO3K33sb8O3Pvh2AxdHxEk1iANgTmK2kT7SHkNe
QM69KZxxYMRgdL3hS4BxHq9duK2YhXXlfQFfPdjR1Hrzf/AeEgiIzQBPgVBrVjXY+OBTjjbO/J38
SfJq+RDsgotFOHYYX4SDF2CfCciK0/Lbrkx5j0EPWOFd5QuPySYWorsDagmwM2K+kr3N8+zYm6oT
IxuJ1KKx56Ths40T1FjWMieXkm4j9nSvHGt4akaZGiilbRDj1XdJkfxtzvva1vhVJMCZxvh3YNOa
4zPdd/ltRQSTc1b8AVUc+kBeIyFy7hNeDqM6elFYc6W0KcKuL+mzgNm/knAQ6BfdI9FAEW4hooOn
T4UcVFX5IKF1Rxf5S2zmEtvOGqfxCVLKDAmfDKcMSZLlbyh3doFqo0fZiRay9Bq7Ka76MFJtDD32
cFZ6qnSRO6vL6yk9FKgCb4rKS5wtz50ydpq1mCU31JkeYEPnh7DEJzTR9ZtTVVL77bqXdPPXAJbM
H2IGly1Ksh3nczLTIUL2YS81ET4AyU1jG0i8cNcyvYdiHaFB1JMYD0nXneAxpebBmi9yzlw3TinQ
NmEDTZIxInxrE4JHLXQtnnC3hFOOXpHCDpDqpcCDSqT8OxvMBXghgn0DO039AhYAs6GU015uMlwU
9D80ZBu7wRnimZ7BPV4cCjVz1YWxqHG9IypfQGqoc/3rjSrEh/DObZUGVEaGtprvRJFqnDHtKthb
A+EdRbRdUuqdi0Z8Rg3lJA/aOmAAjrWZi4mxE2x/9iY+altWoSCcNwcytHFUcnozMTRTdQOkCzcm
orf0Jb20IJgbfa47Ai7LoGVrsr5mpOj4oyTcKx/2MxJPw+oqbrKqd2L45MFkzPt/fMPNS7piS1yg
WrjrSwYHmpsIzWTx9E5H88BEuYOY9zAAUPu6UBTgC2KxvCcAg+8VcRYRDAx15+0AS8NPirLPufvg
qnaldwmig6YdS0d5ApkjG6+YNlsJpPTbg1nXNLR2Riqi0j0C4xepP3eB1no/dksHqwVwtvoQdyCu
jvEIe9D5zcUNTh/h5AHu7YBSZZbazsA4W7dwkxftJiv71wKx4NkKrr8LjyEmbsLZheIlY1HEFqSY
DkRQVWlf+eHtnKsJr4p5hQtJrqMxsMSZXCA1BQT+juMjDw4fkSS9nrGHq0rja4yt9mlzoZy8/8E+
bTB/ZbIkiAgxYpX9Nrw9PeV7qWeW84FoMYS3ikPx2octCD4HyR2llqM37lpYFe6kouX8CGRZRp7E
ETFGBIAi0arse5eJOqvjfLmMc1wSTr6UwosXF1T6epXtwUxPG2MNDuB62XkpYRLGXkzgJUlXSPq5
0aVBxKuhXLGm5YW5QWtWtHs3IJDEUYSb4mposXyvPq7tAmirRUUf4lhrQfGcrA9pNldnXAwdx7Kt
nzMs1Wx59OzbAIQN178XhG88psvAnurjkS+xHx9KGSGwpSLj5GrSHbSwNEXUAEJS3l3fxev4bIKz
OMaB3710DQ/3yT8XN4caRP+q+rvSR/dVXY9Hl3WpOkyv5fNJdWag2bpMV+QsjSasRJThdynxU42p
fVziBHTX3eOshUFWbXS8J47Cx5L6uZVtoVegq93OrBCraslxq4b4lrYGF3Cu8p3LRHHvwLNpsRyi
xWAPzjihPhyZl8IFIU7NAVx0HDXIJ1D81a4RGRcIaRM1QvQyjEYl1LFmPjvoXLXQDHPdYQSR/Cqv
AaUe+g/TxcmvYi+3KQMHpa0qshfx3D4Jv8f1cviD4WbWaVEWbCHNJx6jZt9DGPnhamGvVCh+OjtK
sUB5sbT62vBH8xmM8Fo77TAZz0ZVRR7ER3niroCNI86sv1UerLkXKAtio3cVEX0dHgVBVfQKYqRo
YIxDdUyQVDusPYaidTIgbnSWaGj8lHfJo8wwTemlXg==
`protect end_protected
