
module unnamed (
	source,
	source_ena,
	probe,
	source_clk);	

	output	[0:0]	source;
	input		source_ena;
	input	[0:0]	probe;
	input		source_clk;
endmodule
