
module read_buffer (
	probe,
	source,
	source_ena,
	source_clk);	

	input	[0:0]	probe;
	output	[1:0]	source;
	input		source_ena;
	input		source_clk;
endmodule
