-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qid6Pa6VhwUT2vZ6mzqrhum3eD3GkjtjB93/UrWz7/W/i4u/b8rZu+VSTb7OPmMzz2yA3bAZJWAq
WgKFLlfF1XF7qZvvJWtHIAOaRQiyCZFMIATYDWEt8+PW2XQiuIEp4vKENN66gTtRLvJUvNtm3/Hp
bBXt8Ydri9Rcw15haCpQGsREE7GcTt3RqBUwtAKRlbbGkN76FqeIKifgvx2m6rFo2f9fuU/svp8E
kx9S4qW8s9+xG2enooUJoNFHftO/P8cpLWO4fZwif2Op/3x2bVhIHL3HdMxPrfKwhezU6fzrFgPf
frGeCcn6mS2bphy22m7lOVTGn3O6r+91uw1BLA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
wN/lEFfxOBCW8KFgh6CNRePxzRMwPGxNS+X21gaPathM82zelkrZQ7cTDewF5dPcI22q1cVBDF4L
8uLbH1aQvJ0hiyJBJreq6+1NDoN3QJkZO7deyTN8HH6zhdZ8HB5ncMWlkBuoRusq0zrcVRJLuFoX
Dbp+8vFdncJJFqMJFiiKE65mGcdmPLwLHxzpFu/sm0ftr5V7Bc9EKrqazIjhivj3jySF5x1TW75v
dufktyXbewCSa1ltDnXxJH9PECrmdT5QvwvtqKAdyExRpCDKG1yKiv7LZu7GW5JWYaiW9cQZ6+Hp
WkW8M15EY0uptITcSYPSLJO2EEJT6kiTe2rajtKGbgeDrFF395pDjumURqniI/VCZi5MY6h30Mvh
w5Sn/PuGiSDVgSDGbdP0kBhMqCzrMHUqPaPPS2lF7t/1SxW5tscF0siPUghd3C2v7x52vZOLIPPM
cY9MdvtoXMcMUomYwjdVBqb+0CTzKwAOMeevnyK5nYdwi0+48qiM2ipEts+La21O23R6xokZb+BK
PLLry0z5q3YqMpGfNhZREvEfn1YMcdDGiuMP4ggO2qOeqETXiQzNTphrxFHr7BDkF+xEtPIu0duG
zmdpBgoEo9Nu6yHihl5ZCs5RYUWnP3Y9Z1peyR3FlFpORXF0RPmkTL/MseiaFTLsYi2jcDOWmFNB
XojD41HCDktymVR6fdwry/FcC8d9f5QWtougArIqKvkhWWBaC1/llcxLP2lhix0tTfBGC07Ys4d1
279OI8Qp62pXa4GYqVHIrma2j3fswnWnjGBZebjs9G5pLz2JKJ9dtfxMXwLqt/7dG3Ug7mYP6FV1
2kNLbs9bPaD7Bf7QoMAVmOKRXT27k/aI7AGN+4/f0WFcX0D4KskjSlR2y1B6Z+rS3C7FPDkMXuD1
74Ao5Moi/ld9hDSWrVY1xLT8LD0Kyp8wCoY4NKjUGCTq3L0I5WHOIK/9zgZAetnxoeOUxbYnQmLH
wxytRlYRADw1IActS1Wlrv7AQ95yYygP5UZMyG3dJv/7UZysLvUBEMOEy51PIQYXIiV+aa0CvauD
cv7Qsa1uw4epmf6G+PXSOyzaBCeVnIiy3F3mQr6UZoLQpOVnVbyGLh0tWq9U9Nv6EQlWHI9SOS/x
Kn3jaic8KeTLLeB8JaUDZ0YWgahopR0I08JiPWH72JrqE8sac6Kjlo4MkAI5GFw+bXkPI9HlD+3I
NkM+15VJTTrxIbiDvokjKDIGE2m1fOp+WargnjHZqxWZyXH9z/XmkcDyqjEA37UbiFAwu+nWl/V/
3zZHtQ1KzOe9wminDM6jf4i5bqQ1rsh2f/X+dd1SnUX8GwLgHks8G50FUYO26H7d0rcx4KrEvjhy
WeS9CQdrqaXf0bhm7EvKaA3+Wi0qmbEkXFejbb6XW9yE2bR4yESzMg28BK9okEdBwUEiD4LskXne
8qtWOF0+d1RGzwspOXlT8tW39Zegqf1kQCO5WuNc00Gv5vajAhR/TNRIB1FuN+5/EpUEKT/0t1Rc
o5vxcoUVGLaG9dEOPnNqQRS08P6bBYgr0gdZzZVdRnz+mfmO9ACdZ+Thk70MV+ISy+Z1wTob19yB
eGf9v54rmGF3EgNqIch/+4CDfcHdafg7rKYrNh5S7CDuCfJJ9E74RwC2AaEm1p8SLEPSSPucN4wq
Nlo5qiAyR1YHZLuvN009p37zxiliNpvz1hD1DbrBkJ68uC2aeuDEfRkErAL/FQy8quzTkRRLpuW9
qJ35gCy5TYyJLKPtcTZ9rSQLQemhEPPM9rLLlet1Eg898F+LW0uLbdZTETgfvr8nUciQEUJ6VhDf
/0L6Xm9T+WvPn89IhO+tQEHCN0ZYNs/otKM8Jcz95vur8p//hJbIqDUhDr5Zkwvnab4lKbFMbN2Y
wBtVDhOSLU/ERQ6yEougE6fWWtytvaDq5riAm6nCgoNGixwM70InOxSo/5vvrwtsB3ziii4/AUsw
jniLXi6lsbQVzrwTLIjOHinoCgGDxFRDyWiMzW68c9QyKaF3veoclZM60Lp8aN3arUS3Td0Wp75n
t15CrvHtQvwajf51rRv/hCaeeHDBth2Raamh5D+xhOE9EEIsuvNcaTD5TiGhkb+mkNecqZg0ZPIz
XUIm11BWg/4eqYcBfs5wt5kIudApzmCvUu0WBZHKXpbQvVDcViFQUXWpNDrIMQFvAOQEi1XysDYW
QBpreTei0W03T5pgJ4XTrxrXQjr2IRptdqvX/mITVO15hXgnF7xw4RzkcYP89EQruvBXSviYb1pb
dr/xf/1CBmD+y6nU23ryyd1vKmzYZlRvor7rZj9fAwAqyEl9r1VjpCXwzMnbv5TZZibNOQiPYbH4
B+2m+Qr8DtwdKq7wh3+RiJJv3xV4FJEpqjSmMpMSNIhdIJFMXpybfAGVNvnLWaRNyaiG0D3WnBzA
Mz6K56jjG0JmbTMzPcWJyO04NX1BZUvBuiSTN24hjmRfwBH0BrA5549pku2Lxq/hE5lYnZQqpUrK
7je/npuakzTtDbEvDCGb/5t9F4aiYYCbYlHbTbe0+4O/hQUum3Re6oLMkjdBG2qlQtpw2JZm6/MI
SA3Y36Q/ZNmT0YNhYrVnyn9wKMByJQy2NJiykSiIpm3dUr3pACADXBWm5ihmMzGvHYLScutO0z2D
OLfbRKAbVPjgbwHb8pzb1CUwEURM/zeF3Tb92CeX/ysdOwZ0zN+Edi4J3+aqdrveb/j69y/fTfCi
kZID+1/RCUG4tEhwmh7GK98p+pl2PCumfV5o1xhmE+Rax3XG1gamapWWL71TrpPCq3PbuAjHycMu
dd5kzTJd1fy4qjJZEF9H75zYsIrRe4MgcguaBidvg7Ssskl5kL7j5F5KF5EHsPytUsix9HsaZ3Li
J12TfPRL38OCy3jwixKhL50oiU0F5IlCRIleq32D+sM6ooeYTZoztJEOLP1L3221jJyyI/PIMqoT
Jl8u+eUtD156i93bXNJf6Mc96b+BBswz8wnieKQapQz0co7xXWXMWSERIt6aSVQCo6vPFCRa1r8X
MZ5x1022zxLjGR5tTZZKdXQ1+6Y53vJNzmG/qSH+QOlcxxfNZYz2O1ota4UoPUp2hpFU8ZgJXb7W
ahgIFcIjBmd3M1+TqtCraLJbqU9kHEF8QF/sOzo7sIO/R2DcE0ufXdOBr6AyByaTtY5cIDhA3jAu
s6UIbzKCfdGL6Plhe/hsMIT0lXwlwAlbLFaeVem9IxaJe5x5ZycM23Gbv9zphbjSolDAvBh8337u
TlI/3Q7OAVSEYT0Z65BJpqUNwGujZknSEyPrX80O7GCn+NTVyWOqXTUzY8mad2SwDT/wb3TRjT0k
IFn19G3gzUX32vGTghuiWiJQNK8dlbbC8vx+Ep7WyNPBrvj/moYligjSYZqQQHF7f1DpjgvsfYhT
/HTTW7qgciZYU+Qhgfvrz7rTj+4qs8XqXE+y+8Cz1fzSM247J1G3PG2OXHapdRuJZQ4M2N3DtUoi
9nrOOtKyD0ndMH4pId09zuiCzxkcWGxNnrrd6d1O7ndAulfSZdx59ZdS+dUH2MnntLCO73Mv2H+f
zOF3FkbLcc4mN1l2kbwtFh0lf4ko8VAGVU+f2/euQmkTgj7U0HVoeUaoVfSlwoTpF8xidGbM54XW
XajjnOmoyCNpp/Mc4Yq02kHF5wrWdu+2mrUpRsuRkTzgmv+kN3qsk8ZMBBy7hG07utAC8W5+yKnL
ENfN9US22uz+nbCsbIeL7kqf25AZRQ3/PDzsmAOV8DMNrCNZZtInImlueHOwj44ywHlR6s6Wfl9J
mW8W+P/EFjfmyXdwJEMlXM+U7cthsrNyudYSEYDz0ZcuIgAP3y7bEPtPMAqRrE6ca8Omyq3t/hQ1
XSXoo9O5JhfJMrGixmxPeHwDKiNjOfRIs3lSnYicFZoUPYmw5Aa/ERUrS4wwLzbZGRHHbDFCez21
sRCDc2nxYoEfTEQZmmoJVMi2pyVnmIrjetcKviavWsIu0+mNcTkbAH6Lp6CO/IaSBKW4XD7CHmFP
LHgL4RyH49SI9RsxVjKu2JaaqkqKoMsbStAzD0R443TUMTMlqD5ob0jEBCiMvoIxsvYoIdXb9Gvs
KICgulxBliE4WpcFuLBm0g+YbwWQA7unc90AA7WEqV0Kgd7TwxjGNUK//UE1wADDpfZuFFnPh5ux
4sdvGpi52vWvB404G/B2C02xJj4jE9KMqeK1OrsIxAY32xvsbDWvSkmMBbuuheqJJJX+PKlMqC6K
R38QNauOg+AodiwU3+kEyclXYXGlDAEvnQBSZ/EknqHE3ryLjr3vTyOLdEsthi81WApAduEFE1d4
f59MRHJJy27s5Pd4wv2YoiIEzPCCKhF7ATKQg7wM+EWcyP/8jtfs0STG8weQa5pXVbAW6a78ZZ03
ILAaVVdqY3M/df+6maRoAFiEDKDNx/JS4aBkYLkgPRgM+wy+xE8wGfSQqqxKhvjISTH4AVuMqsh5
PWfzMiRCPpWBPsWczdgyqVkfATGn2+rPbmsesZAsOHDP7uN4L1UI9mnVGPRA/QMsMMndhiTcG3CL
4mz0L/yX/OVCUddCZL9WX431AqhhhE41DGeDx07Fizkq8zb9AVzKgN7we5bSfw8fg5ViqqAZ80Zu
U8Ewnnd6FEVzF9if8TE4XWJCf8WXce+FQS23fOLBRMR+xUjXDgtd07y63rC1tRdpvn19SkA3iuPC
iy0N/j1AtsJjQOMqpf17nSMsKfITJkBSfoe3+Nb4Dfykv3SNrq1ZtdQU1vaz4y100l17G4JLIZtV
3d9QBx56JS4bxPd6WtzDHK3q2qhet0uDeMqTzP6W8pqiM/2afcAOzX3oLqpw/GfOhO5qNI/VFKej
6JNGfZXYX498J/S/q41rTEHxzgY/p9o70J5F7WpMhetCE83qulIpYPpgPMTw526k8B26KMsfRHxT
EwNjSxS7kdpH0tXMK0D0R23sgTYxQebw4H+ivvOYvRP0EE8poKAKZS4/D7yaWoWFXrDrMGyS5De5
8L2PnAK2YRXyn+u7dSFGF0iZFzOtxXufBC4+LZCICI8X//k72XJG3WeSVpqNRs1n6TG85jp5AfTF
ikUBJTUtjvbfQPoqTTDy0remPpdA8fUNpJllB2nsJoEJ74vz+MzIsExZX9F2e5tob/VxHZKOkrzJ
U+CIFhxRcZZwnkWzMdpY+yQteivokmObf/Xt9ElCCZENRycg/liDs4XCOpcaJcT7/weiRaObUdBG
EknCZoUyBvfAQu3HWnVJFP+c5t12Bu1+p2FuAmu8fI7z1SAGoAALGiB83SGfDkTCSRTqIbh3yy3q
/qeyjWC1Vh9cRNqH2j42KC6WvI6EOlphNigsFapio1lnB6fwIHgEzplgUe4N+5BxF0IWC9A3gweu
r1vm4caMNb8GLC1cKw0T6/aShItilPqWcQLsN/508ccdHI1rBGP1aBJ6h89kgW4cdUkkwikVEWkD
69vpc85VZvuH5lFLsgzLXdpmnG1eBSK8Vo29dB3NpspG+0uWlDLwu8NldJNur5qidStL5uUpOrzF
vvWX+XsVavtsITr7IyjuyjbGt3X9Z2werVa+2c17tvn/FmO0TS4S+ShPtBrC64+FubgVRJSSL/Ml
e2QQTsyjxGCO4Al4ORXFUF4EQtvKvAFYfHu83BqvFOfrY2adHtq9+YXBPrIkDWUJIoPYlbZ7ED2j
qzfCYrfc/hqYXq3Jyqf4SIqnlxswt/NGkAJnV+6lhB6B8hPCgBCOWYeLIthVRhNzhPKz1ejO3Vzt
p4gGDDGy/She11rAO2vgc9Ay7xWitcHKd7FJQ6LtlAWU3QOuR9/2DJcjIuqNkSjNNrI7CdyLVshW
0FvARI/0ehT+Tdm3xaL2zns25RZi3pd6/kxTNsEeO5c+WML4Gt34qDLZ8L64P+Mvl+ByClxke6+D
6lXTmMHBoTinugKFuyybQMCkU6o4ogfzA9bdPZtPana09EOCd1ddZ/dFPYUncsIhbD7cWm0sdxNE
jbsW4Db/fJAkGyt2XUKd8xj1Ube+a+i+W3aZbmCCc+eBpvaRQF//6ov7kGQxJ6RSDUK+xmZqwVze
p2Mmtv322guAZPFbEBF77udpo8MdTV/S15PLW7ZKiwJYa7/VonjRjjbpuvV4v9/Oluhso2OvQGYu
ozh8/D6bl6V7HOoYwNl49dSqaopwvlb6AMH3er63eul2z4Ef5un/xX1gKXBwdXATuF+pkgZDfIFQ
Dj9T/K33CWcjvXX8lGopCUsiJgpF6h9cxyKjFlTal+tLf7cw8YvblyU0osiosJW6teNVxSj5e+Lt
EZ557gl5dxj13V5Oc/ogub4mhZ+U1XSCft3F4yyBdeO588mNtmJ7Cv4f5dhoEkh2GXDblLr9kAzR
S1LTx5Jv6t/QuWovb7DIX3cJagwkAFWWBjP57H3IfATv+oPRxJOU/8jtzzI3rfIE6p3WgaT79urD
8FU0+yxHCqx4gnFdj0ABmEJqhsKBcP/y9YQHm0a1eCFg9IO2cDdCYWaGDHS+xlaEjtMQAmfJ3l10
rNWWnVo8SeFizcDZct6WCN7eGxHjVw8TVMEltY1w1w1snIU/kLc/KRF2STopYF4dp8NX9L+nIDUT
Ug4BK7P6TM4aTYyzuLp0JTYeGQm7Nax5lP8AoG127+hUbFa78Y1Bua1jnFBjOTGfUN4feUSx8A50
dbpgtHltQsDsg09VySpUEqkBOX09npqr5PBEJ+/4Xo+IMLP2ApC/r2G9uLfXHZB+06LloHDsvuH5
cukadK1G9bggelBDdqg9OJRJwbEFnr7pKNzPPGeYdi5dwH2KqMTnibhKsDnqs9FS96i704GDPY/+
7mtloaGNT7g0yL+JgB8l1+zU3u+zhmbd0/fLWYI6Fz6Bgo0L8V+KVtBMISQ6v1oaQ0PSqXrzTw+j
MTTwyk+seoeIPWIBE2ducRJt8Gpqh7Sq57potwoOXVlOoknJ1IvfmGDtiJbelsAhtyfWy0H+Zb5U
hhBKaU7Sz0RiXCx0TB/1Qa9lWe4uqhQbU6V0ty7QgvniUCyLW53I4car4RxKAdHG54kSx/p5JmEY
qSwFCMaEpmZlv4P+t3uZ/cbnF1zQHJUXmydayopjbQLSBkL+Av4pbllvaUbadKMvybYyQkeZ5EpN
aQtpZN9adzuDgmSx0W08rD3OLntcLi6RxSRwKM+sjAJfiPIkjZa7TX4fOv3BXj8ufmWs/PAFQNBC
iulNrirCqr6LluY1EES5sfaKcEuPmbi94Llf7QtnXUUjUohBunN0ZqudWORWwKpiqEbZFOhDLZ87
gs6kD0VuhRc02aeNnumlCSji5hC+tqyqUCHWHwqKF3FovQaVOjXK79uvf7cqBf0+PeHuOW5ogYzG
NwjT0Bs4KAjcJ+rAIvHidIR0v1qZ94yScUkQUEek886Qk7CsRDBCIA+Y56ZhEQY8zumYRMryMrIh
B0tzEIGzviqt55yDAnbxf9/f8WbVo763QkH5WLiV8Fy3nzNMI4FWbFzNpC1otaWCw8A1iG/WGEjn
raJSQm7vW0PWP2pDeoykTmYbiXf3SiczTvDGM8J1GgfE63kGRuSbaFMSHgW8pZFy78H9YNDcgIJ1
gkN66b5D7dhdCSc7XyOfW32v3O02D0hJSZf/TaWPhxuOOyw4IDepXpzrZ+gGwurcUo1+SAXOyYQQ
Z/N1aMKNjt0HvO1Eq6TkCOo501HludTU2X9ybEVPIHjqN9ALR/MSiEwwvPOxiFB5RExk4PggmzEy
OXaVQjCadZxzEamW51J+lyF4ava17dXI3rrheIRvrOh6zBDrQy7SRmPd+7GxmOjridRLiJSnZtM9
lnR/lzXNuBI2C3IcNC7vinH4cq9BrZqz1+RZCciu00E6vNhvdXGRdVkVeRTZg9ewFSxX5BLne7IH
rptHqffr9/dFR6Zn0WICEFeihm6LJrYUfxyGgw5NqJVdBGEi+DWiuGZBhPNQbOzPTa2b/EWndTpr
zSuPnLpiYbIbyxGs7fy4t2Xcr7mitrWSmIMAN2+5OOKt7jFa/4qD+fxV6BtG0HobzzYoNfoywBXM
S6kiUcXW6FIckICHqwXwedjPREUh/eQqOYJUGLOIQa2fcwIeNPVZ0FPk3RMco0SvlyL++g9p6TMG
d2b+yfrDTJ6F3ZuyE7NUSpEq9cGdgxoF4S14KqbpZQ+GXGRI5SRMh4Mus6OE24P8DDb2uevCw4Dn
P/F3BQEQICCMzzsgZO1XEUBUJNA2QtoG9S+T+EMSSd+BnHyc8L0BYSkvusyTlS3jCpjC1cnZnvEg
+ooaXiOLQeB36OIu08T0nJdwiqOEPrTBcQgtuJw8tLSK7Jzte1AzBZDTq1CP0ZgjgRGafW0OXTkx
nrJGjpmSQyxZGR7B76cruvogh1xrHfSN0pHXX2jlbxdRGLKiqlh1abb3piZkNOeUPykFVh/N2OLX
pFoVxJ31dr/h6z+O0l1u6NNxrOeAkIYlwPmUlhG0ujVsmuPGMJMwAZIYyu+BhYBqgftaQC1Ti4gL
Mm9663uJHcHTdKJRRdOVYvhtTV84wHu95VufT3ZWllQu/pG8Fn4GYd4Tg3ttncwlxHRDfvHyRfK3
qqYPpDFfh6UofHCOt1LthCzVsISOulFV+BTB18QzLtFIZLyNFzLLkAhCOOvb9bM+YDglH2Oa6YKK
uwwP7Vxt0Vmne0SZsuWv2g0VTD+BmZ2hIODhok4w9X6YV9IYwawJK97xXBYDhaHtyYep4mQ/lRCl
xzE1/TzB69V9pneJ/mSBH2e/z6/e9cS0UdA0jxOAvLbNdzh8RjXBqv2fgNCdgZiIiT+uiWYZR0m/
5yb50mqwy6295Rma4RPPbjO1TTpwXjY/Qsby/FFGe/a2Oh6f8csu34LnM/Y=
`protect end_protected
