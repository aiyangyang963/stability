-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hpgbsPvrB3iO/ERfuMNADlculizKnvbxv/4KvDAjJ4ixxd/XT9LD2Qwt7EOZgC8K7Fds/d2Vzr0J
GSl6yFwq0Kh3x3kZZiPKUYDo6+5VkwJVANJdnriOvpkeHV3GigYW3No7nT2eFfAGN6ivj9LIfjrk
50LjXSAYow576y13+wlouv916gWq7QuqtZpqi+utaX81ZvnZl+SBoMPkFUHBCUrpXzZSEqmkJivo
j9HN2UMGKxKVbcwzC0P8FgV97gS57xBYafCDWd8Tw8XuHGOLSniZ1QLgYMCSdX4OD7P57EKycimM
jSlBSr/nmEq0L2t6cb5yrWrEtd02OwNTEdEeIA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114416)
`protect data_block
jb5EKujEac0mlWQypK7WRzi86oLtdPKYTctKC1frT88JEv+cRguHrpYRS3h0hNrVafBZp/CgQuS5
2zCWsk1/IFmmogaFAbLz1DZfqQUXaq4aC+6erYjfkYqgo9sAOm25kCPWewgXiW37FOCfzMtToV44
LyY/yZNWlzRZFNOfdkS4V7+nymlfgKfNyuVvJBMscU4sC/3HkfrHoR6IGcRD1w+hwncc/xAIR+UN
EYoH68I+nqLEo+HIxSbDG15z1tKOh/07lYTP0LwxEl7gAn5Y6y3dOyf542eKeArfhNQnrJ5qir8i
r5ifjUvr7EkZo9VzlAw/FSz7eemidWMr6W6wQPoWNPOppraqFCU4W2NjyxkgEF9dMJ+r9OrlHjG/
HEVol2rljSA8nWLXKmyXuFBhrj8QMKkG70Qq5C43epoNJpu9aW7DS1jzLV1R5br+g6ZSHl4KySbF
OBLMXlOUmXZcrRbYwWTP2cjkW2XDcgCqGyH1Gr0kVeVKkxM4d28oX4dF/un+mkYCpqpmcFAACL9T
XVO68uGOa5Kn/vpMaZ1XCJyL6gBXtJwwMGp09fiCtqM3bo0fxHvPBflMpEbs9cQEAifQlAQCoa+I
eX2vCsWUYQDFcXlLovAIq1HfD0Ar4kDeuA6xHRU8BH7ABAMj2geAWDKPgfYRkLQoqiVXgJx295Ww
3ZYLjQNLUVeWYUiY9c2z6oYz7tlfZfnhhzvVsuv+/fgkw2r76Uu4CS3PpdECtTr514WJfcrK3tsy
+FkYwlpKG8eVXkInTEfU4Tw9VuCIU2MfkYKsuu77uWXa+SeiRXlF+IBHeuEX7JW7QU+BZtct1+1/
XdwvnIO4hiQTqNQGT4wvu8UZQHYoi0P4Bc6lTIgZGcRs8VUHY74QIHrfUJiwRtH2V2Wv58Q+xiIo
2pdHBAckcr/cfVXM0PknTKaWABTckOluPlg1bPkiKBwM4DJ61/5FVqfJABhiYhZdxKDl/m/9aZaM
HimI35QwTP3rPK1MuI9CqIUEhu7o1N9dNxaGJsT1T4aRc6edgcDzrJJybTY4abiKSO3OiErxmLeP
/iapo/UQ+m4bbaTD7B7QOgqYLfm1QiEwwGsa11ujs7kb9BUnYObWEwFlPfxF41udXq1paObtd3L7
8ZJ4kjn3+RIRmEVz+ZXTqUzJG7jkz4SZcBoPSSfAGmkm5eBHn7k/j46ybPlTVN5nIqgXMQtZEDE8
Y2fSy1ZRtMRovNoxtaHk9aa3bfASB5ARa9bGtqTm3F7BIEmwIWrq8vfxdjFKi4RFW6QToWtJmph4
OyHqf5jzx5iODWtTq/Z0dtf1ZcmU/wh5zoXYsxG3TBYQocLYCgg9NCRMiPMHta2Y4zcg0dSurycV
Y+ARo5YqhxJYwioh6pGU59HA0YTB9Z5HcOWFTLbjvu56SyyEY4GeGVQhcKSpcXb2539YZ1UfIyTU
cLeESWuhXc7xKwBWN5b3BV+LX9LXqIapa3I3+TKdpL4WyJjm3mw7GxPN0YW9y/DakbdZ69aGY2+6
gUSiZvpinYsJUbIGScg87GzmFpOA5+YQ8IX8y9Rctc4DOBxkFsMqzgk/SBjtiS/g7vv+dcz+s1ap
TJQrtz7Kazs5FrD1mviEVaHmuN+ANTuPdwbplPXT+kSW7u0n+tPItNRQamhgqA9ELu8s1/DPaMyE
UKhBM/+2Rhp9yO0wGBid7hz+B21vpCfa6bT7r+DpdZemqiZdaPKobDap8xs0u6FBgKmVdCAhWoU7
OlmpEhoIW8X88vVRl6UItJgyvi+uWfTokfxE3LofdcQXc6VLu+/Wp7xetZZySPjIkznzOfcVJZQY
MnlwCfn+pj7u2RWZ0IpVfHIZ62uYb2Pr46Dm1qSZffXc5EdrfoWvc3j2fI0RI5IDa74CSuf7CfcM
45lNM+NY1pXkhEMxnVkJp+IVA/xfLCmCvSDGh1LwIeEcylmmc+e4dbBlnOQabRsXoOp7MmLRd3Rk
3U3kztd1TTTyOgSCJaMJgtyAfRhpSg01smOJHZZMgmH3zRUpzQ1/7PlmEO2eEN+mNd7pSU/Ml/8a
ypvjKUrty5iYlnABc/7eSbRWKO0SsOsMYqef1dyotAndeoDvr3MGWm2bop2eHnQ2G1AEWuHJkcTD
COJA2DmyAIc7igIod17S1Gt4VaCszqnbvjdhkImUm7f5wVRw2AJCWrqJenWSYR7sbPzOkm3RbMUe
b1YvNOgHqSblZNPnwagwxc8Ya0FMexAUB65lm76tiwtvaYjkcINj6WONGL5imYwe+Hx7ttEu10+z
NfmfK3SfgohDWS/CmjPJpGLLsSsBYpOTMcf3g+suTHpEuBHtLHCgd3kG2rGkhWa1HmRkopcRLGIR
6yj7ZbK21XfNoyVtoaOr/bmfr9KTg3mmf5TAd3J5bTwQzmTfsEIY87tDlIEn4XYSvHxHr8wChFxn
US8AECxMso390S2SfsXSdGLafV3M1Mkzu7V7Wv1RoLABcpJiC1gDpWj+2IRYgfYWlX7rzEF5eOcS
D43j7lVPcbWbruiXvSvRBopbqtZ1oR2o7CBaMkAUkSnxVI7bmgSkhLG692Hciq6JguavhjJ1g03Y
6oqGvX/lcecKqTT35QodACVuaG+4GXSFHCFM+KZ6DMXm6yB0lkjW1xFUpR1/q2npcn9SCa4VXmPg
k9VdrxV8Ufn1HEuBvw3ZG7b7gy+hzo44G0AZOZu/eWwqmc4JElElA6hSDzfnm+ovEYImVhBScsq3
/yK8TuQZd9jeHDHaUMMNcvQsG8YJeEdllSnzbZASv9LCj3nLfatI9c8+qg/QoxSgipphwnweZfdi
bnbTQSjQ78KUqiMuQOwb/8FtSlp/0Qdi/uxTpIWLXuUbapafPN9btx9x+iTwUOG53diSBZ+EoIr3
0yQgYZOyO2NYx1Kc8slW0Wge46e739xViFqzS9+L2O7fRzLbyLDxgUw/CMgZdmZkALbep96dsstZ
PXQAoHKy0hgApFNmIzUtPkmgKTxK1T7yewfD8ENaYFf67zWQKJXz2xwIDRD4aKgQ6425t10IHKOP
S2ujt4pBmJopEzW7K7PeBwWC5f6SnVd/g720oChONl3Q6dwCtEltZMMaKdkSfQsiwGE3+ZVMUWjP
l775/6VXhJasHwmmMzI95El7OOCHRdGvalIW9wkbXsnHaQ0YkKMv/liVKyi2RrlsEdZLKqTrjy+V
frQET1Dnpq4i5DhhNvT24WgYMJ/7vOZhslhm+HNC4xiQiT91J/0ofBmBOtRNaB0oEATHCYU7WWT3
Sli2PssGF5E3UkDEEdlOKHMQ9swXwOYawinctXi2/AxI41s8VkL4cL8tvgmvdQ06DrvYoVpYr0xT
5iB/4gO3TtzsU7JupqN1MnEE7wd0nKCxtK8Z4PF2m+TCd66oy1ddtuIWewMFSWNVPdAaomHoW/Vw
KFiCcC5J/XXzFXaw7SsH8eA3rbv+lfxqZB1awzTVU5t8e5NMdqs5syDi5CUKUUKvPwUCuKeOm/Vt
w+JAGlXiKxIdjfg05DBWzmYIS26+Z71Qk8ow9awk7PQHiungFKH/4ofctDydUj8XFiNEuWOfttX4
bVJN0J+tfXONO7B1qZUDsIx2IWF48beatciFsF6r7YVjzuI+S8uwWSu0S9lUbLQlBK0y43QdjyUq
pq4qzFsEYMXsJ+wDLM+GmvvO3VKCtX2IZagz2uXlgQSEfUlcAOU4X3KNmh+mGvWuRDVqyeolQqnK
dI4iAT6iAbLfFkhxJNaNl1iFzYjkM1d0tp2XiVVvh38ikpvGGLk4sU306Pexxh3iKGL6xFsCDWo8
5dQ1GMxvFFrReIW7DOBuagBb/t+m+HAisJ+c3eIdTVV4Y8rhSzpBPNON5DVHDkeBOxC7TkpsyUbc
JQ+Cz7CUbfoRlZfRylXZcG/S4q1c5VEKY9gOHCzZXy8XK3TvVSlM87+PmWgo6fhyKgg1CKpWJvHO
T2qHbO1kGoMeF8B5n5Blz2RETGVeGVJ+522ZGx9KyX/jVeBPO8yx5P9vYqTvZ8LLg0yynsFf5XEP
3BUi1k7qIsSAI1ZYJXBHwfl1WUrrDIiOXgHnntb+zNHHWwD3StpASLjY0W6Iua4iY4AIKCOnQpg/
VVxljf/vJKJuUdDF4FHnmCPYSoKYqIpq/m6QFwtk5E2orBdgdi81HmEd3ST/KhZaPmm/P9WeJreD
oyt6TNlczRcGDUjvdkjeIPDjR+h0vwhq/vA37BRss6HG3DMACUZLKN5XOCU144mchQsLq1ju+Ne1
0u8qY0lkwVqYxS5ohehUVga2LLKyRU9gwft/0kOCMt6IYnYISCYddWhbTlvqE3yIHZWozHMjSCC2
wAw9+oeSr3G/9lZ1HHpi0Ieyh9vodSOcR7ksV5B74x+5g+hRJDBPxqSSfngEivYSrvz0xF/6CJ2J
BXhvq4zJBqo+MiVDFCSslbn5Vkgr4huvRbEtVAqwa4PSGf0t9zniIIUgMr4xgHe8COmcjyIOfEEl
l4rTKp0gatLbImZiUYLDDuPzUga6tEDcXhQzilECznvsmcOBsr/4j846OGKr6VOvraMrRl350Ebm
e3shRnfit2EI9YHheV9ug3guwMMeHZBhZejgiLpJxxF6hzMfCkVFMyxVDeuLBy3Clz/GjKx/vWiA
nsqwzCewu2eZc/hp+byeTcUpdVbZQ/QSUDhvxHcP18mlUOTM9E57yfVL7PvpFSmLW2zUp9ixeL1h
EyzKY2wvC3A18ngfbT7As8tpsaEjdknqGb0svLHZRWrS2IGq914mSLfZKYCJ0IY1TXCnAiMiBcX/
p6e52DIN6o0FeFGcVJnCy8b9TsJjgj9dUmExjF5K6W2pVqJ60BNRWlJkkGI30S24JsYV+FrhJCiU
NW9FX9wh6CP0sIhIo84hVUTw4hyF3A1YzZXJbXxYhaCHQgAPcvQRODMMRr2ZE6/WJZiHomsyJnWg
NAQV/YgHTmO5NF6ey7fm39uewXET+H8ITTmNeXNe0AFnIcc7AZ5VzIPtvHnovR6o0FrWUCSREHUH
00Gr/iOGXYZqXaVvv3MxmgqtmrA7EaG2WqHIiW1t8De28zmOF6nBG6uRh1Y13NBGbVkU+N2qLcvF
lid2870OsEBjhmET9Pog4a70GSHfkz7f6k63f1mIBBEgzh03B0yBvzXFSN4joPRgnfLT2M6uMd3o
LGGESOG7vMcUvov2gb8JCWeHNgrIuyCPc70nURn+4Ncpl2gK3WLCkx6vnkaq48nI10omiRTlSu4K
D+p9v9RmxRZd812g5pb/jQilOW0oRO+MYp16982M/vYcO/rXeiF/KQHG9cokrSz/ehSatrQhO6Ym
bhHiLdRpH9DuglIzbEzwEMbKxD6Lo3b2469hLr0dpn+DDMubhI29Jn9Z773qH6g/ye5tUipzyZKt
ftPN3477C0/IIrLmMUq8XeXjGhn2Q7NvKGP7OcWIoMfvOH3fZqokWB0vK3iq9GbmOLehIR5x4Mj1
cX2xaNbz3R+osBdHV0WMgbu1IaKW1n7df1VH+Skh1jlGrybrO648mUoacnFKcR0Les2HEyTyBivT
hkT3rH77P+qPBV+HtAMtDCNAVclLF58iYkEWgSwL82G8XWvkem3CK/cA+dxhs42/pOpEK2FDnzCB
niVFGoBwIi0yF+xkDGfeWyVp1oMBUV484VAww4L2TRsfJNBRDOXP7KhwoANGbdNtwqOYFMTDn2g7
uUnFLaDO3y2L3rRAzLCXZubSy+8JBK6ytX2RkPtXtoOb4BhPGBNJZWS4uIH0Jkx8cpx62LY/t3HD
8oBTjwEYrixL4mAeU8DQca4gnveDvhYY3tLpCh1BrHl50VTkwTO5M6F9hQFpS+iFtjXfLOVm9LMc
Ar8OTLMQfop5cf+FTy3XFArzTmeRHr6cChEiRnKOPAITBC8Ax1yyAp8GqWRHt/1/imd68fHY+auC
2PzSOj2ONdOnW/xc6TuyymFOqsFbzhCsxdLFJYp4GfEl6grfxFH7uarMoitl6SExl43kkSFn/L6X
2f/wdh3/cfYJt6nBhsFy7AY1pYMReD1AUEZzDkANNO6AIK5bkitnpcKG46qwknHJUae0R52l85+N
WEi9vgbsUF6236fzSBD2oXNItYgedU1ZMpmhrBKJ6neh6twKoxaKVssuhQqKZEmVpTVt6w3/L+aq
3Wj8PhZsOVMfD2YReNVdO+gxn1VIvmniwX3aLjcI6HuXu+l0racAPgTRJ0ZoL0S2ynuQApRgGAB8
wRpHoQ8KaQvKG3XtFphaeV+McecKeOwtjzFLqjIxfEtCm/HGkbY2ZnnVBZFxT6eCmgrsWhV8usxB
TEvQ4q7rZiQwcyHRFGiZOXvVvaJf9uQKAOh35TWZsBiqQU4h0aigqUcGt2eQjjiOPHINnACAjQY6
tk2rG+PyYdQRXXOcWch5WXDaY6dNoA3N6BcS5TpG5/wC7/MkL5iSMGQMFNMexQZjRWSR6U3Nc828
ZCMIczJTdQdHGael4qrizekyPFSDUXirq+Swn4QUc3bAQYC7yUT/ThRbarAZOmWdIvyWIzFaK5b6
vrU5RbNngQXjVyB1Q3qaHrJKPkFxZHo5SNd4j1jxne2/qBkK6+KyPpdb6y48WAfTnRdPDumxONTb
pj5m/PVdzmPoP4+4eA8sBdZbzzFeImTvckeSr/rniL3qlzYd+UTowPDNAubl3U8rE8X+t+7KOhsg
hYIjz/ZiBsC+/T3rlUXnIrW0FaOS8BiZ+24PCSnSjR8evawV0UZk6MVOiZl8Hj2WlA05XzT77Ax2
X0YuqlvejC84VXuyMVcim2asCdkten7kY/08Zz7gnsUR8WynnsKZ++h8hLIaxHdPFy10YDx3ohnQ
u5Olh4rNpCWz05mkT+Mqt4glagZ2L0CuhtjVi0nBRcpWZEOnOVY/wnhTceM7VHYIgMM2Mu8nYG/a
Fyqxvtm6XKfGEQhMNemAh4V0r1kdXXa/k6p7xN7lOvmRsQufSnhzW5UohhqS4KPpFLtz6lAD1ZvH
nNsVMpq0u4vaKExtsv+yFDZhRF5MAw0IZod0/aQvcJ2d8bdZjoN/1cFykcFswBQvtuxokK7c+7f2
uJqQSRK/jOgv5fe+1U8d5XG9PBzIVTG8VGcuy4RHdm7T6Uh3Khu4UtCPGzhF8xAFDZ1XyNsspJBb
DwtolBroEw8NwvkkXRaMhzz4r60096qL8+R569i/hugMakGpspPZsj4QG1tew9KQOE/jwS+f7t0X
NBcowCix2nhKyqpaerAl/LWgbJQYVhIJj5iTSMx1pMR8Tds8HZU5eoEplCxsUmAMA8tTv/dy4c78
7qfHMqKuV3GFbSAojzeUOUkPPy7dFKM66VftKWSPAv4twP2IgdyM6Re2bjJ+kHibJiU9WP4+pK0B
sgRs2RL3eYqRQXKGQav/ZEH+av8FDJwUT5kOUSE2rkl2P0gB1L81GsKAvY35Odtz9C3yqMWqazTo
rikHLzIm+oDRIvJeroo7YJNR9OCTArU2E0tlGfuiak9ok0V+MBj943sUsankhCt1xv0LEnDDcEKO
0xm/jae1elLCxnz8Y/XYiTpQFmM+mcdMn8AsNRmc5d53kRMg0f/YDf8ycAaMC6WH3zKiXluyy4AF
6vNvKHg091UjVH2NBGbmeUZkEMUrqO8fmct/bn8MHRWd71PI64vDgrEsAMqYhLfZ9i5S/zz0PkZ4
juSZfYLOg2vPfon2rysu8CNSdzBCoPTcwDQ93Au1ArGRg2w189CzyKgi48x9S42aJ4HO5MNczHcc
60WQN5k8YyKRTxpHhMkMflu94adMQdLuqOK6KqGo8K/xReqxHO58uxm9RcWHgLZ+cHj5PGf74VT5
lVqjsM5/PmqzdrkqwF3zphQx07fTpdhgF/YBz2gJ2WPQFczGxsLkwmLj94Gj2Z4OibCSQl1zjgNl
6vnpAfz7FNeejq8v/5oMPSuyeXbcTVl8Ttj7yMIsRnpQHLlYdu7eE25fglJQ3RApMHhyBnDSFZUh
Lz0nIwjWqBXzTDFyOKOLBo0QX4VViegM/Mg6zg6+B7/7wFPHC2TYzOH+Y2Yk+8totNRYQwqLZ6JR
UhLdO42OQ18tFzKWwFb36hz2cTWEoAdEOtWTubeO77Qd5LuEq7f5ISitF9q4QfjbPiwe46Z4up4I
FyqYwDmjyCABgpYzM7jhSRVN/DGkEp+nPAlz0uL2nq9/RTOOiEcsHOJRDlOaVFhwB+6GImtq3n9s
II7p9OSD0Gj/0DrZm4KUCXInU5R5Au9mSDeYmhAMBoOi3wlXB7gXlEdaAJEYYrmRkXSGrAJYB9yI
RXrx8571FilXHa0Z0vpZzpkU4Q4ntF42l2AO4/ooyd0xIm0hZhUuzfV4+VwN/GGTY+svn6OI5yO4
39CMzE00AB5v03AvPpZlGTx2zzEKM9lUknNV2Xw28etPtS6S8zTIHIX7UzDKl+pZ70Mugo5mFlEX
6XF/4vKtm0SeXt/mcgTaHajIBEfEt5Y9kwg6W6XLucW4izSe7eMvImDKZc7+arZSonJDM4tPq65V
JQ2lgPCZGU5vikkdw4v8AsRwSGTqOJymvv89kElNtYS0FoS2jjQ+8LDPvyznuHupXBoAvwbi10Wo
EhTOe1M5lZzxj2urkPAMfH/iuEkZa6R8E74Kd4B7d6OE5hqJ+6cfY5Xv/f5iFx3hRoFUX5Cj1Kro
4Sy+3JJJsJ+SnTbNacBrj+GX2hBKcjADLKi3hWpCA6G7lUNIb0/oBcQsd/M9tmlsg9AUDzV17WxY
F9AvDI3aZJgLHljZ9FSTXeO6jZuVthY7li+R5D86NbJ/5vyjgoPxssc7BgjLtST5UxF8Xvk9VKDy
MiLG4/s9wAsbelk5NT+Yn1qtZDTIZ5NzFGzA/g6slxfwX8JJSPKYs+IgtUrnxylg2pr+eAb7Hhmc
xbj4Eeij0emxT8tO71xH7xFsxpktFWcnScP4UKQ97T2AtnV/5aJPknLyXCySFfoWyDawAobJOQFh
zoPCYlKDb+3K++q07Boy+LHwgC7tTh5IAi0s8NGrekp/9Prj48h/vtFgOJJthJ0UWeGQttoQNLR9
CI0Whmh1MKnfrDMsDcareGlrQcCaFYnRgQryMnuPz4HZcaeKQU3bCH0pxRQkttuhb5WfC2YVomFB
Bx6Cit+40UaFUcKjKhPgVl/2uUJMjuWrLu6/QdSjbzDrFy/wZyq71GFnDJr0Z6vnSNgZXmL9m1ut
HGH2M8p/19yFe4Preepl+vb6GoWFZcY1p51vhwIYtAC61ZTzPPpCdWyLdODrtK30y1aWXJaFvXdd
V7T+aOHT3uYxIvzChCk6QM4KlYCDW7/tpfave1A+Lbn3ZCaBlCqmOyh8YwrzpNqE7PFkhe7ZwNW8
niEqik6DgxAqiPB5LVh/KKXLFBAYKUc8/0RAOao3t3FQVx2bExX89s0bk7msWg31PRe1Uw4/Fi+E
T9r1hWWTBjP44RtYLVW1hqUpDzvjqUZZNjrK07nALQnTKhOsTgOPvahEtLfYYWL/AaT76IlVpNoU
3MxZIvsiW8ACjAoOIKbBVUhCH8irkEuaiUqiInrx9ZbsZoFfL6I1iYLIfvGXZ2tCjxtimq5ccqV6
czPvv3/qE4yiFMPohk+mgKNmIui4hdemaX6xewZsKpDbss9ZxLmOAwgKLQ9f8CqEKRaMm43virAD
TXgslUMMmu7Lzn9OpxnmbbSUvrbJ0Nwz1gKJbbvrtle/w54Nxn8uqNPcGLDQ3/j+mbu0wU83Sj+1
zPXXhhjpV4ItKtsSW0ta4YfhfRYcuupzqZRa/g7J8Ufz7J5jR6x2je6375iEqt7gih27PLyxoI9F
CK6bKWOTiSPzRjIOBz3A9VudSUpr3KiPBh+Lbtv54nx/7c8F2hFIVAlm9UgK6S5VDyt+bHF4aKo8
kzKSUtzV2G9z+TIDUWsO+d2E262q6GS66vnuJ5Wc3FpzS6Bt8Ca2HG0E6sATcE0VY14VFmKK1xyQ
dryhiuuVslqJwRK616UnDIqopZyYGBMI/uFwb4LL/UH3TCYk9OxVYozCZlzraSzorgf57XxYg/jL
OIANKWHCOWBm/SaA2ULHmXQAK/CX2xIyRhiR95PpkJyv0gLqUKRMaSkALADLuhaEKIGgD7J5mZFF
xy0EoSFd0v8ym88kMgjC/K67YbhJPWbB7zFggG3Z3/Y1AJABiiNexN2EyIEkLbiOuciuLFoWxy0i
qaLuLfODPKkfsSkCQbM1ztxSMYD4VxUGQuBJUndSPIIq25EbO2M6FXH3P1/XTiFzeC5/YYiDJesm
JyDOB2CFYcXprT5dHNJuF4cxWe8ZIwCXQnTE9MJ9dUQ0am8nP6dgLr1ygX5n3sa+dWBVw8e1o6UY
4JyWZelWbv52b1uCSAyQlzP0qRh6vmSnhRQfL0LcJtxrMaOGoxbmXUTnpKqVfDqiIIQn1BSj8cby
OuCOs7L/ejzEJFc+j+v2VU1ztXrwXpzhG6wqLoYqYnBGtwberpJh6hcjUKzSSjIGRMcwg8M4lYFs
h6zDxS588S6LlMKnI6lfv4GmzC0Y/5Ym8DvnsyrZtkBnCNFhY46YatByeja4c3klaefHLyo4UMNj
3mIiT9J6VZGAgh+Gaend8ibWmsLaU+oFo4c6/8aszM+S3F8I2812ZJhHFfShsRQYgmH0pNrx6C75
ksCcF82q9SENfoywovoVJ+9GDRo6nn93pOd8KgcXP6rEVF0ndz9bg1lk5dfAm0aiKdpTl/sXHAUd
0s2UB4fosUGK6TrdcfCXyukKJJi5G8BgtFFRXkfRYrpVpTd6WjvS5OTJOw2u5H64nD5zMhb4rBNp
vrLJTYmNBGn8uYAJ61b5xxKVwPS5CWd+lGAf062SUBOQa7wXxXJVJH3aA/I5LrGsUrNj2ZGievNd
A8IOrI3Fls1Ik5aSyFSP4uDQoms01+20YQFe4jdUHWz0gl0N8YaXNGXFSG0q6p78i40oi+FXCaLj
QOr9vd9VZ6CW8w0lkYVmtWhcC3Ri3ZYj+cmsFLeiq74DaZ8RuGNYE0y8EH/nAD+FMC+OzzVbAc2q
ZL6CM0jPlpsurpDtJMVbhe1vK/jn5PvoDgkyVdS/3lgEuqyK6dBYwzLjbenboefp1IdGP3FCSmEu
SsSJb8A5oNFsh1Jp5xJoNSeKhYUBZqS/AUacmxdVxC9dGPeBZU/lrnMOurY232hWz3/8JrTx7Oxm
8yw93qV81gxGiNgs58MSbY/TAlYJsH0JgNQrczPBPkpy+25Z6rV/GP9ofP/nXHkUNUB9EQ6z/prv
zYzfppPlV36Wu7JnohF63zIptSLuKlmxj8mSFthzQh0ptjRnFd6iRhu9RaQqCtKqZcpYdlxsHPxg
Nse8aAQymkGQx8U1e1hlhDHSq5EYBi+rakZMSTQW4P3zoKK1N4zv6/BFtTuFuTt2G6qgoRQFDxTK
cXXibCETfGes6O0tmxKH5LlbU8AVrmnFqX47ClDuT60wdrCGYGXDdoq8Y9fU3iVzxBGFWl189+Ia
HYRkz4QeysuWYll60Y9Vyz7o3F9H8sRJXNlg485xrCMSeF1nCfqUxlMppggXgZ4xUiXZQ/vn3k1S
QDUP1PT0xk+fT55qCkVhRYtlBmGMURHSo4UqQOkHXN11pnyCUC7VhbGiTq4KwI2hB2fVvnPf9ptB
ARuVCyyqay/LbknyR0xkUDcAn78/mqscMCz8JzR+o3m/pd84EmcPtXsBqEMzk0BQAdFohdw80qaa
4yavjoFahGGGOZo2KzYno62B1WcBf/5qvtpzzxbbt7g9P/WV5BJfrPu11St34FP5V51XX3GJmnAH
ucMx29nGq/noBIGn0yDS4EQ+J2lmPn8QCTMWsZIjgcEw7p0uhycnTbu3J17tLr+d+pHH0qFZAovt
TfwGM3r7ix/8PsPJW18rC2sUiRLhB+vSfsGUkTDcZybcr7TT6CjdeaVkzXDrgwuy6gp6fV82rZVx
gVyEDBsfGr5nQ4875P4G05CxSsIg3cO6LI4KeewKW1TqOz/IaoKSx/P0lY1QOYyW63ktIy7dNgVh
/QgnjiIQgdJ1Lvyo1abMJHeql6cgi+q4y6Cl7IpmeUx/6vATWUhBuiRBnxDSxAg8lsqxUinD9q49
cVhivxj1B/14zOY2mPKsJps+IOPdsLemiau75ujouJwnq1l1nh7BQ9EbTo1Ut2wOhLNTmWah0RMb
kTuAt1ORo4IMlbbnjtA6lpRVa83FuxsOxNhXPMqadFCe5m9nwL2RNvA1E4O6dyp3DAktXkWCUujQ
+kaPT8FxZ0P2k6gNWLgLh2B3Zg+gjtph0yGAKH0z/6wiqqBPqQDJ7XiSsbT058yNj7/Thm2SOw0b
Ei/aJrbhNIKIzqP2pf0wxSBGbLZ0YyI54cgCSvk4CffexbTnxRPVzSPJ3SZoh+Bkb1SR2NBEUUSh
IIQp9a6S9pNbfNOvzdC6FSXuOIOMQFNz8tltPiSYKmz+RZKuNrWy37/A3O7yGX4lzUxo8yd4o/zu
0YKkhlrN0bCXQ7b+luBvHClZy/U/9MV3qBr9NXvSMtp9S4LwJEAlXTm75KtloCmvycC/dZ/AgdI/
Y8/LkV1bygAUTp039nM6WSXBm/r0XMRaBU2IlwD5LjRnmAEJ2M7rvmCpzPfISxGw6sSsP+EI17Gh
HzXdDCzqhgbseeEfQWJeW/Wb2ab2k3LrqHwFb5R9TOpMiBfrY8RNlDM/u/Ih48HYCOydqwo1gm+l
57iRxRLcSQOlTV6MhDBzWd++H2Q4R3D0bA7t2sWltJTRsysBTmLQVYbdI+GAyRchy7RdawKLKOJx
EvNok0Sl0OdaMdD8ZLnNw5KlIXWVmQmQvft/bj3k4xIJLbOoG3Y4a7ARzxSVBmiu7QeBDZsco9iy
qkW5WgzsZArBEokmQi/V0+6AHyf2emJASsGKPZ3Y/C3zOjdG3Utu2/nYN3JdehUYEXFQtHW9rAcW
XePtWxhZeGiiJinUkWnZyeVORY3OxrsoZ+Kf0qft/E8ix9dwia4ztYt0EWDBgbQE/DW/RLOmOBeO
JIpT3ZleWFhFY6bA7UhRuhcKX4SpTR18XivMd2tPoVrgLOCatuygZUjGlWP+Y65Yv8HkBXopKWHq
mR3E0zFxn9W0pLOlJAopw+ASXvTUKoNu5moQelNIX13mGY+4L9MWMfFE8mMvRF1fZv3MNHyKr6m+
5TPXMDXAhJuQEUYS3it+FkSAcFaLKQtAcyk3tYFf7Ige+tMGsxV1/QhPzUKvWdCKfHAENTho9bek
Ea1x13BqvUuc5dp0n9ScXy3Qj+ghxoMaHlypkQaVZHfNo7LmVv+by2odjEp2UhH1MBi0T3luatJ1
gXbEoG7Ci+wjCyI5PrGEtX05VLBofcLI/zcpVf4puZyVkNpOjgHvXNY/MyLHN4+piqZrpM3wac59
txFjcDJGJ9kUXULsFTIgIn/c8LqQwq9R+J2sDwwjNNY8Qdhp6bsuOZQjD2+PSBuBMMoxwb2LQazz
WO+amPQ0khNkJr2YQbzt7wuTD4KsL6+LUwN92GN2z3vOT2N6tXwHQX5jrK045mcvLkeNb/XnCOqB
g5pxBzejVbv+GAdmYIQzbl5p7vo896F8hiTHtCYgVwo5kbaX8s7zjHrfLD/DMX7GymvRJytwSkoo
FJa7E5RhMH9YP5hOUvBhc1/gJQHFkmNy0aRth/C+U6nzENpeUjAiSjmpsFUcwPMjqrI078lrfFo2
cCe3XZfrXDgI8Q42uGe6t6nmuwgngC4kYs38kKV0qNcdVQOEpy9PDKhUvGQBkb4JRy7DSTnARplJ
OcY9/8rvmjs/VAE1N2MAccJFyShNMVnUJ2fqzuSa65yIa+yBdeMOiO2b470aeGI+Z+EOVa5S61UY
t2UN0iIlbbzX51yUrr1vwqhTBqqXdtGnKr7moGnXEbXYJCaMG8DwrZjym7qXYU9RT9t9BnW4Nqg/
4AHFULIBsNumpon6pCxfaguT1J6AAaSOegogjWs52yaPpZSj0t79Rj+Ol6FG9HfRftL4YzzMHWUP
vze0RGPKtd8zuXEUCqXiGO4Vs4+d+p+QcZhxi7cLm3ZmeSF/Rm3+oLC8z0GHcYU9z1rdJVcbzTMu
xQNis2yXp/Bqdj/8vlv1yqbbDzj5IIm7nYj2n+AMu268s57UJmJkgxyFE/6MuzAoz/IQ52cwgXc0
zCTWtEfVdLfd1DRZHRibll5MVTHZEZ6DrPacpB5t1OujOej1VtygPKWk1GUpfp/P9XCDGL6oFAq7
8LOAQs3sfDipqeTNghKdBN4U24J9W+jNfPvQZh+qkSk6yyLyC+wT4J+i8oCUdRZ/GPRmw9399d7m
bxsyNIJLZxw94YN6IMQQWO8/EsK5oiODKm0fV4J2BN+CLOjXpM/CcCI+tz5UUXqW37A4qzWoZA+W
nR7lw0Qws74UiwKjuXkavCB2WMIitdLnkGnrLz1w4aLZXXayfq+gtCdKh8ERadFY/jttLxr19kML
aNMczCqKIEsA58wB4As1KysPdmPrirzuB1VgThSVg+EAWBy9m4zJ7v0gz+XjMB936u+1B3pIeGDC
osbTRukNNBKBIp7XhCTCqz8bygUU9YF9Q+ZMV1+2cVjFQS7SE6W28IT7SpfwBzoomoEmcv5T6NEq
hNx0Yqrbt7Hzd1ddBn4GTWN5DKvtHQMxoE8M+Ow7YmG3QaV+xSdl4OKF45ApnRijEGl3bhnLHurL
cIKYqFCMkn70aqfLUPYnx6V+2K3SUu5OTbZPs6xSF2TcihiF/yI2lt0VQOl8EaWaaLLnU1wGpVhK
Mw0OTqQWT5fO0kcrrLdGLyitm/h9wBDfmtYzkFaKh+frdIhJWL6PRHR990K7OXpaby7/7/SGrlx/
efoWMuzyf+riSLmf5yEaTGBZ0zWatr6cCrHmXQQCVVch5t4Gm5iPeSaAC+wiFo2fCW4L1hPxZdXR
Bqrg4NlsYdfzGGZHlQoZNxLGI1NjffwiJnIAqxBdokUkQtzvxN6VNrrd7pyVAIXxAcJf7EBWtWrd
pP13pvpVtYxYJZhMuHXQseYHLhcNxxfqfI12kPUXzSWQ+f153FBfn8LZKlmJWO2Ikg4DwhR1dOop
7T5hiAMyPFnfJn/djGprKpH+3XsYGxKKVeXTcoFlJBuxvpBZanmN6LrqejvxkLPfl3VUtF89ys0T
ULN2PmYvdGTV8pah6M+9xRu6hgjHi4SjTP9mOZuZFpWAlHUQJixvvslva+wn1GzWBKugl4kipJeP
38q/V7LdGUhKAYJshqzoF9RXLBtl+j9OWffuqu1XJ/6KAypZgj8D0nUEsqa0F0oY36Zpptpu7vAW
lzxXRBHpg1WT9nXry7hNIM/Ej7fhB2iVIzDHYkOHgaVBfHgpR+N03S3BsxEM6uRxu5Qcf8/NZnw5
vsGMVj/Dk+M9c7GleGtfJsNLcnwGGK29jQbrHk3fKZNvplJwqwB9rBH4MT/gxwGo5a7eDUw1VvGo
trIgjz3KNhH88slDgwNSxKmykS/j42tniubvWUyevI2EjYhYHh6sRkNyqzva0YHJesE4p1C+p7x5
qp6jCSljtLAOXU6pfx53aQj5ljFPRcwlrQgLMM1AaueUKd2B6mF/cLha2o8eCRNYg3SoWVlSQ7Pp
upFoUwF33fqO74wTuvdPwNrZpxrWJ3dlI/5wR0ijKey9OUkulScA+ZiE0uLrsEOf/e3QD1Ly3lE9
jdi3YGGeOMZC5igcSV5i8+2NSAPbLsz9gJjjbC24XZ6482euVlnwh/2rqgpJ7H+64f6OtcCAUGM7
kgkP72krViM8xA7VVln6nwa+IRevW1HDJResyYh7wmf1ZNehVeWjJ9vGCYoRjnECc3iZlgQgISZB
f+a4++s8MLJQ9ZTyKF8z6VXTYDGAc3ea0RIZEbvU6RVsWlltlfApQAJ5d3M6pWob3CBczvajxdoj
cozC+2BkWovbEwBnIrfhjZ/McMbRorWqEuN5fzpNnHWBQicuWaw0QajfnNnYsYEf+02Us7Ok4kDk
mxT7diMi70CbMw7MEN76CICrSS0asvgBA1A6bdh4yHyZAljaqJI+8RYqz2CdnKMoKxJliV5uZ0M3
lbojEdri1l5ief7NzJ7n3hpY6kLyQfU20Xa1b8FhBfDVRsagTkCB0uPKpUpBFJSWoYScBKW5it0x
/2buyLkApyg/cXN1bPL/0KVRz0HQMSCCZYH2bjoDXktAOVpBPMyxH0/+JqI7lom98UAnbZcNfnNu
8nYdZ7QVsOrcHP2upVULn6dCNaCq4Z6BNhfNlsxy56hBDW/KDhdgnEZhJW9ULES+h1CRntVYifIJ
Jo8NZCXKeBiwLpS5LybS6LNOPlzo640pMaTbVaPE7A1wwHdN+9HvCgzt2ZcwTzyBKLNRFeX2JpaV
PaiJ4ZpxOtXYOo1tqqvJpj4kX/ZT1YIOQhnQmwHCcTNU/6d72IsJ4d6Y8+3aGpjvyspd7ygXpvyA
xC7DH3C989ntC2l1ip8w4H1sf36/wHADzKAtJxDvlWUEhwyD0xLxoHbbLGgDM8CBg3J9TIje0r/e
BhGiVA7kdPM5L3SlBjxJxKAdsZ/vjyvaBcXpe8Hc551mV4WWC24BUBrMMGjk2i0BNjRM3NRY9WUe
gwKLEp3uikKH8o8K/pQ3PVIrcJZT/cpVkEY1QJTsdRSXcOMjNdZOTHdSOsYHW77NCXDZlE4UwzjX
zhv7i233m2HrvS2NDQDCE616NdnToxHk/U8qdYm7VbY+T570jvwxt+ENK0af5pZa72T7F9DsMyY6
XkICQk10Q9pQnnkOLDXV5VweSsvq6DhqhMw4nVkpQQFyi0yc3z12/n1pCMNufor5oe8fOx9e73gZ
nOzPud3eDYgOnPsgA/ZMQKBAS5GZiANwRtFb+zixe4cfYseC4JT6jKMX329wXCS3//HKbrq7ld8F
M6lQtAXL9OcGRyGAwCtdJJrWOD5KbMI8mgO3md2xNkJpOjZjP+/Z/9Pcqxk8BD02yUygdVqLmt9R
0cuM41l8Y5o4iVZ8gUSWQh7o3PjeTDUhK2Dly3xHJf1FaIWQMwOUDy+1jMG1NmKO0h1D9RDDGxwV
oRz61t5aZWwT3thrh1ArP/RlQ6xUfYap4RLJiP8D0UgH51Af79DxuD4uTPVS+lpWYwmGHw3S3MZG
sM2mpVmTi96T7RpWrxYv6ZMX9dh9kpRN1XJywuXda3eAHkbIpkKEJokhhuKWUScQZbjgNyX8Dljq
y0YEt5ndtxEiN38Lom88d4TWdEs8fzVVNUcW26o9Beii/mqMAWrmMv7dQxwCvuQVZ3Bk49iuSD8F
wa3Km/pgU2RWwj8VeIq6uZf5tCiONuphnFOn7eKg3PLyhT1X0wYeXxC11Q5IIL174BG2AguPjGKb
HH4umHCpCzAb/oOKEef6GPzz8guYjwvQYQu4vNtGMrKzALejtdhNDAcbw6RDbv5o1jrukDKQ16UB
giDyzvuzxCcE1FQg9iiBYe9uGkUy3S3T95/BQWr+OjE3b4kDONSINsRoLwrVAeozbxePN7XyEaGg
ZLHvJORsZBcWy4DwTlmVuckENWArLYixCx8nvMPV/rXD6a0VyLgEjSIXLfy+4x31VP5JLvl8EQsa
k4rsTO0IWFEX0grBKichzN4X2Sp5q9RKbmI/Do/Ni1q/2Ic4lJGTKrYHnDhY+o0PDf0mPf4w4mYK
UZJ6o2jAEaZe6fHhpnruI+MyDU9V3FiuHAOC14zQznkjuJxzbJihM55Ph1p+KkIkOuJkmf5QxAyl
+fcQ7hbMvJIsZ2opvyDicJpf2AGbSlqZTuO2XM1zegfG74N9LZOd6H9xSoXahDDi2d9iYY1aXtqW
AM/gS460Nc4OZ+YlFeTXTHd2bVdgS1Gek19bcfxyqEbgr7ofelml9goGzmgPDJQmSvoGUIyGKI+z
/rJeXkFj4JVcNJG3qMDpGUtRgyQ33CwgX8xwzmQcwb9SCvIZzkVLGSXkpgFzwNWVEW5I2obJg8na
9s6tgLuVXeC4wBdHIkm+TabVdxpaecXvjLaUJNh+sPrD/OvKiCPDw2YXTkFDFtflGPgkr+39ndNR
NQp+G7LPglTOeVwHrfDyaey/ukqngUMVjWM9yZXUKrcQFnqW6tRO3xq4bbzWtWkdCJTq4JIUQzJM
3st4/qC0MUeu1OPfo9ZiRSLq16d9s2MIQRCsQlQGqb454oyrw+RRhMNvdqIqPNHY0EEWa2HIQopC
AcO1y5jfl9820Fbdh1RsdKo4mly49Tsi0HauDKV93oWG4ELEUNyyq/tPRymlZHZGx7jpJwkR7/SY
e6HdTTdGwUBe3oHZzJRx2VpIuQE6ledsW3TV+EJiPUFiVkcY9Y9UkKSqdbxiIyfy3LONwrLEbE0s
2MlyTuTs3akb+8prIsyTJ2eHiUwEMOeqKOcFvWXQc37eRUBkYhZK0O5+HntQ8XDLWZdv/AqoyvaB
Im3e95n8OEeVSnkicdb3/xTUHneQg4ilN03K4DGgqm7oAVsWcDpx8Cc3XK3LFqBzRtgP6M2RPfsN
CJAWqLMvkHuszAd03ilKGhWZkc0zQmuSZMj40Vhrg/xBkh3VEt+Bi6yJHP3AIiTyiCRO0ItNNp4O
O80UOWXloR2LOYfhKr8IPwSsEhsIxBzDz5PnbWGBQVlLYMtUGJGJt07zgrpnbGTrXhtskLpYyuKT
BqeEgrRXLec7Y8lC4YqSg+6FoahhtISav8gmpZbE8Cc32mbIgnRza62cv4FDXVSucJH11yJ5p5RG
PxJsBs7t4pftfhffQV1AKjpN/K8DGBlEXwpQhsQHy3lGpVmS5aeAsECFPyDUW2om7Knks1B1xYkK
SKJa60BOXeRSVXhVuebb+z/eMc6uEIUtCkJ2/H7xWJBmqyX03A6dc5K9wYPI2CeMJDfi0bLdOeQp
/cqNqxWer6zANtCsc8IYa9yzPa7saploNp5er7Rq/CogcRqxQ6G3c2Q1HrQh1/RhwjTOEaBtddH1
CZqLa0oMrcDssqEQwcEFWGgedO14Xiyk4J4uItQdEAN4Q9054J+8kzqxctxrNAP9AIKDwNs+8MQJ
R2WI6Or+lD4PYygAWHAvbHu2DW5fYCGm1oZMqz2U1yY8e29JWCHKiaBKGm035Q2K8ldE606QbglF
hBy6Xsz3iCOJsbEnD8sTIQ5tw65Oaj78Kvk6sPVuGPvu0SDOgB4rE7P7s6ixIoHa2k5hcGuNq6hr
+Z18zWwIlkUjrcrx5f8ne8Q/BOEVtiZKUp00X5p8rYufQK6IsYDJC9yFBLofmaNFn2RQ1OjRYBBn
tG6BpcrfHycSeGeJwzxAPlPUN5lEXP69vSpFRl9X7+VOGcfYbzIK51eT4rSu956zvwT6Ng+m2xpy
Acc5yVy5tjlRgeKGKjHEDZQVH21WT4+EfgpYvZsV6Q95MVGK6my5sQaAG68bhm8sytqfO14OeqgQ
fkyrvTV39Fjhje2B0GCF5dVAldWCKd2elJC9XSFYr2y/kJsrRaGmSIhawr5X10yHvIcT5T8+rnns
kP/JvgPYbG8AfLjYs1Is1K0pQUbohWPEw8ZWDk15BkyyveioryA+2C70ZSsls9GUQyOVSLgp/zvq
fjvjM22QUNPPPYPQel3bGlmDSjUPYb1xpvasWODsTkOq1uPQ/yVpI+GNupkRBtvEn3KrF+vRxhoM
VeWx90BojIzcYai7HuTBWQF3pfeMFOYLka2kRyR5kwnr1LEh20dYpwrAedJ0MWAiY+Aw3IpSlPro
rqI3EcXnIBRCMVIxV57jXi5X0GDiTcFu+JExUyjYY9/xjMd3DpxRlMy5ArKKNMrgFUbtlshO/Yv+
vVCgLIi6CUFo4QpQRJnHMi5npTTmTjLvW5+poHqbSp3MR1kcBjjB3Rg6nNkmLXVqAhi2T6bbeJYR
k0VZ01/+7Gt6H9ZnlB++VGsuQo1QA2TV2IGgYawginIQpW8HOcnGVheoksKFrMQHfiOuq+7DdMh3
jrLrNOk1AkbxUJoCSOWjcBGzRFsoWBNmk9/EzsJzQQBTkouHIzs043YNN9p9U+4Auxs49TDyjDF0
6Hmo0b7udazyPx4C2HASOuMbannDkaTTlqwWgwyGMXmqbx1D5sUdTOnFeJZzr2S6J63jwwU8rYd3
YRT9A/fHX3lr1V8IVZCZV9NsoUwA3xmfVle5KPfMvdr0ZJ+WLKT4MVRt3VVdJT0lDZrUnB8UNOxE
9LJCZSgGnldv6kSvliq3Ai9JT7EzTy+HCS8F7DmGJG6xSZXZlXwQFUF2VF1D1z36A5AXl5MshY3T
UBdUn07/BaF90WHSyHwOSudpr09arjsV4FYaN2mbDSZW0tyxjsViwelvs9vO/Cu+bSRwWC3n6PNa
tgiLpsDfHmU05fp9PIDdWsXOBC2gt9Z2OEJhhmXArmxS687juJFppYX9idAJeLG8g4cmWSJoAbYs
mjpx6qFVxsNEnmGdcKX8RWxK/rerY62LNXSf3lXhY9ektIubjpv97QD6V17T+U3aXBnIXAOAASQM
DvK9y4Fqtra84L6+OaeiqA8qxM43oiftYOUdefrEwAh0ggSo6QaXlZaEl3RGSZwmfOJiwxGdIDq9
olFucKI73JMIir5vdR5LJ1vqWo2iQ7QbtnRWj8FIIR832tGGwHRd8Xd4bX09FDpyj0K+3ANlUZOQ
P3qF7yuDhZV1je4QXg9BKrO9/JRLlSyoHndKqG2onfZsu2918hVcrJyAq6pe/FVDOKbCUot+lfTM
4euAA/p8DghAAQZ3FjisS49qJjfAran+YYg7H4qUmWd+t7Ai+HmpGTfXZPozGpb5Twil6cLPRoo4
iXWthSo0uKzYMaYC0pTs1Xv5EtSZi86AQ8cg3UnOX8knYHgZSUX0FNgyD1v6EoVhRDBPMuP+s2aL
kUDF6GcQWR6R1f7d2zi3BVPbSn5qsZazGtiBiKwwAWfhXpNym2b5IB1QZXsm5M6u+gzA7exbhY+J
RJOLOj3SjqNKWyx9ytUZkyCh522ZQjgW5U4nZp1EtEo6NUKOLuMee3S0BxeW2zyNaPVIpwjGDQKb
HIV/L3fgZ0UezPHNpmYztCz5ZMZ6shxf+6opmcv/20BjS1zl6/KLYzmmXsn2fs0CZQrxLMXABepJ
3N5ObzPt2cgIdJ4nmIDhK/yKGPHFyLngGXCXEcBApL6qR2Z7TgtlAWqbQdmXlMbyJ2MNtrCNHhKG
wHHsxyufuVNIREYOGw7lAOM8vfH0WPXNtRCF5HVLQPgZGGC90Tmb59SJYNf/hv+VzQyzm6KqJV9B
Nl2VVutBCJkhu879JvrL46bCGH9U+WaDe5tbzea/+Y2CFaw9tOLqDpOj3224zxtCAnZ9UkNfx6Xh
lx3eq9rsUSHUP0NwQ5dxNAxSJyUIT+uj4pvW8DJdqJHNPULIwbRthuL5KZuPnqUNrB0LGGpJtlnz
hu0dcNY1JccUzAWhiZnh+sDXqpOCDxzXEyO6OqIL0sEdGSH0sKWT/IzATcuqVT2Xec3XFxH36Bl4
2Gr8VZXE9jW2qBdN1XvAO9X/q+cenQfvQPfGbp3Mn8g3tinxseC0TplH6B8E9GtkmKE6qaZ+SFLX
M/aHX/Q/vhljsyUxD/FzJapYOwS8Yasd06Jxs3p5raW2eSMA5Q50oKZTZM4MXikwMMDG+vWVKEjH
sWRRpnMSRCx7xIoaBfhqFNTC3PsXhTzu5Co07mV1R+bM2d40Oil36XOmfoy5muuJLiA7sZGwuJZL
R/kaaW3mvKc4p3KqgBvTri2fST3Zfi+CimHBU0bjDxLABzO5KFDbgDApXDKF0Np1LhJU2JFZChEW
Nvq/j80XzeYYVXsn+7IYXuvfjCx7Gouwm7GwxpRhL3RehNkMFhJ/E+50aZbYd+Egmd0d/VexcFxj
kKLpnzVyx1PSFWYM+satjybYbUMNwm9GLhF5tf3XwADfESAAC3CKiOWf4UdQBGzPiPzMNOnqmHgA
cs+0tqeYcz0zMq6+Gll/r/5vJADMv/Mzn1Qb2kOWtxTVFHEDoutsLLprbQouR+jVjarjdzV1yjVd
sXRT9eNpzhcbSsCs262ou3f1qGpF30RMKHkZQZHcq1pzVYgjiHfXP00jvVfdyrglZfaz9TNLwqhb
+aKGyRWyqzu/OvVYfVcuearZjS7z0Twy2L/BNzcQWCHY2aBQrNHp0kdU7V8rj/H2bePK4aXeIhTH
1lUC/omwrqGoKtV+i+4oZrc2wCG6b6F+458msdRXhZRVdR3WVf4pHV4IvGv1NZM/LDbNA90VTsJf
Mq7bODvgw1ZeJ2Lfyc2CD7rQMMKWEKzYiD/hyYpmW9Z//BgV6ES9X8oKMXUbdVgft9fB60WuwnyG
Hg1GygM6i4bSDr9N+dIHsEMzzit2FVHmx6zVwbtJ0TH47ProeNEqZqzJL+q5LOn5fMws/qVwnvKE
E5ZOHH4GirsxYqlffUvK5IE8bVq03idIwJ7A57v2E6OXreLsw+FGzfDWbmk3D5t9tsrwX0lGFW4y
mRK8csVj8KePU+ZfQH5cxNmidDhMaUBttzCnjFmcorcqIEv09tIc4TeOX81sQW3HGddinFdshFq5
0M6GpwsazfRnsFj80KdPVSOP80duXdiikWAaLgEGoix8lM1xDDLxn+SYbNDG1lCYcYTo/5EgpIjy
hGnD4rqMIi8m51ERk9QTgSAjMYQqbLb/acIGHj5wKQK6/P2xH6dD//Q7cqCFlCilnJqN7jUlwVL9
kNQmIhfMGn/PK6iCLjS3nGi3VEfO1+fU+C7CeH/Y/cnmbn2IOpJ6/dFufD4b5oNAezZLlWWk1pGO
9GQls0oY6QNZvt4eCycoqnMea+OAvqPhGnTYUPR0Nyq8WWQaggcNh7zYuOWmVctOQha8qhsqOy3H
2Ps5eaMW+LLDfWMcoaHfrDF8gyh1BPKPOFNhKmtmoNRMxKufoQacbmqVfEJGHJupud+OKjta/92Q
e7TUvV/jyiFBFhP8nr5t2HiXsX75xSvEw9gfneLgOyqyRdz3lvb8soTMlxTW08AmR0+Mo51j0pwv
77YeEfgmknEewV+Ugdmf6ZdBFV/CvBZdcHXN9asXytSWyJmYTb5T3YVHy5ne6FQrhT6U/pA3p4Yh
GqhUfOWnEVO1hna4Zw9SiqNKRI7jZlp1Bj1fmvn8Q3kONtYYxU0w1Sr6GMQlEVRzyc11/XTs5KVX
EhBqWpg6CDZ+joH23u7zC7f15aRKwLfCylOtgHG56b0K2LsQ7WnoYFQ9QvfBzQvnhhyrrJKQyAZ0
2oRvPJM1v2GgnnlGZVAGdg319blTZYJARyCNMoeKqbaGTv9mk4RVVFlo3HjOGOwYNASNyyH4DZNZ
GsXG9SWVJyo7cqZcS27txU2YRcuEeRHO3pBL35JFZTrooSFrgV5KvRoWMvcxqxkJCdml/KirsMUR
R4l6f2UGk792dqXRgmq/iKlp5w52uVD0/Q/M9vMg5zUHKJsQyxlEfe0ld416AQo/kuEcxreXKome
YyOFbMLpv0VIjSmH6O7YTk0f1OaH3tA3zfyQ0ANYH82Ol3Pq0VJBavJU2sAUggIDm5IZUQqSPA3y
omTdVmX8wF7vS/iebMfcLwjQRgiBlnLptA0kLyHFnQbLDA3dbznKghPgHCLUmgY3aFDgXkIRCv0h
RTXiEBHeE6zmcar2JZxNAmj4ShxwqvqcNJyvpELBsfJ1qUYKjb3NnKBc4qUXDCPo31gERqHgvX40
pGYvmbayk01xHSV8+Bqt0EddJT6+jzBvqu/Xbdgy8UE8+/EQN2w5pxsSAzf57MNhAbvNUsqPAgn+
TOY3hI18/dNASsuEmIG8xpHy4OoxOOqyBH/q+9oyactCxsqypzqcT6zH7UihZ/lVuqewg30B8DIE
RxeKI41V7Tw8qxZlKe0SkkzBar3WZxBQQFj30BeDq3JnCzVtF5dZbuLDiFGy0DkW4uWDIqgx0BbA
t8+CHFw96rxo7Rl9z9RiW3EapemWmHwnGkEon4nKN/nZq4jtatNVPtF7pC0wkeh9DzK9/byvj3Pn
hTRk24OKHCLTIW8MI9/aznv/eFcFFYifCuN/lK0Q6Jdh2FOSCL2JH7pqptib8dp77QjWwnfkTVc0
f75rrNu9iXc9glnqzizcz/bxzfbepfG+Ug5TTAp8QUH+60qQY9BvaTxNHp0mAZh6dKGz2CkGKwPW
eTuwb5MrUh2kQEJhQD+o0RfdPocqY6EGpsHNYgx0ZI+g7tqxYq8LGr6TgIyx+OhQdasqv3Lve/Mt
vfosLOqp+Je1VJwbBzoLXTyV1DL+a0pJwUIIMw82KDdhKSS01INckd+i79LpninVOnRghGr+JmoB
bbjF3XGVqIRrZyoIBbp/8hAA/Xv6sBE3L/YTkSW+uYczhfzmn4gCLEKMFB7jf0D2IfrbiPvkaU0X
97Fwdjh6xhN/hXEP3FdVnz9inveb/6RxNVHUUHjx3cp+gWEV4/xSey2ld8gqs8zMQP5Il956m24I
3AkeBr/WOBDHAdcRRLsvu34kIB5NdaYyAJ1Pta1Znru1n9DhA7WNp867xLPKpBvhyG8wDRFtODBh
ZlYT9g9cPtuK0ZjPhD8F2pPzshahIcdu6OrljtkOJDSJHJ2E19T6I6v95DOd0ENAgxC5Kpdvub4v
TyYhM3pOmBOBMu3CXqROkZZwRv2iJm1W/9ewt08Q6RAAOGwCtavYAqyi3S/xy9rvbXc1p2jJVabi
1hxeOiVfA9nW4LvBvJG7CeLa5ar6JDmJMhjygYkRxVXOmh6e15I354nbSGDwwvr8WntKT1d+X7am
0zmHlOlh98Ok6AuGWByIY7QbosnEK/dt+ltp/Q24Ncqwm3tlqHwtAYQecOUv1dtzu7wiL4m/SHLk
PIw0LPzaQTL7M3dzl4ygKIVGc5/N3MgcJ6Ss8jAwOz2KbYRVep2HFuCCBQmljNTtBTY3mYreFWsa
H47HMVXMU7Rzfvn1Nr2aXywFAc3g0NM/rYwmEQasUz0Ary7XqAuzwShtbEeq/J+Hs12j8QKvoQYN
qmd/pFl4Kmz106VzzEMmRIedXbt20GyaK0p1yNQQV8klS6BPPu74L4XlfidoycnOPL/BRc40mkqj
bL5mET4fsLgh1kWNfwlWVsDaYKv/e4sZL17tsmkokc1nmtgTFi6x/fiUxnRYn02N3enI7v/UsTmx
3AbkdhT7hwlt5UM8UkXw+zhOQUngdn9MSwU0lsOTfinrNxuzyJOtxk4dYiiys34AGC9HezXNb9kK
GcLJnsoCbWoB7quP7s8JO58sta6n+rgo5B6CwLd089mSW1jcmCE4PzSQjpiqOyGJvFWXyKeP6EDZ
ScHjM/WeKU1AdL5hcCqG3zalqJno5dpttbbxwcuOOfb+XwOWqnsBa1O6jhyrNJAc3kQPDpxlSdRz
CfdPJSbwIoeIvP4AJU+2R7L5buG41N68LVa50meXPthwp6fOpxTmt4vsQhGMCc6GRkjEmEtxjIuk
x+Byyq21zxnWFwlo7HafE0fB5PDRhIUpen3xW7QD38QBrz8s8IKef57CxNU2+1sqIK50Vpw7zR34
++ZSOM8/6uxX4AZKQqfnyq700aQ1f/1VboPXKMbiQEMTldez8k1RhTpLmL9rhANv15xv+fcKVDfW
jKao5s0c8mjpkwErfZp/ibr5cPkMe01SUvi+Mxg7hewE9afR7e70tP6wjwOEBWdGnXzBdVAGpnnZ
IFgMmQW0G/Q9RhesB8ESqDQtBoX8TGIDjaxQCB6FzeECLFlWH4AWA5/ni5kXH6+OLgsAPeRPUfnM
CsbE6JcMd7MSTbTW69+ZxPgQBucvQk/42oEbEXL6E7XPnVa73Atw0biwJpws1HoJww8UwiL1uEbX
VwbYbJ2JrZkomSXsORm+aU0Xn33fNNbx3rEG/60dPtRglpJvzjo5hTx0E6iDo6bcUDA3SzvzLP+A
v1OtRfG4mNW32VgG2KNrUyPurHNeNZD+7U5WzM3FgnIWGAddaEChAbjTrpdm6Dp1qAbqKhjlzDEV
u5NrALXuotlCnmAcqIPmqk1+UGl0VncwDhYcrtnT4phbyxWevH5CikJMPTWp81rwDyD3rK4dYot8
hO+7HD8mJIRhRRBDzBMLOj34XW+q+2I5++rEliARoeJP9Mo5H7E+Lj9NBjrjbTuRF8EVWujfusQv
/rKG1OdicwPg8Qeik/KrKkk1V/KNs0VNd2dLD7VKNpyTFO+G368ZdKuhjdSU4s3nyVFq6RtYnwwO
xKNuShThahjX/Dq9HLyzfk1G0pB4WANwKrbcAQxhOYy0Kd1PQpED6S1Gt8jRtMGBEeonqPNp0Mf+
TeZ04BD2YdE8U17mMg2jpLn4TlXCfNV1LBA8CeKLkzaKrbTA8f6d1CpuOaE9tY930SEMBI2m3Zs6
YTfCD5P+ge4vtGsUFCvLrDLwCmUNMeBKR90oolmhd+ocyQPhMSfEy5d3XUgWxSGwIgHaHlloLly6
WuofAN3ORGy6yfHU+lvSO+Ias5t68XEKy9v8znIOISsi69605o6BSAm/VJgi91xSrP6gH7CyUPD/
vmv+M143ruP4DnNBD9e0T6rOLbJHgZVaivyyWDzGqHf/EUI6U0KbnBybfEdx0b2nJvtLr67pUVNH
h1NkOaNeqyzZel13OofYlQAFpt2T18ljSJJNuiQ0klka3qp23axVMkpVknhsmwJS7petbC+dYUgz
RbPRiKpRJQFYTPfTThjjTYDucKFBsKP37nm1rHbRujucHf4AI4kMYxbV4JxhWbY7n1meJzZD5NSr
xnfyxLYb+I3k9EqfYsS32cx7GsgBTCHhD5ViEVSqdJ+NEAFgyGtnR2u8ZcWFxYgTPWxOOuMfhSfK
nv+QtkXVj2u2YAbO0ZAN2eDCTbzwZWZ9zl+Ien7JG6nL6Kbqe2qmB6yVSul29lBcX3mLIWl8jJRe
/ZgBZVCpDRJErz4uCqAZVPJ53UxvmwbIxFp5a0oTNm1Fa2+/4AlrF/TPouXv+vgQyDf9Ti8dbtvJ
osCm/tmCJoQFKOJrBeRmjj/R30isVD/RQPFK/HoIZMLO74O3PVUj4UKCJ7HIFjTe2ut0I9VYVkKr
2QU+dh1H9ntc8DOdiay+641s/BoG5noan2vh98tLyY6d5Ay1aMKn6SHAN8Gj5gDS47j6TteTSYiT
zFIg8O4bf216FlezDnkazNrV7lkY8FA+jm+hIHlbXbdCyAVJbenYUDLxaxCyf0PtJqk2obR38DTl
3WhSQgw3qOJKEQnRhwwYKIE0Un/inPrcwL97W5KZOk7eR5QsCYZb7eJvp38tP213z/CL/AuS1sZS
NzAZZ/+rH8XeEHapRZ9bXE+deLRZAqFNW6ftml0OEfc6v25tv/pVDLNYBH01b9upw93iVYcJdXTZ
wm9uj3cJWDwW6zuy6AdJ1YiX3FvDPwbqMZBZFBG0vtxcEEIux/B4p2cC2Eo9pNJHb3xVDLk0EnvL
r/93iFQFpYYNPTCIsbwkgraqyV/0bTOqe6tEUrtEjYqvyP6llNfBNmCfCh/HQuIDbVSX6OYRsMtp
DvNfc51B9oiIfGhkowvH1irz5zf9k8baY/p1t3cD42q4Hs/hfuHse9HPiyboJoCg4mQprBmaEXf1
KN3tltfJC3XF/NZBIym061Ayo+wzimJFj94xQzFYVVN5CNK/hso82pO7tC/AlZnvAqR3Iz2E9ltS
8VF7JiVTw1VFWP2/hIVedxxgu5dyNngWFbzOHrfCAwr5pygY1NlcQjTCY9qUuXNI45MtUpDvRluJ
P++k8dmAGRYRw7VPrelyV4lbrw32OUBW4hLMFAh9ypBE8KPYYAw0YiSZqqR9ydZuwQe6z6+uMYSY
gfE5HjfAH0PSspD4R5dycmUHJoLS7MDsaf8EA8cP0zx6NsxtPdSZQarMxMHqNIj833wVB33p2hkL
AWldmvT9bRM6HDCfaIRl5pEqfkJIoSDUyXmSOIyFkdNPUPh4IC4WnhFs0kdOjIphHDnVHiyNpzwW
lOi3bVtiAMLQO765Vd8haWKQPxK1KIxtsUtLkEGSpgrXQvI0+c2VD5ojMtJTHFtxD0ARO65KybCx
MN+JL9incaDs+82EVfsn+iQumwhZ1p2xrkRUZVxDU4tEN47MFAB34Qq9fp8edzYHYN6Z3gkv9Mqo
IxUIlIsFjpV1sDNumoh0H0HcSuTJwaKxsmfOJFg/jEqgsPkotwdoISu2dhNGpLmo7wJ1FyEcb/++
2okeD62t5AfDHjIQuxuTlzSKUtXYAixmYHb5elLhh1Sly6/Xdbyc+GBognWfwQLDjoVNmiguo77g
07fIhOYVJmvcNlPsBtoS+kQkSZUKhya7MWw/KUhIYlVWcTI7CmfYaVm36sz2ocJl1rYelL4S9G5y
lCXUOM/3nnXVfOEVsCwZV/jddDoH1HNKw2vHGlwUmWE0Mve5Fr6YUX15Qkv57m8f7bHfvgUNAQB3
8inRpREOA3p0ZOAAPvo0OegxqnlqGT/W29M+mjpZrS7GyhpTG7eWTOVBr4m+VatA99oK2u7OtAWg
2DZr/IHxTSiRlyqknOjOdJriHfL3t0ssHhphWeBkv/bL4bbGAMCQFKHqQ/4rtdQ2XrKF00yOt9ug
VXXIPggfRqCmnQdx/EWEiYQdfQVaHHoTCPRGntFYrTdRJrrvUw3UNmefxPBSDivBkEKvia91OAWZ
NwqKs5FWPu2svS3jra4rRGjJQcjJGEcXqZ20/O4X1c786NLMEoPnWU0hY6o1Bs0r2gMGec/xqPVr
rlTLkWgWrPKXy9BcyZ/p3ma6QTzApJhin/zE9F7CaylgcGT9Yr2mGk6cXDYjQYVIxGUb0YWcQt0D
wt1HzXnXf3N4eEX73GBqak0rWvtNMKlvs/kZA6eqsupfRnqRvM6d+Wmry9Lk+oYdLmjwKfnm0BIy
+eUWOKs5hAmj4bsGCGFIE4ZHlEk2ORDjHgqlBv9aTyUQ0OG9QEQQB+fPNqrtRGDb1E14MCq7NGL2
yvlGylF2/1RZiD8zu8uj07+vtoPcrCf5xguoPodzLUst+hOxKDFduBDElV/1DZiCw1K/sblK1BUO
MqqZ3HefBVaMejhg/FdlHJc7IVbMdlrlYxgZynfc4NwXfLUnJoBjvNb5akBtCQ5g55GGIqcGZyfz
DhIrJl/8GLBZ6cqIyaBRLsKg4eNcSZtNmvnaLS9S62iRkIDTInN5tTB8ZWmcBTcVTrbybKtcDDw9
02QdGstmiJZucp0Km/V1+sXSS33finoENMmxFlKVMpwVFp2kPZC4hj0xDCdRmF49jMemW0NG1f+e
725gDFKoFD4NpdtEXfZDv208iaowtUIwShWQKGa4q7pHAW4Oj8aUnnHVZq7StHfP4rRyjIhERrXH
5v0+3EfzW2cCKJW1ctLciITmSgxSZ/YXN+FEeKONvS76IVig1OEfCZHdy9Wi8bRPV9yffEZmRyQf
Ykz8qylDSdfzXXcbQ8YSBBDzf99hmsl7hc0rlU3wNWbotzGpJqcGqQFykFPzb/BOSJUbKVThLQKR
BwPetF8JZ5xxUZ8ViuT+YRonnaV9a/Pu8wHwXtEyjNNb3T/j5gKUsa2D5UbikBSBpxPaWkZiMXTm
4Rn2QIPRsujSk95SgSEZf9SdCeIvgFYUVHuDwQF9T98B/Pb7k+qzuJ95D/J3OrzoFbbv9yQmAV2H
5yuhhTghHFvmO9PeduzaXjEOVXtsc7jSX/R0q2uRyB2KVTvbURzi9T52ELWZVYEZNOUVpyzGhJyj
K6HwTifp9VILv8yoUo3Iqzckl4YTJI5EMUGDL6NcLkeQ1JGOchiNMtf9wNnqzSDnZtGr5LRqQAN+
RkHKKHI/Va0hFV/4NuHx2+sgr+fO97W77jbDaCvQDhx3qKFpyKc5jd2kg/6itJBKdVi6iHvP4Uql
8ETU9ZbKGpllK93aQwJof3TsBExO0FqaC+Vu05FvMvCsdlu9LY7DWoGrTBB/FhmiXgEVPin6ctrb
ffU6LXDeZwg9AvApVy49nAd3MTvGMbvfL6/yFXZbajrctBKEh3dRIFayVLmm7xH34rYaFa2RGlGM
4b3BgNrLqJd04wy7GK4DYS/vRbb/SzqI7N6/fh9IpRG0Oj9XnY3wXw0heX8HvNTgW+kK4ykHrcvS
c6ZA6DnSuAZ3ZZedtYyQmB9XJYjFbsFGT+w9+t+x1kXzV3fvxpbdgP7heuQx4TzxTVJM/GvjwGmv
lAmJRQsk7KUaVPdLXuhfUEK9CWs46JJLKG0tx0nQ8ZPkb1NzEo/Y+K7iNhl7FjU7PAvBZTIwjeOx
opT4kHYi0C3VuLcw94zL5dfT/lMOFppn2UneNGthUSp+tn8vtdqKX/FKeezdYncmriI1BRHOmxMT
LXQGWINlB+fcj6Id3iDDC9Z6KVrQpAzRgWKQBWGisI1JujWLxE/pUwRCLi/Q6vMrCewy9Gt8K9tf
1oa5Gts0RAPhBkJbVeADpdvIU0DMbwuoETI9+Sa6zhEBNFXqFD3IYrouiYifksYd0oZlCgAfMN+h
EIDYTaLhOn4ElzbIKR7afYuiC9OiTlx8ibgIzpHyV8LOPzucyC9JPpyeVqhwqjpT2QllNFo02CLV
kGEj/K0gmyFJQn8OH4ggimecBmun2tSsEwTErDIQ0bizqyxsRTDa0kB3RaKYkJMq+DhsH3vwj/C6
Aa0e8FZwh/rqnBAO67JbdNBu1y7tUYlgogPtWpBpWj+B9Nyk+jz4Y5MpDmJWYLgqrY5rO2NR2i1C
Jv0LLzf6Q5MNsMVHvvw7KJOKeVd3O9QCXs6uipRWZqdhV3E3oIsxLQprnFuTj2RrvRdVf02SJKAF
tD+rcx7fIsZD11q6lBSVN8HCjYwSLEHSiV5QYJiay+7CsuwcEJxl0OSv//BA3WhSbcTj1l38v11+
sz6Z9Iqi1W2GsEdeVpuUwJfDu7nh5kzI+fYAEqwhFGLQt9JZMttQEiyh8emxFaIqgRWRiexkNnPi
iEHGJRQmZdpClqrktT0/gcysyt1K0Be6qTQ2kt8xqxX5qZgKyJU6o0LHmaSlDCpHrcaUrOx3sl6N
OAxOIIyA1LxOEAdvyd4pEMbEcLXYuGkvq5JZRanpq+QEo2jG6Aq4k0E74S2sW53OJx9+O0iLfn6q
eJzIGVWEh+lYE1CvsASM4Z/db9N3ctN/pBRi5sq5wpfFJBuxb0itZVDn7Us41+6j3ri5QJAMQqib
Y5ljUUQrYtpjIeIQyXtbcaSW2P0ixIdSTawQotXknXLY7cnnOqWFa7M0Div6EFzLKJ9/LN6ovlgI
wpE7BXJZQ/nUxJCoblJYAZr+sF9c/Kvx+/gZhjxxrBI+WyjoFvieNrqSaRsQ2mvfwhCfDFXr8tWE
pYVeTDfV+0w3ICRVuBpcq3NtqkmjH0mOvVQuDw2Twmkh86jvZk2yyEXDUOS6nLGc/R4hF0zwQU5E
8qy807cXBKzwAm1+qbgXhx4SaX2cW0vyG4Vb3Svnx27jOdyNsreWLIojZ5VkTxJYwcJK8wPYfnSW
r5WNC+njaXtCLv8FQYmR3C5tDMuvTYQiuo4C3lJZJbOY1NAmBTz65qULlmkESPH9hl4KsG4tJ4iF
kaBxRl6Nc3RzbKoYaU6Lr6c/jMvPNSIzhnq2tmCyiEMHBfIfyJd5r4gd4LrOnbkRJkjsdxy+OTDi
5Ym0r82FuB5b5eFlo2e9ZkA15R15NOQcc7kliP6+21HFfosH3PPdN4EybljQvwCraWXgFUAtsd74
9hbDScsjWRk/j3bMX/UCtYYiRzL/d+zGa+s0kbwQcfYgCm4TsYl7PBwYqwGAnCYv6uVkuBPPWcYM
ybAIEc5A9tDJDPBzV1v71qYyG1p3POgNZZW/SHXkt0B+IuETjPmFIbHT4kSyr+dNJ6GdJdxJagqn
+14UJPdbpTyr8sBsSTOWZwf+G/AMhAYenSTssNuWbKDdpHokzLLItL2FRRhh/dqVR3TBX99pGvuw
vEBR1/HXy9Y6gW4Xj/qNJKqiSvZa6aiMmeeglCcXm+lMHSo2NNPMvaQ5hiThB8QPFQC/rGD6eZRl
ByPpduFvKKddC4clipzks5WrlmIwdb+N5JJOOKzdLSnMebo1lj3HKDIPM1VTncF+zjzRKfRzQi74
SsagBuu50d0LuPyTaeAd8sc8L7Fceh9QGA54lERD1E+zGNBYeFOTExvaSoKjw30g6gj7UF6dxYji
GYotlUU++ePb2rtgG1jkTXpppanNrYpiujelb/NFgAzB1dlvyKCYyY3OruFp03YXfZbVLfGUtTfh
GrcaZKmmls9ICwVEN8qjag5Mcdw1mjnCMdopqhgYPDfGF3I0fUJCUuVsD4z9ZVBZPJFDJnvqbsjm
UzviIJyWJzvTvrNljnPtlJiR/T1Nrg695IICm6cfuO/UYs3M1iBg1VO9sJOBEnYtptyaZuR2QeGg
rTqMM+udcdUjJuwN8RjLm4O7uu9i3yI91RJgKyDtDUIWo7vI4w20r31/gNCfIONlLzzHWklAZq+4
ppOgD4JsNfABQUs8uDEyKYJAYIn3HP/z1GLs0K94T4pt9WxTAvNx4AeaziPmE77tfQmEhRLUi7MH
hpSzFqB5JI4aHIjw1o7x9fnG0pdEhtXViZcq6rkCppRkY5q2xYFtoAWexSaABttzdgyAiQccrk5G
8nbiTRzxC6iom/fE/bJrIGaprQRBzN3nbskInTx+DR2rIN2E7gY2XMchsJ1MwdZMOPksqXDQkuJc
J3Yf+JfWfUQ5Wa2USqK3O2E2V1CwpL4Jli4fDc0WdLgluWSmOnpY4EKKshevz2bbBZHrSDZ2orGs
8auhLriqdXsCB6mbcMDYiswHrjJU9ZVkwMWWWGm1z/VjmGjnPWoqKKZYSAjKOIz7/YOOiIJdN6as
ND3JfWbfQAoe+i5fBFNiXqlGENQmkO45R6dE1cURU3awxl8QGXe8LcFMzJiGT39phj2FLuj3wqkd
jHm3naIZlq8j7WY0EisxaAuviam196rSnrRqPmSirDL/Szy57azTFI0IcALR1vORq64xfARobnvC
hDKKsj/b3U5A/16ErBFQQTPdJIudksyNQp+QaRFK45X8aXZdgCKEbJLmwEQUEReTC0YeiUF3427d
fDUIoeaW5ezpklvSVww+YbcH4zWVYMnsl/JcmKpkNrucwpSSv/V4hebwnQBnfcBymKpt0jzLSE9j
2njPZZMHPb21KFVl1ZZmkjWooqOkGhdsLyb7k5LnH1xNeVaiwxXj0iC6OXlhG7CWuAGLZCVUr+zd
TblXoARvuw8dCe1tUhOYBqc9sEYDaNIC14zMG/ZGHltr1upswUagrqe28dvJeK/fxBf8LXECcnGL
0cCZ6y4beVWqAnTjlG1NWnNsm1KnoNeEQlI4LfptBfB6Gbh16hKwBs2X7DFmUaX54AB46DigKpfi
1KQh5q7YziqXIO9Lqr+5nKTlZ7gESmUsDRstOkSdKZJVSRfTO38kXpn6linrSwNOVhJnCr/8+F8D
vI6NwpZsNZ9WWPwgd4cfytsgyA5sJG6RftXXRP+2I7q+WPRuuhcgXbtbFlnD2v9QZs1fH94f9V4B
oEEPnfd0yR2+erT/F+IQ+b1+EIz8Xxmhvw+VboIRrd+FYxp/99lP+JIOFxi2w9vZr6cm/c10uHEo
4lVfti6OJV6UgFnwiTitpyJQArM0NydBNbdzVESRqSwYAoJIYI2VoQ8yKCbG13IPijuRaI1L2T72
WCWwpfbXyVU6Ep7wFUI9yWUd6FPT08Df4DpGdEa4CbkSztXHaRx89UvffTlMvwXj/FQQ1h3O6zaR
3Y9kOx3U/1jiQNYtQfoi49vyHpGN3T/hA/2MPij4kyxv98a/9I+Q4GEK7JLyf8XteNM0i9hw4Dns
r5tKLSZ6109PeeFCqvd4IovknFX/iD4yusLpZ+JYXE0diSb0A8zzBE7+rnCORuaKP4tCQNeAAKsQ
W+p86vciV9+iXNmPQPPwHo6+h5taQVGTi3xDueWBvspXABCXZpvCkK78YFTJQc2/AHDHc3yCEkzr
cubct4/rN0hLch+VXfo5aTZNaNtr73E4pOHe9NIRn+9WYMEce3cNURpAuWrKZ4DVJWwFPhFA3hXU
CKCQONl+SGQ+eS5E/enFP8cDgDS+DSG4ic8xDOalmph7xy07tao1N45y9HbmZRcUHljE1DuozY0J
2HqBIETWhnqdIRbQjI4cI8M25TTNQNskwwTP0IVFodTpvt8SO28boQ0ivLsu76QjokaG3YLoJX0P
LIectXv3i9FCSg997aBMEruXlM0ucGxI0YE+bSpyz2FYv5CNzet1h7vYavG4NX4gypC06g7aRp0n
Kkdaic35usmyG+taW3YbFQVXp3R50FiF+7DcqBGrVkQgz8gf5MNXOCH2EIdCVBCkXKF4k9bqNbYE
zNNaY87Xv4V/SekoRVRQM0GRJR7B4S8RzWWeb3qjgdNRbJmU2L19PIlzDrBCEdRh55bZFtyqU8lK
fYrhy24lSh72KddxD8eIOcJwJNMcviIIosVCuVu4Nl32b5AHpJNk3Zn/EpQ5SW5yfQ/lRLoNonnV
hvszsrLSXHILFzlvxSTU5d3VtCnVsmPWs2qQPkc/EbiIg390Bc9CoV4j/lfn0RFasqw0ku1xPYdQ
GrmhILbyQKRXYq2UkskvD6K3jHV17zgcw6smxnKHaYgtClCtkiIjbIShBbLNnS1zLhrl4FfkG+JX
extviE1k4UBPg2PgPPHYTgYAuXOqfvrJu9qYtGdNPfzCNkllj1WevJQWpOZgaSOYXgXmwE7cZHFp
u4JfAFH6iQ6CYuEUgPt3ELWSJxGl/U8wI/0+5/CPLJkgsuDk9tvdWFsM1oHPfW3TC/6FFNZ0r9Cp
fNl6qSfiVODml4RuOpexHYHFAF4Msug40DK8p1S1U6CgKH9IsTLKMEY7+6wZ9NRP0z4jgRPenVV6
TAPnIyNgAxnH2HzhDGH/xaXcmszzIu6hYUQgeYLwT4Y7P4kK0GZ8bORWGu5DBvoY/D2SdqcmA3B6
UVuZSVBudH0w+lcUX4MTLm8kXnlEAXXBKdwy6V5G8lXlP4qyEwYqd+spx98UBQR0TJX+/QXgpjf2
dBUgIxdOqkNEseFj1X0ZiLPOJLSw9JPqLZ0ddUNyOTngF9q0T+EvrLDZhD8nQJ/9V2Tz1ZkrCbcO
+PFOngYEf9nBKrwZrv6IeaDFeo97/dZYFe+ixkR66o1ztdisjIdNP58Gf4SpBUnOvqEqvqp8cAcS
qLcrPBAvgCHAsyfTxSG+oZWrpON9FJGcQ9AFDkKIKZRx4PjP48mV+rm+PuiJqmtaD2JMRC4ciopH
xqLIhT6xvFb0vpHaWggXoZh/MQGNinrPc88OwBSA2qgmEH1QD7U4MLrJDQIpduJ4HeRBTxoFAexe
BsaTE1uimzxKiquNRDF7abFhxswir21jyWdi/oQEPSrDj4hAJm8x90cK8ULGGUeL2rtZ/jNM0VPP
uV8E/lc0x7SF96iL6SRb87ff3FhfoBlcHL2npgJePeTuYo2CmOcPyjbm6v5e67Vb52LltolCsPpZ
s+5ptQ8/BHKy0iLK9xdltLVbVUStSZV2SqA1k81GG57BKbKSXl1iA61wlvxRWJFsxq1/aiaVK9+j
LD7UGR6P4xNDKvhEGX4kvFS+YVLbeZVehWcS3BH8c0Fyqv00XahlpaWXgkcWHhVeDM3lmngN5ntJ
v3KvadYNX0NwPvBnzJyK7/q37ErUM0Q+R3CSnxCQsegu6HIocrLGoUfRjBRDargKfrp4aOKPYLXY
IzHwdulzjE3zN1/9pY5wPRldrM3z3wXtZd8BeHgauw7cpDSp3GqA7tPK3z3768u+DKJmrkJ9WIwE
MKLjFwv7Nu8n+iRXyI7/Tl/aeWx9jTwzpg7fkFwr3x/H4c7WRAndp37EJrNmrRTws8u6N9XgANLP
S/w+zCdR+pSb6RQQqG+mQKBgSEX/TZMuVVwVzl4yqrQdb+1MaaLDTIGnFEuJJtkZMvGqFU1EwlR6
260WZdSOZla+vS3UA4PZfU71GGaWraVe7T0cUtW9IagXEuGrfx4iSRapxzc7Z4fnsd496qfZgeD2
fb9wZUpydVQ7yP160vxiuUyzaoTlKY+B2XplCFfIwgqqPy09LsNhDAvL/6DdBTI/hKpCU6HdNoZ0
X7fZGMl1EocTqsnuM6FVCmgOis3bDoLnAXthWdOGe2vtZ3ZNFspCoOrTE/8SitOeRxrF6gFQ8G/E
9jVrNp1lkCCbhIWeFjCzpW2ruw0shdq/4fb3FAYUKh09F1rd2e3IMBZgUII98YFYmBdoJ8fBPWUU
NnBh2pWMWasaqS6+lawJLp3hBNWbowxMYo8B5W5vHxrV7GyBRyAYeJZEpjaKEtyrEucfb/8yKrGs
gbvqod1IrtSbjfXdlRLjlnJIR+V58VF04iGDlaNAYcEI8QdiZwklx/MdvoKj3gvekJV7RChjH2Jg
fuc3bV3AtylgLaVubRZASiRtYzUBMYo0Qw2P1shMeqJSPaaMn/UCPy9zODBxtYgqeAeEx/uqCPTX
FyR5Lbq5MWmazhGxeH3pvESS22jKXLgqsxFsAgmbOK0IUpQwOh+MxjIDA3A19Fv5wSPn2Mm7U1xZ
PmCaYQnOFyppCkIIk3U/VRl3mfwjlk0YwDCj9DPYAfYuItD08p3nmAnsBVOLRMpZ05QforMYHfEK
DoDi83X20yG9OFN4FSHNqEZy/huJ1/wm47pU+5M00eqdL8zMA4PSo8ei9HD6Pei8Rq7KEpu2KATE
jPJzQ6zZJzCdGPQvqwrlrWr7FbBevGJLf4Wof81fRZY6iorpCsOKpOOpALVqOCYdcPSuTr7wtpWt
tCWnlXzl0wRx7nAjzXWvOOG1KuslP3GCqX5jAZLQ5dlvdyS1DglE1RYRqV9icomIznkJpPIW8Kko
5s796WchC6jgzzP49+Stsl9dMno3dg02Fh07ON7f1v1BW4R4IbapxH9DHVkDYEKCpll6kRCfGHUV
c4k3YjclUgmk4bi8eUT43gY7LeJSdtZ0dL6qRJHyfienKJfH2sBsyvQ2J2UrgQtJndFMJ0KjDzPK
v6e4mJ9xQOnwJK9++jKriIvT7sdDyIz+0yMkP00hz9unb1d4kpaL7yyhpmHWD1HHKfO58Md0ANTT
wpO7cz06DseAFSdeZwAQ/x9qByV/e2FHcoSLUBksnDf82O/9OphtfMJ1WkgYR0xsNB7lP9ltXHsD
vhmVp/A/Krfl8L7hhWWMQvF4uPmlYwY1VSa2Lg/AHJJu/PJ+MT+wZikdWL2Hg28HVdX97LctEmc9
FB0V++NZJrkRDVoWnagCX3Gh0OG/QjBOCOFDXohOhPAKWThNMunVKEs2D6HqhQK3yW73D9yBXR6e
LR+EDC0lx8GAKcvodbPJ7xF5PkaHxfd7GxcTYrm605GD6ZOoA7WMRTpHtTBIm5VaoXjIZxBRvpJe
gPCDC+sShNpGBGBcHHOGVrPNhPqYYJplsQq4XYqhuCAamfWkL7zLyVEaVX8D2mqMCxyQxODQ8o8A
YTHsl8rnbUDhlcHs37RxZNHuBRvJiiWWva06LhqbhoCAsA5U61WBGvwVXf94g+vc+4i9P3QkQ0Xf
6ZROwN3uvW6mZ1W1yd2KoS4nkgjqwsVmq0IIbJOylGYOot1FfZWY28S2VvtchssKaxbI49m6l9cj
Ma44MHHkYPo5MYO5dzKTXM2F4qN/5eBwh3yuIscghTfh0o6DuAxBNwiww/0Rgqc/J7i21ww4f38R
tLqafDGZjaJR+SKYxpvHC3mtQau0FcI0WukuvONnevkAKk+Hq+5V6NxCKJkUsNVhTfrtwYyBhcBU
AR5iYEiw8hDEJ4VIVJuqkkmG1N+f4RMrvon0COZaQLa9rDgzI4gnbXa+3q0gvpJlPduSGYw3Eeac
kisMfKzbk+g7SXxPytaiUerMJozFJfXualMkfqH5NYq/hd41KvvWzcstPAXR4PdOf4pODTrNSLlI
Z6sOXoZaTjfxNj4YR/x+pyrGXrShV6m1N8uqNSgY8LJb1An+owyA+jx2XsV1+yxqJNxNQB1WJ6c2
ohrfL0KcuHOXY9hzrjMzeTauBvrlETAoGG1KDyP8cm5aQQEmGhEW9cCyF6IyGdvW4BRAJUwswv7C
kmkOVeRQxaQDbKmRegrZoLwHU0n/YdDIHoDie5CnxY+CMQd7FG3MrQdIsOh5fX1mevoWJQCjdx2G
YWXTn8OxRe/4bkslbyE9NOQmyTyDpxp6p2HtVogoFW4RkanCy5LbrXOcLgwr5L0TzYXUVVUVgP4U
vNSVsEVO8qQvRXFtaCNIXzlvdgTxAo6LAZMwnSSSiKIClxzUv1sQNOAq4ENtyBd3eMVnsNP2Pld6
CUF2u5Ikz49blnE1MUk7PSXAHqssZddAGossC+UzdDG8CUfNo2+xLFJ4o3JeD3uZrg26Z8YrKR3s
0GHl1WxjEajdwfqXdkvBH2Jlvfl4lfDJN9bSHBVUur9dqB92u2KjdqAazHOQTvmjCVUftF6tz4O+
UIBHRTGv24dPpm+9koe8jAVMOAAR92qzF4ugbHVcYzmdAc44H6Cgg6jUAEehKIpeUu2hptM6Nz+h
wAmwlewtWm1NgFdMwxhPgY08Uj9OTRE51fYYk6fV3lnGvM8XJ7Fsf4IAi5mgA3VgZZv/0rr2U5ms
se1U4cpoOTpbeBtpFraxP7rRDLtsLkJJ/gV2Fi3czZ8vNimX7o8px1eyB3UPqvC7IGgOB1dgHHWg
j8jTaTwC4PMzbxKwHWO3+IrFKGnQ3WY35GeL2tY+UifPVWug2k6TTZBRsfh/qliKi+Mpsnyzf2LK
VI9zFw3LB9nch4mYmgqrEEztWzbp9uhyW9UY0ej+5FOdUmIwSCT0OW1I/+kXTAqIsHf+ax0WxMYQ
yda6m1c+Ncw3CDlqAUjhf4bPBXZk5kMR7nCUDhBbJO/Jv3Cra7+1HyH411SuGs3a1GdcsPVAUWq0
vR5AN2tsBtn/f/p3/DP2gjZ78Fl4bKGz7WJHk3mHLCCuSUrX1UfbRaRylaTQUhHP/nbJb3mfEqxX
c/p782pMFNAH1oI5z0OKLeQY+X7EoM9MSGtBxsKe8y3tWXl0asfXWQpice4A8lsNRUhNlPslWFf2
Ohlg0UxyzrN//XAWC7e1IO4bDkapVRokWxqyFXGZVlsg2ho0BBMvAbpZ2wl9YmYll/dD0tTVqzRk
OnsJvHbrjpwImTGoviNDc2AVV8a+iaAtwr7C9ecoJqISPaqlCKaE55Hvyz/e8kIw3Rlv1Kk60K3f
zae6V3M2aKoE4urY0zTU6ta57hLXzfKUl561xacShaFvcxEYvFDeoVNEVMTRtSNtcMFhFCp6jyrq
/nxP2KdSmNLSqVLPdi/aCFT70XmbEzSpSRwJTQL0rUmICx8QWAeMntEr0+/dSMdX7KEUph+vlJfV
GL9BlIovQIkeH9q7nrhh+tbTfa127uxorhcWBhj6Kayj8QfbV74BFMafv2W0oY9nbQktrP5gZKuK
z0haq76p7MSiH6Og6RbF/p1D4KW7p2G1Td4Bag60hKodT7wYU10YslW3oOuB7DJxwK8NJp/Lg+/g
umqVlJ7UG++hQVi2S7QFH08f5s6ks812O7rC9nGj66/IDGqVxvkZLFPzQd0wn1mVK+sUIn1hAg2f
WJLK7ckRvkEWT8QsyQijgRRuLNtQo0VMSB498d0Oj3cpGS859BMZwLXre+6u7M9k7BvrPrYGu/hu
v2vKy6nUggCJHQIs0XP62knHvcMGiXwqQIkSJu7LnKpJoTVQeY+3RygBnfswcVsBzb+0GrtfxwtH
kT3ZMDYZtuCTcvFvtltr9JbTI1kISi57XC1mQgcc1EqvStF7gIQ6YDIKkyMp6C5WGUc5rcpB+DUf
NUnzPZOIWYLJ8Zo3JASW3NmykpO6dUvz/xoFNMot/iFr5hoz759QIAfEbxwPRm0zxrq3ho6YYgTV
Hag6PZ7emh5bsBJ0tUKlkIr99N7zHZwP+mXp+IFQ4ipyNzAekDl7hXD3xb84F0YQRs4hneLsBKJc
cW99XRMQLjfJFo9atuYKgUmy/2LOMAySWyFM96MoCjqhqzBh67nzSidylZI/WNrq8jHvvhlvve0q
zN910jbrVN2Nd/rpEFjxl58fHspIpzBKY4TAImndKVBiRBxKN5mMZda/q/uYECVkM6mKQ+Bw7FfE
tV75vJhcAY5+L6ujmRFTJ1XxZGEkzqh4ZZqwhQJi9gWRVplwmtFLuXBwwA+SGdKdXxvF2NtRTrpv
tVLNaWmOIDWt8EzokTGKSlMjttmf6DyEAQfsjxcInmtJw7Cd8dxEN9zd5IF88uK9RiI+ciGsM0iB
GIIx1Mk3W7BYWN1cYmaXkh0AzZHTHERLWDULylHVZoAyHJzzuuXPV5Ih0iItZ6GS+f7etg8kxDgb
1p2Sn53s316F4vpMTjA/vC/NkETG87UhWfru4lUMs1FVHcoFTBoAHlr6vj1QSfywS827XJAbF4pR
1rs0qsoeINKKFPOo58fvkOJLXDo0O33ldHnTO1ZSvhtsj6AMGGqUrSpVPTxDwFHFmcwla177EpGX
a+rb/NBz9DlEHz1qhnY5o/es52QuQ87lrvzgAgOLAKd84qzFtfD3lIYASh9hWK4yT6ZXe7mQ6qa1
dYZ816XjnY2QJAvBKkWHnT/Nq5OnI6Oln6ahNIMSmZVbdXBqKWofAhKhzBtuXW1SwY08OQxnRdGs
G32UGErylnVpEvs7I3Xax4bMSJA9vYpd5P4rrwt31s9cxJp1pAPgdRCgfiHIfct4ZXUC6WjpPy58
qlgTabA0PdwGa+qZbFEsiaFq9tUMcWscxLcgMbOk7YICM2bAaLctpEWrqjrsQVCJCYkW7d7Xcwwq
QxiWQBN1FegJ46a6QDtwTfxNFeR6J6oaXgvswMSN8JrzKY4HFW1HeNx5Vz5m6S3G0HAW29p25AL6
6dcMxi1GdVTnGuVFSVO6P3tLk36ooFKwxILPgQCDIfWVxB4mo++l1LHHiU1Q2aVgWWMJZ2obPVe8
MQcAmNSxxzRuOrvekV3Q+sYkfK8uuLOO6vwMwDOs22lAHRgDdwhL0B60ZESpKYAFDoBYe5aQMQYO
ElOwwS6ZpsCc/7qg4xlAnZQSjtG6ixEAUl4BGE2cBd2IV0kiqtcadG75ofbmOTOjbi8QkjEPzb0L
zbTQ40q5RCPfaNa6bmsT2BWpo7n9AyqGzDoBV32CAlTXxNTFwd8FvKeqQzFe+skphJ+0O4H7Xq2S
oDeKzcQxcRsZ711xcj+lMWjHIVFSqwuu8SZC3vIj8nvl3Vibi6b2jU5Y5rWo+ox+DssyOAKa3r6b
PaL/T6uEqabda8qsGnOcjmzP5FllhVkPPFI+A5EG4pa7vxr182IpQU+LKiJmxzHvcSaOVeAm2TjM
xnx1TiJDXQr78ekeZJHXuN6jtzZVHzvNRJf7CShGDDbKhauH4kCIz4M3qAUO0owNb420RdKq5tGi
41REHTftlkkXdKjoHIb+FG1FwPilgViFunDFPDt6M9Z890AMfozkx26IlNtIfU2yPG9cUnoiFDHJ
tpOc3LSWH5gLeOeOT6pG+Qqx7mb9eIDF3da2+gt/BfNe5vb2TGm4Yy5AblZ/AkHN4YlYnOLa344i
qdsWrVagv+50P7k+A1YTFW2ksQdX+BQlbxaAU5PSuYlU4wMfqkuTe1+ncYr4J5zoHiyIAg+BQlh6
jh/v8Ub+y707sQideMhpyEWHMnfsbXf1N7Dkd+wVlhB19ROwdVS4NKOP53UuvdG9PnqChCJx5D6r
BU7nkyPaqpW+UsE52imndkZitPSHgH2CaMkWnLfe7LvRFaGOOitaC/qxo5TgLZAm4/L7BJ2nT00q
kr0Kwk7N70ZBHWGh07sCBCJKU+HnitC9AoYwflsnIa/+TePSJi3FTaToqGfI5DA3ufWnZFYe8xFM
Vn8Tv1vUCeq0vgOWChLoa0rL1yNEyzLTBsLPXluDExztvDhisvo4NE06sI5qBEn1aITSXocqvyiK
R6h+RnNXtWW6fm103XiaQKa9GNMji5JAmizXSKQxL3+ELQteJDT8qzSDn4QQMjZOhSXe7UAnuTwB
7HFNwQXY5aRIMGZ39AnykHWqINP5YttuiCrP1xy8dEVFm0/sKIkilq9M+pg++HuNcyYYl6RA2d6i
fNysQfDMWhRqYAZvKY+7O1SK9M9oE10rdN7J3oFsVIzx4Pclbu2Yhz+kfYCCLkjSc7gJmPwLA+Ss
pMEjcGf89x+OxC5SKhfh5kvAZacEZBL4VIVi8cxgRYWZE8Fv2xRKIn8i1kBvm65BEoSGc5yN5rZI
1cQQs6vw+xi7nXxfElfajpk81cXHqvaux13hggGo3nsky8I4g5Wc4VOK/dkm+JaaFsR7doz6TYgW
wYMylwANLzcq7LkNHGhoE0zhRSXx4NDi9v2JUT6kUtQASFDwPibHEvCf5v8L2GncHOB8rWmrJID/
GhiZaWd24Lkd8UAcB7hHm4xKLeLF0fXGy7OoKPNbeSI96KEQImRXzC1zQJwreLaBhV1UPXjxE6Jj
ajM73cLj/InxMfTcWcSYnH3tWiuZok3e6Md0qH/UkAFhBxO3bXG3DvhfEzmjVDo7Obn5PeOvHrGJ
uKyCuXPYrDDZpAv1ptL51hjVSs4zLzBV0SJ8pCWyFh2Xj0dgWTQU+PfM3+Mg5mG600B7ff+Sxpqt
HqnHC9UtOstOfJZqud+L2HA3sLTJ6xIyUZK1jbRTEVuq65gPZpZJfwzBnSnFYrKHY0QwZ3PZF6vX
x3KiY0GobdY3VV5zGzDndFExQL36yyDuIScOIqmT7ojLKEdQV5NYWKWOW6FmYbIDlQ1gTIzRnzZD
C5NVApsoCtE7YwPfvp3M+l4e9XMSsXwszQvPKcmcPd/HCT51bGNPPgt8hq1xD5NVoh4uwmXLNNww
chtODRP9IXHnIBKBch2/yWWhHvLQ8PGLGi6UY+9XaKlUPNk3mKR620d6u1RHRNiOEbdBX3BiE63Y
eP5utH3JDM66f0YfToTxmXC5u+4p8rovYXSI+yxm/5vWv6rUoW7xvkQawGuk6OmMrtNq6HQVybMT
DKbSWVLK9tnxYDsoqZeKzSqUbGT3OjdtwSIEEUCAdGSgN+56nVHIx94HMlp5SXqXwrmrfiDtNwkW
sSWGs6THyA0/LSqDXpjl+9dC1Brf5fSIZPvLFWl/JRlDvzyc/l9CaQQTmobkJZ3MwAlcMBFpkXtM
qwzHwc0taDvQr67mWPc4VeWlAs18KdNMS362T3sqEWgXmGem4UkCXGwUWAV6B1I9i64WY0RsbXzs
bws3YN6/pGpWvvxbEfKOWvvudH691+q8vZRj0chlSkCqTUr9hlyJhFCr6lltn0PwPber2Imiszeo
Aiw5mKo4Dq4cmknU7NIlO1NqZMa+qsxpR5BqrysDFeLrsCMGXj3dpSoyCAIspLCHLYdvVRrsi+Ec
/Fy31gNmyC847u0B9UVNn9QcheCyj8ZBGMYfqTIVYqI0U0P60dswv7mp0ybJ2OM2UViLs1MGtSnM
ETl7FXrG26uqa6k4DkbtN1zhwhMdIkoin/u5BbuWUCmtik58pEAtfAg51u72JHmJMNL7HwJVyw/E
SvxgXype93X+jyuYuDxL6ld1JkEmKOn+dOG0F+/h8F5fkxcG9vfTFvx5hCMzeFw2egzY2WOhqQ/d
pW63lsEwHIhDpMKb7B2RnlJSH76f+jgSNT5+2X1CbA8S/EG0ZaPKEGGWn7xGWoc3S/2bYPdQJM6P
G0984tM1YJ0HTtmxKK/dx8X4JFCCLO0hvcXKLlvrzUgXA17XYFHJtSIjKRDJACF8CkgBiN75iynz
zeSvpJgS2m4XaHlQOfYxlChAdueihlONY3Ewt5jj7wIPtBiCImJtRbRRDGT2+Siwnh79L37wQ/9Y
vT8wkEt1wYLoU7+wrYcN8YHQdRAiE8xc8Spy1fC8ozIohebOoAoR+ZKJ0UCyViAuJm/Eslxwx6Fn
QtkiAlIU7dZJ36a/k7tXtQsqzo+1nqNROcCRQJwDAugkYJG2G01VvUmzvmcCQCtZ9+aKOLo902O7
ffX8BPO1+obYEu+WNTQbnprXcXynh1UmiAoQwxfkRAW1UNmEUr8IyZxKw16fZn0qqgCpBp2UtDPX
cQYjWdm5Gm4M74fEdleVt322srsOpfrJNj8UtLY4kMBZURA4uYvxAYL4XcBWpgveCq8uDE39NsVx
1diPAMX9kKRw9ulxNnNSStSVFPf4Uf20MuXxQIYZywFtRvhPC4Vsglwrr4Uf2uw9WuZwdrQSUKRJ
bz7c1UtrSqL0N2XLTdPLqUT2eD9wd9i+3dnxb8U8xt9ZGBBAcqS1TbhgwN8O8+bSp20H5pHB2oES
4BJLW9hgS6or+F5fxnGSz3NGv0zR6LGZvYXjP2fmQ6donIR32PwgK+ToTiKsQo6Zyek86C69bcN1
v2ktAIj/gmb6cvHJH2T+a2F/vZ1NC9dpaxecWcVNkVKUwd1ssrWhBrTCPn7BnPmoE167dDXy/ght
OVAro7uL2rCWXx61cGwYmxUJXCwhRN99gx6fYSKkZXNRryTTDbP6hk3wRy/Ks80hgcxjcqIDKlKt
nEnpy28Eo5kaCDMlM8+5ZUUu7of/UNJ0yPcWdwb2EkR9ig04qxE3ERzyP06+8t1DOutcm4tbkoD1
t3aKdAP2NAWnCTE8RyEb6i2vZVtG2AKkMfhP+FyR1ltuXQMfKe6kKuXfCEhc4R2ljpRJrBhoLzFs
5RyuOJsg2ps5cbne3KsMZN1YlyYS+iMkmayTCHB3kvnstcm+okTcnK5oPH68e1lkuE61UmfJ4Xmx
tjLqmNayL8LHAuIAQ6kwsCdmL6ToNohS9WFbK9eNzQ2aWQ2cfF7LpbgrhYMqY6iGd2PA7Gmv8AdR
eT3kr56c6/a92gZ4GU0kZlhKAZ4n6e79/ZuKSCPGxEtC0dIBjFpq1yHUjWqOlP75u65OuY4g4hCt
yW+8Bm9XL+0ujmhkJIfXwDJVud8ZRrrFlTJ7k3gMhXObo1xgFgAUxINNzki47P9Dnl+F3TrWqa19
RqeFQ1RKMERX+2zF1gpBcWfVFuxaiH6MrKZHqU0QtKdFFx4GlyMrPVzA0Q1Yj3y9clLsPSBjypzx
HRtT2NNj34cYc6C4WTtIfD2uUUnKUw5FXYhBkEXVp7pHXMtzDZJnQjU5VaObBMIRYH6FtNGjy/+9
47UuoGZZBXlOSoZgfaCuSzJK55fI9hyNZNynrqwPtai6BNrx9rYLNOO9D4DwhO9BtMJt4sKQikYa
oWyIxMx3oBkP2DbAuwlh1HDoY4FsU47e55ImhNIi0gvW65DnJYmVr9dwA788SV56iz6VaVax9K/s
CYLR8wqbthceraH0OBGRHZUmfta1VlcfgwceV8G08/oWBARYIR9xWIyNeC7MagAZmntx1kA/eSkN
VIxfO0Sm1N2SLzoh7WAG2WQCpsyRKyjKANZNNLMoZyKkAZgXnNoKe/Om2qUwinfEaJ5d7h/YLFYP
CzAqDzLbpJAgoUjRjihpLyKi0xtVyXjGdycjcLvfBlLo4yDrzGxAyjsUIN50nrX6cNEchLS2dgz9
avTpiK2pZGcXRjcsOC/2FOy8EZojUvAolElGC0Qd2/4gCBJmgxXu5RxCP4unaUqAi/mNJmajR4nd
sZHDYgQ4dD0LdvNHmwsXHf5obMrN0E4HjYskWCyIIX7aazbBSw1TUkwC8Z312yRRCL6ejWniNMki
W8WI8ZW1T2ppp0oJeNN5rO2PAUp8DFpKe5Xxr2BLKwBj+VUXRyFZvGUZJfFbFwWmXCWOpJoI2JS5
xhmZXh3uSgxEuJC5AD4kobBn0m23VR0z8yQDdTU31azDoZwCXKRAIpcoZIGTz2YjfHKzzRi7itww
iMhhr4QojQsPa+KEnkkKhGPmvlEtBNT5eE5bUdGftiDq+SxYLfkUIbigzzlW+uPylJMGRm3OGx3a
sYBd2R/8GaHLzgy8zX+3358PxCPCuuPbYHq8IFyybJYSeT+kkO+AgwwDj+mc8UAVdjqqPfY0EVKk
9moBrZBlt/8xz1oVZxEC+kN87Ner8mQ/7MZ/+tu10bdLIm+26pNYpflTuxTy6a7TIisGwwaiLs9H
mV9SXdqyGZgQzANnpZiPRJBGP5w1edbG2qd72q8KjxcZKBTlbh7wYpYJruD1Pcc87vxZ8prry7lt
X5c2nZmjYAacM1Mml0hbHgaxQO+s5Znx/ZyWyKkU+ZDgCjN9V0O7aOAlhXUzLINaCDuWNO2mNvUl
itVjRd4b+11Vn1Jz+FkTDf1BvARWCaMCu0ImgL/ZHr3yiinDK0ODVpVBG5NamTYKdD9dsA/1D+sF
mV7Zw0k3feCApIPfge3PU8FwOqhtEuKHAy9pHkjMFSYWSNkhlYcoE3uWRHUMQOFdsDppAAMf6nSG
jO5hP2kiBzGESb29O0jShdjWrHiwddsi4DXp0hH0MABOxmqdW7SWVQQcomYxBA0v3M9BBz7+xpTR
GJCcbUTixa1X+Y/2ousARKEOqFk5a0fzHPFYwrSM8fmlbZd+af797qysGlq3e8obED0zpAYcZPqG
RpcbaxYEi2/GHblT9gurLCo3/o3VxENPmJb1A8EvOCvW3t+UXlefJzpL7MaSDOv2d240qubCdCPp
pnP8A8hweqxVdI6TfcRuTNkSevV/gXQvpbwW4hhKUMBuU/q7yrXdNBIvW02ZyGcAcSgsA8Pkz2M5
gGqT1ZQtHpNx0rFvrYTHVpBG3eFjauKufwrKCTguqsm/YGKCgthRyLEOkRU5xUc+T65nBayGnCzG
Ip3nXEr/gtKCCRjPF/FDeSAvQkWZPg39x6jFTEsZAXLlZzHu1D87ZHrgcgrxXiTrkmbdZuU6DtFB
yph7ZV2zmQIUoJokWhU6NS/7kDDYgkKaUMD3JvegOURjwVIuEF4Z3ZA+DuFiOlIBjpWeCVXRwCPN
9RUuLr7H3CzaIuGRTdTheL3vcJYtkadDWfxQVN6VhS1V1hhPSNHQKdLFnAy88P6uObBmEhJDyZXl
c/rMRdoNwOMT3PDd13c6J5fgdMCFSIBQD76pM9AcAF3+luuN8LAsJi7qdvV288jGauCl2OUYSn1n
saO7dxIhY2w91LB6Yy2H0UckVBo0dsVbmLHiCj0wza3WKx5vtaFCaHc4RxzRFyg37shggcK35u/M
AniRndFGD3tmwe7JfabrB7otieTUdyBEYA/pim/mJ77MdoQNUcXIZrDBMyj5UOj/YQvAb3S6UZ+2
r8RQGSPD30CirvTcDGrxM8tTGI2MmBuhAPKYQBe+PAFLldBd9xVqp8KtRn33MlNQvGxwpZ7mFi8Z
YgtUFjQqyP9Gg1G/SOrUSwGzbyr6jJlDp0CQZo6x0jm6g9VWMD6DcbK1csr4+1ne7veQP0WFyePr
7ScoZosGQS2Ju984Kjtvaymd8qGb1rtp5y6DHHKp/b3FanIeXYjKhhCit8g6o8CaY1UmjESp/TuU
qwxGRC1CD3/CmoGA8CJJ0L/w6dwflJapMdxrQuV4180kssj9iJ3tyBbZRwy52nvcUAKmg5IuZHGE
dc/wFDWd2UhgPC4QouKukHnjfxqgoxYrswdAMd5MiKyTDeB/E1G7ciN9Q3E+InSl2vYyZEljVyIQ
/wPQbk16uZ9ZSfQNsUiG36YnQh03PTUvAY9oBjI1ucRRDLRIBCzc/eYKvuK6XRl1zEyQqFd4m2kY
mFMelBJyveUe2UPwMKEHvJzY2GeMTJuzfZk2ypMwjOiOcSWyQ31Vwd2jId+ojOp/Eauh3tZz2sHQ
ynckMAMKfvlRR09UMGMgSPKvfgEl8jPVt8tGEAVTERtkkAYcF/w0pvqzJjqOt1RTYiJnmFpGFR3e
Cygnlg+XKi/W/tcXbUxdsn8m9IYETcAClD8ReuDftBlxJTDGKFzHvWVczRUdy8Y04OmRN+UrOOz8
vUG61HtzcJ67IdP+ve8FEe6vYO57wAasz9AMHA6ymmrntp/E5LOHxrbIOo5kCHsSEfljnISnTIjD
CxDakZlI+Z5SqoprgSZn+Zn/BXLyg8Vz/IyzdXK0qPo+1dLIH5ie/WLUJvoEyCdLfzi/DBVy7Sqw
Qy8kHQkRt/aOtthNlTGMYfkTMeQ6FSVggO9y8KR6Mn9bJzRAp3Na2XLppEUKegQHGhKl7KWEoSMx
847ZHRs8MuibT0A7oVyyYCwPqWFYBgur41KsMAia1ofOlTeutKOr/pQPNrXaRpAdEz9EQPjB0iqL
XSrftuGSiLizMiplpQOMVqqVyy74VJzjukdv2kJ/gEntakOOpKZS5q87vo7O4c1/Vvj0hEJsp6Vt
oGCKD2EuxdYYEG9QhbhiGPr0jUwqdrKQlpYJrvzRfJH/yDV0wIQ8ITdns5s0Us9oZ3BxJAOLj0GN
y2gzGA/R+TrJ0DGzf9HI6cU9NrI5PJBe9FyNpWlHLPgXmqGBWz8Kpg62l6aAXLTUjT7yBSdDgniD
oKHhu0psW6tlSldkU1HxDHPbYfU+3kFtIff7Z/efFmRjdrIIFpgZLkOgSOBwfTVJiN/2hygi4CAX
2Om9JXtUtXc/f7T/KLOO8Z+w9NJZGmSGOEP8vPfldET9LPcRLm3XE5yCVi+SR5LjLtrxTdRmYfQr
VnI0jXoyCGZnjX8iGsF25wANAcmYWOU28tmO3x1aSH7abWaxYQTIShpB5vqCXaUlGKuHX8fD42wE
IWtD8tbJ3whO3j9zlW9xPJQ3kZCxoN871I/K625NysHsn+M9RvDsn8I0RJnxvDfmqSkOFOJaLQDq
fPZTtlSexZRKySVoKeCZtZ4xMnPaOJbuwsNFCffMNiu+ioF/27bo5xkeWJtfKnu7QXljFrkSX+Vn
Gq09KrG+IJ8OnWZeUKNp5xYVFDdkEvxR4XQFndq7PoBWSJvYhlso9aAA6u+ehCykzrscFYO+AEZr
oFWuYBrKnY5ZZZeEI30SamfI3iJWVAwYfZOTBz2RBKNacPtf0OxeLxKBaNtUpRuYJDDXMg6srnkv
u8h045CqobkClKPj0nq355JiOA7NLNYdHn1QHTroIhMXsWrsIV8vCpvdCQxdGkz6jQl7RhoxoCqe
xg8FGwHK4bnbpxD+zbnL1qLOGGZY5PJwV2wt0Q0ZiOUxprk24zusaIx7z+G+AAQZhbh2CTxh65jJ
S1cjgXIp8UuJ/1tCh5V3FdN4o/xbw3GY5FGFKwGnNMM/5lvyZ1sbCa3fVty8AMkaLEJDvHNr/u4j
LyvRLcLEQ1rXjolGv4CtF+v9qePitR/DOt/oWinjwiIHVQ72Q0VzBnYn429uJsiyxWHV1nJWgEy1
a1ZreQap3ytTa3Yy2gm/2j1tr0VZJDzM04FYGDtHmEexgxY/w3mGy68xHfHPSLC+op36jgkGsfyT
Yj2kkUX0V3lE/qcp/MJj+vVvKQhD2PGI8Dw8g0I0dHQS1kQnFQ1MltB2K0vWXG120t5pywj7xoIt
P3tSfHw1EHvVXF2TmzyOYFAO7qMhjO8G7S8501Fg3bvid8igBkdAmXPHMlFYgZLIhHkQnjIFaP7o
woTHrgUy6/c+HdRSmR3e3FQF/R7ozeFE7PPPwK8I24WPMiOARADbujFd7OnC7OKnL3EIMWfESNAw
+B3uJnwmSFIbrmZ5v1p9lfqBcxOEwZaZix65ob8cpd0NlLFR36jLeyWbdRwW1Af2lLgN79u9Una7
UMQLV1luFQiic4BbMg0jUT2YOO8dm/XSoF3C1fWNnMehKiUxmQBTSOENWRODLV+LlmNQyOA5x4IM
54f6UbetgPXJO/CyH253zcBRLw7OSNg4HB9x49YG4tIXW5e9NE6IXG129GN2ae8NVZqnLrJnXgPP
RsVQMTM9GASpSLmxhCIiymx5AG0RwhEGCPLZBbM1LEBtv1vCKkDK3/rSHeooDMIDhkBRdJUiX+mY
q3qTOIxUaKx8i6NYUG94TkjXCb017xHb4Di5SA3AuW9iw5Dr1p8jJtC9cd9Jlo1ioZftoybpKDnJ
/LJEiq8eCba7lH0iJVHVmS+FIIjE85wcApaA43cDOmsD/bDGnbeEtaI/Ziy0FVbsRz8fP/gnFhIn
jKwTM7vSbKiPlzfa0qgTcKni/BPL0bm5t6oihcX8ZidHmYOjm+tPkBo9RFDLojDN4i1884sZK1zE
R+3VKknPu5Z5zb+ZfI8edYrF2z9zrgTuEkTEJ9iWXeJ/mNjSCAB2fvO/gBAftmIiK9tqeoNh/+f6
wpC+0V9NswyKojsNcNtaWnqgzPeECHkH93gjjxP/G927nsripPnoR92GXVmzUeaGYHl3IjWOrZuq
CBnLW6eIGu7q5AOedx+Gw3594x6+HptowR3kQ9Xxv9xaVCR2lhOpbpMuHn2C3qy1rr5iyQVNlIpd
p5X0/cG+bM9VsB0Z77aZ9hBI/4zFXhWLaSe5JJPRJvjUDadvrQqZSL2XHGKGXjexDULP0nubIwPR
I6JSbD0HB4Mk+0gS5Gyw98zZfJElo0H8jZzdE3kvUFZMiIdivnavddVrY5UBuxJU0Bk9/jvOFDbW
+oUc9JLyIXMnZFZl64zM75d0og/RyNEBvGDwQUA8Jwc38m7St5e8iaqUq3jE5gTxSY+JIvQxbI0p
esuIVgW4+81Nz99C07yGHR76E5O6jGK27JTQnZ3C+LTYcur/vAyQrMCNUOhPZVUeKcD8okdOevIY
gj8yzN2mI/BUICbXiq/bOUYEeHMAhr8ZizEUnm6WaumKYdAz8zguow+uZIG/FYBGuEldxk7KDinw
3JNV0HApeL0QprrUtlEeeK3jcuhOkYq+jUnY+s6cdCJkckqP2Oyh+/AtY57X8/AqVbyIbaTbgJFq
4QMkR4kx1o7F38x3j/o0eN24P15BSMwbKV1LL+STcmthNpCDSxUJEL2LBtg1/+DfXMJ7GVoT82KR
rLmgRrcG+H64KDFfaeoQu7wU/JmThBITi4JwyK+obhJWdjM+2CIm7hPtXEJlg45OYGtX5cy5vNvg
602dYTzjLT98Gb2DZqRoI7AUDqeyQh3CF/PE36BjDKbvotOOk3GQhtkpje3p0dhG+dvOgnXijWgB
kZIvSIxK1Mpc+iK9NNu73L7o55duIctIglB2tEMblWUXk284h8SwZuJ0pWF0RBd2OXCY+XhvrMV5
G53hIf7mVmWDvo965+7r60dxTJZoAaBkWDyFLofcJxKQJAAPTzFGD9b611M6cYyuw3T0HuA9j4tO
Mi35UDoiywcjTiRnhf1KAaKY7K++vSo4bLGHXQSG7WjboW+pTjsBaO1Rjn1mMKQI8MtI7nOcv0Zc
mFKWZctHreY1BcksUXyXAo9xW2wfA19OxvHOdYU/i28avDVzzP6FbBEvkAQ6sjNZgYESnof56YeA
ZGiFpeZc4PymlK6nLhJack0d3yzvTDwyZWALSjG4/gROrFL8uBSsZCl7Fck0err9UYN+9xc9XTRm
w+rmAAaWWrbmdGhCxFbUNCK0sYqBPw5qDPdNmCqmrdgy5NUqzik0M5DZfSae4dhQ9iV59pY0rMdp
U/FIVxrBRUrYBqc+KUe42V1xDMVX6BpllCumUWZgnSG3YOvyWbvXhfTOoSu6PRslzakZwl7GwwX6
9Ogb04muEggtsLxI/cRSgeAl2g0V8KelHXr/KaYJ/w1EU8WmmLq8gtncJSLI7wX13QmWb78CdhNy
hLIovlnOFlRW2aoyG1bVNifEaKuea64jVLJKwveaEOWYVL9QH9/w7Xs+0xpOJJalk0PtSgcxWOko
i4jOcQz6IJZCbCTCgeiuvFkHwS7bd/U+UJlCUOxGumD53d1okoFWBThGi6be9ImSrpMngwO8x1hE
HeDLmuer0Ev0f4qhZsz0mUPkxkGXXZ75EQV0RNiNhctbYLT5piZn2gk1Z4a0u9cnqmyii45JT2jt
yoE7/ZzqNfeGySn8hk8aOAnir04HYA2imwno3XkNmif4MVwf8ZknShGFoBpDYoe0uh9Lg30Oi3aC
6J8dz1OhXJz3a/Oz6U272AoEA6khpVwTo1etjRn8vOMsJlP+eVP0HZ6fejdh/n3/1WOhMG3WIdqW
R+5AAjAEqQBCJSVrgC3fxa/+0XRiKidINzXfLXJqzi3tsuTm+zj3Adoy1A3VuGCyzVa4pFxXu+gK
tP7N/G0i56d6Lun9xC43EToY6j6F15kpDVueoAYZqPNPknmUnPz/YXjmpA5j75We7E+GQHcf+VGf
stboWMG1hqQn5sWBoZnHiiaIWSE7w/j3mYDuyEPSL4T7XLVsxhSLM3l70b+9sUsXk56V+MS5k2aa
hww751TLg/HlUQLSE8uBMZo1GZaQtbaOAe1DmXidAp0XFB3mnPH5Sj+eDnDusutJxPSkTx6Vn3dz
8XweHMhHs5Ey8JB4Pnnj7VzyLggsFJYmByPIyPpwS8tQG9BXAGIgpB+idQaiZEFXXwRS4H5azGh/
Rw/EPXtoL3Z0JHIBoKjZi/nTVsvL5sgdmfVqRWAjGrjT1tK/uDDNiPIwvzxosG3YFrGA5UsOs2vb
WkT0ka5luf/9n9PnEy131xuaT3FM2jSPXy6cTS9Ahs2fLFAOCuiCqaBq83a3k6UvTMzI4gm/zZJg
bGTKNOEeOCKvGnwdJbhc1TRGhV8xKkmt4P0+d5v/gf5XQnJ+zz/9g5Ce9Vpy/MTKm/Udm6uoAdKJ
O3T51ZmeQjqoxKDJPFRqjyzmgTUgl+d88dY7KqsfgQaFvxB7/x78PvJtCNwIGudCqnZji20wsgli
4PjlnVGzc7xILoBouGOR/1Sg61XJjO7YLUsNGNxpGzmtV7+6Xs8v0xMZkYpBAYwsteh3RsSgwOc+
rAteCqwy5+1AkusQJsvcYYUdPMlXU8PmN+TmFlez7AtCiGiDfEEgtgwq5AI5ZJgftDZqyd5G8ODI
QwNG0tp8uAdoMokxkpuQUDguzGfGtF3HqmNHBHDhj2RxAMCv3J//34q2R2QE7pSXpYE7UL97e5gN
SijUvlEY0D0IB5ueic/DpF3n9Al8+SFqCtpTNwuN8KOOPTchvSh8pcyl7OzjGK0Y68oYnGI3v1yu
BUzUj9wjB0J0KEnVcJuQLU294U5USZg/ylss7TgzgT2BMWUF7IGM5I6FaUZhcKsFQGcm07h2/DMt
OFHY1+0narkg7H5lI33WZzCsVpHW9LPfS9S96/6K8UpqPHqMgLGy5Ct9ZAct+fRdDo1XW0WbiuLD
u9p0mzftmUnnRavt/KNgGeHRttVEEngYp9+QPxgsPX1pxV//96jb2BkGQ8XgbaC3WXCEA6SorLAY
1It5ObHNxgeOMKj3QDH17pMkqcppD2FzjyzRqxVyyC3/rOeOV2qkGq0y6VY0hri3Oxm7kv2w52iB
RSTeIFjVONoexl++SD97deL2DWoDqA/4Av8anw3zfWI/8iqo8VlFFThpHeBClxd+OgdoOEhvLq/P
tiU362hbxYVIRpUuE9Ld8WVhB35BzTYXQ59JB1mUqw+XElU1Cmz2NeTrYhgtny+uKgwfD1tfuNAx
qh54wQx2ZTVInuk+K2IhwQd7MmV00SdesAvW/Ck5+iZKz7jd8Yp+rrMfEY78jYQ47l4MRv1bh2on
UE2ZDwJDAYBzODqKlfR4UCbChom2/xiiqQaS/71AfFaXHU5cjI6EOmiXpxF5mQwVJ1LKtDTvolYl
MPmDn2O9/Rd6K7CNrAoDk2sIhKYfTf9bL78sXQBqYYhOTcyZ0I4cPd2feKiFinp+WWgV5e1973aY
eNNlivL00WKRSQvyrAloUfd61BW8GdiNrWyWFD4tiYsewWoUtQUCK3ewPK9Sh5haKd0toNOpy5FR
P0Sja7fsOk84d3Y1aCP5+0sqxkMGJTCN6vbdZeSg3jASVEWwhjRJOI9TwW+6qKp6daiyES45/QS8
1HSBIyPCDbybnlwrmCAkpY06cb3btl3VfCJO34K+SUFLERvcYYiit4evnqafWcWgOU98gMR9hyKt
URX5nA4NQB87hlkrHDO7DhoCghcxcn+/5SckxOhxpmh5+4lhUMrgUgb2leu6bKN4c8LyT7DYdAw2
OjulPRmAeFspcu2JWpn/P81DvY37JAMUiXnBcD1HBljWP814c04FPOfkQ8bddncIudWqqNNDId9g
gszvvbv8+tzEzjB5zQRqz80m5QG3Nse3759dN7Hwr/bmhlE9ZXKB3mUB1hMJKU2qSGK92jblESaJ
Iq5uSscjy7ZwY60lSJDfyqlDPce3RlaBNdV3135S+3tAhPEcPWjYqPP3/g9+rCh1ve4yv9aINJ8X
Z5pKpzL58kl6t26j634pw0KksiqjQcmlgo2xwpCitQY0gqwxAAFOOu/k+Wbnnu28rZTxGw4K7R3c
iqWiRHLftPV0Qq1aGfYZHZGs9HhSxD9vxQ5634r/xzSAEc7rbUZp7ImO36JtZ6tHC4T0qSALsQ7n
n3ryNU+GY2AYQ4kaDSYUDGLCRGz7Hf7/yNUT+dDyBlUO5wxK+jE5co6/aOrSyhEoLBj0JWPd+1fw
VhUA/fVrrsrjTszRSDwNVB4mg57JVJtw02tf5uw/Y/uzr6lX/PheQvxSXKctSRWZyA3mt3oIzsQA
mLc+d0HTgT7JVkX8zk+L1nUpc6GAt9/dzbP9BxTgiKa5meGDtjxHUstUyhByYVjcmHBdwRx6I0+1
COTWKo2umS2SKlWjbxuBldzvdja+6Dbm+tPBfg0SrDVYeSfwkvdmRfkaKBMW+2yc0XqwJVTE9MZk
xBBWBCj3nV5X+4N5H78kX5DbN5T/i1+UMwV9sLJ5BzXCGk7cP1tbkybC72tX/F/wf2B5w5t3ZRql
t5azk/79iGxgn36v5j/vzLKc2aTt7PizqCo2XAQEQNVACNZpJ4HqhAP7Ia7loIshJefSs24+cHBW
Q/YkTGIIKRm9SW1cUTqyl82AkkPYM2DIsFEF0Br/X+5LOBASlIrmCXYtkou8S2lrgLcglRVaEpZl
XVIwpJeqfNR3eMxC4prIaq7VVHFCUSSohNHRJmhdQqXKsQzaomnBKmwU7X1HOJNcLyACkngjvUCi
K7DFfx5tMzwoIGj8RDIp2hDStObwvJZs5gYw8rujZ4CQNc1vpyY4HDz8A0DxkGXiey6ID8kHIapI
6cvUD0IXbxlwr1GZdgBeAIjyerbkWBeYhIiOblrQ2KBp2PkDeOHjUFeu0zzksJSqo0AA8CgMpNrA
87GichcNsn/aiH9qgdEf9w5LZmbWhfV1Lcw2chnpsM/67e7rO0+1A5+dS+mvTgic0Xrk1jPslEHK
Fx2DSVfp31AMGzW1qjvgacbgOWPygMSg+G1ZMuaI/2F9m+exUAMWPwmMWx8xCNa30cX4BvvkXbdb
Op79QLjIjGRB20EFqp+zjrE7JvxgHhp35w4ooLNfao6uBTd42Te76MTXC2hnS8il9uSIFKOItRzV
zsq0rOJDuIyj8ivW2uMm4sToxyxIsTEq+yYs+8GZW2jOiXNlZCNrh6iMNHROYH9p7XGU47ILKmvr
FUlMMDC4OlS1cBB25IjanKb3B7StyEsZSZdDMwk6TiX7UyG2oBKoYyZn2G+A/0E6cICkFTBaSeJN
YgRItosvoMP2Qgsz8cda8WibFqbKTY5+5R6S+/yDbavN5XHPunfNJSss3LD1eFWmHfpH+e3FoaSR
VZ8/jT3sXsxSrgR7gyPhOdtrlmTt8inOQv2iqNzcXQOBQ+AfwB5v+swDDHe+CowmoIER/3bxBDfd
HT0gLjztfBExD2flaP+GcUGNudfX75atsXaACr+97+Ithiu2bvimq5h0zWCO4rHLugOuKkHjovah
9uA9Ozdh7WBRygrTy1pQfmBNJyZ9Lhc5ins/yzU3TdISQyiw/4pL5HC2Vlm/ueToTxsSU/JZJsaK
+rf4mtPCqdJE3MCK3+h3gXTlKGHJ7dtT9UtUNhgWcmOQ00xiT911x7iQF/vscropGZgMMtx6MXoO
fjFAXGH+kRFtutGXI8h0HdxZZCHnKotyDX6nqufPIxPElDFnxLCfWSAIMHOZpH+wiCVyoTBlUF7h
z6M5AbFVq+WGVInJgXTxRemMyjM74mBzSJp/SAekiRH3f5mUIKU6X3q0xkJXr5BUowNLqMJ2Lg1a
rvIbH610CebFC2/YzTwxHoosCpCX1K9R3iu9H0l4GnXHeAfPa+Wgn+tCi/xQYlZFKxKYbk19bahY
aQIq9c5JRTCbCAX/HN58Zda2eWnX7v9jTNOGVvk//SwZXuLyU10zTIGerOrF25mJtpI9i30EtRPi
k9jUNLdXNd4KNuS3eCADHTSBbMSlSAGt4DoAEnxoJVC9dZTAdl0wSFWneprwiD23KsPxCCeG0Klr
93Oz+BiREk0YV1vshA0Q2N4CerhG/qsz4slLons05Uh1qvmUho30TOwrPXnmVEjRmJMoOv0zwvhh
2gccRKjiZg7Nqk41MkJN0CZLvqzyIUU/+88d7TbMGL9NsZFxgT+OmIISfJ+7ltGtJHOjwX587GLj
TYJm6n6I8q63RQ9VG0j73pC4uinz4C+0aKph1T5eQ7nkbGMfwa0kgb5wIEEIzBFZeKisNYD73URz
v211r5XbN6BRB3URU5mQUTyRaPKt77J3yU6vwuOIab7WJ/aEEP8katR6mPW+0SGIh4iWNqJOUI0m
bgL8i4Fpx7CJ9PtJR1sIUDPlT5aYjaa4JSgsyR1WWMBiF28NS18+BVYpHZ6Mh0zF1XK7gn70z63a
SfzYcCvSCM19xIwHMSPhB/H78W0FNXSgcgZqZJJSqEP7nf2dwkKZBlX2aMNc7cRdK4ci2W58m/pm
vrlkjgl1j5G2KVVRlkLIcfJYuk0yxLGbQWL5645vAtjKiS4kbAzfNodk+K5QufOafSA9nE6rBJ7m
3Vvu+ECEjqrf6IY9Yzx/ZVsaS/Ay/ptK0jYliFO3MWyKdBmBm46yoTT3VvhzQkSB5SgKEeFOhjLo
Fvr24qc+PEq1AVtsmNa7cpMrXaClZg1czwXe5CzAd+/J/Ny3RPr+DSbgjNif66+sAOC57skLJcm8
nYQSNqNEkA71AawDBLQXyFu9sJo/y7oNExY8cI4zY2m4GTreq7rIrLjwzq0c5R7nrIjw7L49w4DG
KP35jS08vn7M+4aCbBbrJkG8en33YAq6zhW7T5ZwfC+UT/gYTLVlzuhNQ6ptADK2khIZk7ea1Dt6
+QmJxSP5rVJTmT0qnsIjnC1PusRveE9VC0z17AePQEynGrrQcHSU8hQSZOz4Gta5j5giYlwDdb+X
q4bS74aVQIcfhH6fL8CpZlmLD0sdnSs9baXYBefRu54OcctvWeuGKSxLhdI5erHIAjf0Rsj7RRPv
9hG8m8Ei6vl/CBliYlGt4LbVKeKuVCMNSNgvYZFvzKQzeB3oJR+16LJudnVDNihozk4IqwebIaWZ
nv0jTvGTt9LtWQHMGocpz6zp3/BPneEnduQMSCCZP/nlHUzCXKCOEzncOaxPB3mdCNS4WjTNIQ6l
xnKsuqdXjgOSoTvLYf0NdSDfSHRiGjhk2kqvQDLqhmXNVygxt+YvhcyCwlHakJaEUeqw9oYGrRae
AiXgJ7rDa9mTiw57d8WhWYgxOowLNTblBhQs38iZqh5zV/m/aTNICbLSd73NtT944rC1z4nfLJ6I
+fdObhvz67UuNK5qk+ju3o6E6zCl17msn61FiSJv34O/xHbzv15aQrQ1rnGiNM90qZRX0pJht4z6
jVrnyprOkv9xJOVXsJ/A8lIRSPFdlGD10rj24AlFc6nVV0j3x6DKE6jopyXnq6waw+6WVDp2+Fvp
hXYVHZqAmhlZX3Lwi81buNnpKHrRFZmWrbLOhZMNcmmKrz2osWxfTCu6b/GU6ysayDpxNdVrbbpD
+QREDs6pr/r82rsLIbgtqNWsLFH7JOcquj+sLHOlcEnxHCrZFs3PC1vm35lEwzHptbBhb+MaUrDo
zAtNKPkxrYO/8f9XPFqduTblfaAkrc6rLxqEIJ108qOxUAZ2Cs+DVEH67J++tZS18/U7LfwHW+2t
+I36VEitT8QuHGxcorV6WUcfNHF73/JSGOnsVQHuZedobM6422444zV0eGuYiXSyCkIjf6WQ8VBS
UzR9AVDcWmrfWx355obN9DcD6qtHSc/iPWgJ9zD5QRLnu2pYAiFFFOS9e4Dt1OmwN45HYxVPI2Zc
6g7XaUIuVB0xbM8qHEgzNPC2Jc41YuXC80ZDENybLT8zN18mTFrj1loy/jYq1azTc36qreO4jV8t
Eq3nsY/NDiZ5P/bcCAFmPTHo6kzWksG4z4EHz5Nzw9wTcz9pWxR6pr4bOCdQ1w0rOTVvlurvdzX2
CfAeLE2bW7DJdyRaRmywOECxeNW7S43qWGzs06L631l5YK2ATq4bNqOLjHOCxFNr+Q0u7GXRvoz0
fMSOmuKEz7i3Ou4OKfN6U5dKcSdjkY46E0rMdby7Mb6E+C38k7lClv3ldyfKh/W37ln6AgjnqnV/
Cr0gcCM8fiXZx27z0R4wSs4ev+mfR8JWg2syBwrykVXGPQ7MyAswOYmAKWUebvkWmaPv6Dhn8Pbj
72Rt0yz42L7qa1SL/v5UaX5QQPN2NESak6pzs7sCFOY7/iouDj9+kMXqG4/vDLop8x95Y7vkv5Rf
ySdEEsalgod1TjIPKabuS95yvX0QhwNlTspYUHoPc8m/SnlPAr7bOxpkakwfazIzHy30ZWjOXYG6
h+rUfmC8fVOAc9su+m80xkKue6VTmc9ilYzBhExYSnRHBqKUQ62BD7+Ntentu2m3eOX3FWk6uSpa
rx8FSvIHJQtm/fCE7HkpaT0GhzDzppUZziAeOSS441x9axgeZY9T7z+D3SdvpQTnC7AKCT7s4bsN
08jY7pn/AzLhe9aaK0tln9G1eIF6C9EDyQCZZElcXDsF+nOY7DCuDxA4YdySuCmLM+Unucos+ren
CoHQFzPpkjBMJmZS6QDApdhi1bl5nvX3phe1TEVdyucjaMB+SFBMlLaoXttDdigUv++uZ/OgL1W4
/BmH3zoA28QoxB1Un2LJKxYZCE+GQhqclYSEVNPL8GzsIYh/SbgIsrvNHta3ygMTIngEzimpp0WT
c1QM/aZJoxAIbZ/nkCqz8ZP15JrIL3n8UI6y2VcYMEXdyhQfzKANlOmUyeDLmyISlj5JWg4x8Rbt
Ug5jqlW1ECvdOTmZRHJsvowfWO78JMmX7Tqw3PefzjEIrbLqJpK4tVtD13cFiQD670DZoUluP+BM
ZWOpjeoJfMl6gDnklAqQnH9STCf+2lKlAMM+TxyafCjGCoY+afmIUszflSxPYvya+A+tUFU07jwe
yFMv1KMQ8+ON1T7ZT6qb4mRPl16rxP/lpllTRGbdpiKEL2B4XOKmT2cLBCzOt9cKBMMji3kOyLBF
hSdUAdcNSWh8xhnbyeU+m6J2S3+gKsuCj3D9D4sJbbMIEsxoEBE6jjAs5NTXquFy5u60fBQtpefb
pCk69TlJMzBucxGNBtcCd6qu+kx9+PpPtKD+r37MB8YO9Ywl1bKm3E8MMWGzJaAKPUYc0OUjuYrx
wgNZwc568xJHcMlaDqNk1X7eQJ7MLQeL6zdzGa6k2g6qf4xZAvDgHUB0tpHDuAz/z9GNIGNbhZgM
4P/Br2XQVEwnhpUYIWbGntlqMzKvg7iZBSqQU3vQDC825DlScl4QcMoGLQx6yxU3zSkvs8W1qfd3
HxkQHqJHCFe/xLkxxCf312fl02B0I3/99v065Tt8H9f0Msd99GfUIcAKOTnkg1W7Dyc4WVApXL+5
W5baT1j/BkK3yvJXJ+nMZ4QOmCKDrWkEGZRwnyLVEPMfk15U/irnn6r4rFWXZ+nWRPaWjslH3FgD
a6BmHbZjkEV+X7AloXVWiqNdG20+OfCazPBH97YPghfeV/33fRayJHtWtLnIYqQVFfSEKa0eALVJ
wVL4562xknGPQhPPb7xxhmR4moIpFeEXqLFqdCdxOa5mKAfPnR+h4G2bzk6oy4soBf5qG8YADC6w
PFlvO8JivTq0sWtkwX2egA/1l4gtTzute9h7Dj80M0BftxHfdRMwoQLLTplNB5ZbEZqYd+Gx0PP2
eRUL49UFRl6yQpAwZStErIWezGNkswLa7vEIO4dbsoX1/KmsWfPOK+3UiPoFbWjvrTGW5j3irjrd
YkO/nTD6U8QaTlfe9QjRI7tGT66YYEvo59rF0DantPDqMaFdJ7W/WlFEyYQISN7MZCob0MDUYiM+
CoFZ8pTna3mFAaauMvTC63AuwN4591e3Eqzdc+9ZGrXWCxiMGBDe+E0HN0jNlgngHYj5HKBJBk72
9E752WXz5PMi3k3LYuknXO6G+gTZIibnr696bpqzm7JCyIJ/qOyZ4GSpHtyKlUF5k11jt+6XY0HG
PhJLHmXjHFNad8LP7jOFkNT4UJDX80sMcoYs36cDz0zhbqyUJXcw3gjyyXvkydtJ3t6SyD0SWECp
yyFBzYMkzUqB5r8xLy2/23DU77fE9nNmo9tg3CJN/eWFdI0ppuS4skh7cZCIvFkWqvGu4LwoUWfh
F7uOdP1Uyg/K61blRf2mC06nRIsnElm8rBJMPyRry8eaONXS5YYi0+Zm3B+vkLHm9Bwqf+WuOLtj
OqhPwSbd3gwzAifsgrUL+k6M7tD8uXD2pjwqgXPsQ7fPrDci2reECxsCiNOYNcVopPK2Qa9xogrI
P5x80Hmjq4PI46NLr/c8S3HPpUMnesJDE7uKFsyq0A+cjyz/CcnGx8J7I4em9PAl3JxnmPqnJPA7
J+gLv9MJ/rsdNuzSbuLA2XVNDfT2+WZOIOfNACtGf+aT8XLd1JiEXCUp7B8o3B/vdGixzcLxOnUN
oOpyP4f7tBxr5t6mRjkbVXKxVsbh95hVhmStz35skQBdnJOBAbJ9hoPqwsMU3dDJn5vsdMPLB4a1
59o7Ug/LnF3Up287wGb3/b4CiCOluvUf8cwc4U3aFzMVni1dWNikQqXcZ/vS+C+hkPfvIRjds8kF
x804Sya3k3i86FNDdM3kJMSXHc7zTAeHOzWwrMoS/mkxQs0Kbr+bflTmzTqmOSMtvGez9mQJoEwN
f1MvgAWBArwHSpGQ8VmHW+I/gW16SVSlBbDtw4JpQgZ5VNSYdwwZuK56GttKmWgPbU39ZHOl4Uyt
6DDt04thflp1VTSJ0+6pDlWaIAdRUhWtAmN+x+WFU5ft4oEJsQwpbZXslZWaNsWyQsShd89PSpqP
dfwrUVS+LKZQ3GNIUkWf5GVcBBhMzOmMFaICMoj4lhp6vBfXYfx2/2XifrnX5LLSh6Y/Qgky7lKF
ymKZ5RUxXKV8N0ASW86aHdnLkHmuAwrdO6kXXOzuaBMjR/EWb/p2zYExRGH+plxsTeR5QJyl04Ev
Z9sPrRvha3A5oZx2uolUr+yNKRxs2wy235EUcD7RlMqEz3M2z7j5XyT+Pj8EhdbgjLo4mrNj9VuS
eq6Nz0nywcwZ83rrm4EGT6AeouAirNN1YhWzm0b+LVMdsxd0flFFW7xxISJvKFMH6jGUDV2MDY+0
fUSn3rheFXOBwNbryjbMVO2DP+bT0OSlBGXDOuYmPOWfjACUEWzVl+BfOJMIVPEGMoh6baO75z5a
pGFKdVwes3Ovshkd7CjWGHPz9shEO7jQFxG22u0qRCcXfdfY6J493kXe4gyh7JUN6ESORuoVi6Zw
OkaEbO/a/KN+hWKecxpX7qkwBlAj3K68CrHGvQBjWU5/110tfeBtpsiQ3SO6OrTChb44+SFGd16o
2aIccy1F5caSeaNjGRF2tWExOGVcVQLhId4rlfqlKpTvatGFxGTPzIikmdBZVfawJYSyu/UBkc1C
5KNR/YyxGG9Rw07WuOZ2MpxZF0i6QTSo5f9TG78KtrvpqrawJ3hI31To1l1ScJDaxbZIXC0n4Ie2
P6DoLgXt3Di+oj8vXD7G5GIml36Kij7VGXcM9aE2W90L5Lcvonc7Gy6MhfciLjAmkMWnc8F0Cwg7
ZGB25I9gsJ+VIeAFHel9HakFHkeChl9MFVjC6jG/QS6JjBPa1AGCdrAvfAYPqduGpVmAqWpgRn8b
u6aXvx3SPXx4+kTNyCRHTT2aatesaSPSV09QAqUgap3ofH6kLn1H7bYrlrf5gfP4yHSzQc5HHbPC
mSfena1Vx3yLgjtnSgsVykTmWUmkEtRz41dIymL59mUjw+TDa9GaK9hddtGLDVrxsGGa/xN/Ir9N
7JV0lHakE82KvduCz5iP5/E5QgofU0f63tH1bOK+kSgJ3y/eTX6hPZwvUOwRKNhk6pw9f6E9cYLO
PFDnyJBaG7KsT+SpWi6G+o7rUHUk18hq1iyQMvyflFfbXS1/oMGgfA7p5bs0fyUpJux4PwV3AYc5
2olp56Xdh69aMvzp9PaBTbydzOfW2B0/hPKZyK9syBFQ4zWHDfLxc9WYp/srWznuCyZpoPNIP7RS
pLEuYF3KiuxyJueGncF44hgYNtTWm9PSM02M6oUqhcM+JuxmpuUX1qZlZQkWSN8mX7pyYpevAQWh
IdoHCJp5aSHbGw7MJDPVsjrhtmYI2k0/ZQwBn/rhwLhVx3+HPI3W9EARg58xOKuIwydf7RIumGKM
OwfI7XuKxQl+kNB5ssbnIgJ1xr+XyAQUzYZnR6eFFxSbYw5rJobBcTROgS3U1ZskJt9vPiQfThDO
c5P96ZrLOZBaH1VzXDIm7GR56/twjwJHqJtORDMzMkb3cLvqULP4k7fSrcnj43aY5ptoWKVKxY7M
1fG6XMbjXh7yCYnV06AgDqGtiXkAn73rK+ZTOGjYRsIAmCt7yUxlr41qg1jaFfhnQOXnYgGpvtrq
XYybTEFALRrP8fzHQ7wBRMCscCrK01W1y4mWn7FIMvrqb75lTpq2hGnaYQ19sK0RWnB1Lnr14oAq
fni5gcsVSHOboCOhMLJEriG6sbdXQd6/zI/H5UsqatzKoYh2bOCptQ29pdCY7Fe0aTsp4+2GQ3OS
6xwEcdP0bxiKxPnqDYtrkUQNnKE7NuR2zapzqrxqM2U99Dy1XGCXyHAjY0RkAIMYQJwMizB6Devy
jDjCafpBanAN/VZcvgKM0wcGkVq8LbxmxK7hpGYK0uf6SrfR+NRuoAprHUjM1ix4Vhmp2yguvHoX
eX7qFY5L6j+uOb4noLEryuuLqHzLhCJ2d2Fe3VWeYb+WHzOrwuKtV4xhJbvsyi6md/NqhnE2bO8l
Btf8IJyYp9VOUslGmjoZk07aQ7kgZyopoRvYnnOOAGjMc730qFC8PHO4hbFNJAJCghfrZyT/xBOf
OMvEuUcO3sBjGV0W7oIof5KUHR77kUJlPOmpXQFReYN702c53u5L4J4UF3QJ8sx1MK30BbpUo6XX
xt94FD9nTzbUb7Sdyi78t2F6XBagS+6Z2SP8mpSlQiuBGytMzhudJR25TRSX5Gg2emy4NbBmhfBm
oTDag7hLpDBqHot5J6kwV5RgqOvdFRMUSDsnu7GyNgEaFpsES8ytfJpkKK3y44EXWZ2B4djbtQdr
JEREI4hmbIDIDnSYTl/Au2A+6rjIQ8ITRsc2r68snWOaJFVyq5v8JUUDRuexG7kXwBUO25fqr4GW
lu9J4vE8mqpBOJZvAdQebfYp2Eoua14h57qYZDeua9DFeIk4MGfrtLfurbAz+WjLknx1q3dyShEa
aaj+dBezFmd+GXzNLFBoSbr8SBqwFhcf54UWn5Odvko5ddwklzITHTPGQAZlgxDAq07uUVAS58Q5
+KFxOxXcoUgcyTadB85qjqDRlmmUV80fhkFzWIWP+Dob7BGWeg9lu5vOEVIaGgMfF+VFJLGHg3Zq
CXeSHMYwz4/2M4gEeEm7JvIiB7+8qhsRa3JJHqeeNpT3qr/hwysOBJh4OBoyvYYjTA4lkEhfNshO
/RDJvlXgHn2bZaHubLn33AQrGz3HGGJmbDbQqrbSgOf1T7esXIrweuV/eNLxgWqRmYfAWU2CxUqZ
YX1+E5f1xxjelMSbXIRc98s7XfAlziXbb2p6EuOuBjn48yK3DvEg20uwQb7zjLT0zcla/O4D9UM1
lMJsWwA6s7NSpU/0CV9AxjZf2pc17maMbTZzHHOTkkz0NmU8jA8Xu8KV+ItPnKmGu/Q4jEMTTK4p
LeQjcNyoyz1L6RRH4JZ+uSJfuNfHkY4FTebTnithNbiziTClBYRO9V9V+nSXyT3yntq3IllWLPQT
XQuDK22zEUgqn7eOrDTRmMA9CJxWSymfL1eQXEKjiLqzD32xoNH1JIR2iAr+TobsPqBUr/SboCEx
DBQpDW57SWfZyv29ZaQt/Xs83ddUK040o0m715BaCyLZrxQYmJPLBxzmF3n4eIY2pHPDVP8VhcUm
F/3cdjkKMg6Y0soN1UDKl4TdzgMigMgFA+2sxKudoOE8QSUWtLlklQJMtooRt6sRrZGHKNtE6t9C
p6X2BJa5SZMQwMaclXHuq7onNCFjIBGPgo0d8s4oycgObNz6hIIyE8iQ46EwsXpWKwJABK+EP9Ok
JtYYCpg6/aoaznhQSpEGzjr9w2MBINOs+R8mezcTU71S1OZV/gqnKxt7D5bkLUEMEBkCV1Fe28zz
yTAWfOW/P5AG48S2SyD1tOZQp/0PlN/TWtYJmM5VqqnFkgFRhmzVw3Q7lR+NFMH35UIH9/0wyLnM
zUqmpB/8ULLA1NQGcpjQSZIbb2bpnaYypSk7jw9G80nMprTaSTKWSe46uw31sUUAXgGB7Zr+LHCy
3E2X/WFMwT4NahHMl44T1lfEx/T2n6eMqqHmBuVpyFxEJXCluj/USBbWQcFUDqn/FvfNPiICkX9x
Zf2qfRqR9uX933i4PC0ssNH/NDV5nPDC1oa9kiqgnlqOBNt9IJo5NNHiCNaUid3uLSGDbSDb+b70
RoD2OR1PK8EPjJMbDdQEJiEFrhUU6F9G9i4DmGcqPWGaMqgl/XT3K2kk+dcu54xXzBtoQWlfstEF
UvrXWYvUsjZVAF9iCr1US1Vke+Lvs4Fui+QtMNIDp71qrCMyyYls/+3WLvPGre3kXO7VdR49bnGy
NUY/Gjzet1EvWd6oObp9o1c7vT7y2IRbr0F5F4sSJd2N1/XGZ5HUG8je1W8gZ01z7r1XNc7yKT1x
M8sdv+eAfXKFSF1ZOjMB3rBBMVCDBAy3ELuXbi+bX1SuGfWTUoj3s96akzb2+28gZvz7L/OHbX51
A//bDXw3jCi+xgPNtmast/bI20+4X7k5j+z0UHAuqtVX6F3gX+KchcqzOqW3tivmKzP+sXowKkM1
3aZcq/4MFwoEuyKvp5Ky028cC6TzAlLbAiG1fjDvd/UIdpc9Y3qY/6uLA46nCeMc7E9K8iLT3dMG
lsozquannMUM44I+Cmx1TTJb++E2xzB0HvIl2Z7c1z5ikU1SguqE1U0cExu+IA4Tof+YmLXxGJ6O
vbrRVXfNfDqgqzibnoU8uOuO1TylXh2kANYRVTskPm2xAVyGqodoqUaNo5RrpQCtz6FSdBXaamGX
flJWiNCtQmrs0ZjKvJovTrP3Gj/86TQMUjgVPsWbvc/hBfCHW1TqA+Y1hcNfsWmglnWqMsEIF5X4
9bqaeRf0bQojwI0vxcu2FoiAiadxgDglhdBEzURAVvflyNzFp60bItU++kGPXQrfVR8v2XGaUPLn
ZhVfVjdF8ObqTiTZNfYem1qPwq1v/H7U/8OKgzLbi0tQIVpqgzP+4q5I1CkeEJ+IHuGeePxqkMYP
zXyNaRLKjtYVOvqyiMmRMQdinjbAmzehMIZBjLzaVk6osENBA1hD2iUd0KbM/wjM+hL/pzLo3lUR
llWocqjzO0OBsBRJzM0AuAuBrdBtKlomWKqeKudTD7qY9DQQwQ9zCYaJNvcSD5G1J2fRuRPvhC05
6s6CqraVKzA0xVva1P2RQtjclxegRV0dIXZ0E9bb7RsL+NR+jf1qW/W+y0d4t+ZCul4/+pMAJsNv
QeU+hCokYh3hkt1e0/4/kPiZXvrR/ZtHYinLtgMj4wA9llpCB+QsbiIHY6XZstnRB2Xd1KaHtSzE
UGxXicNN88bIobjio+GjFJVhKP8oB4Z0p/p2BtILrcjm+7JHnfjn0V9i/cbOUap3sSnZgWYFnkx4
TRj7pYmIWvvCGHZ+IaYwg93o0/T9i8x1AjCnTxQcZxu9dEuucVVEmMBhRjE+DXwO3L0nPFJhc5GV
OGFuZEOmfB7iinbQDpguknQFwcEU3Z6bJOuFiIm39rpsE7eC/284C2AzLbDxsmDRYMLucT5pxbnS
GZcY1M/VJg19/v/J+J889YSh0b36QefkKwpRwccTd7iGjEgUxUsAtuu42NN0vIMYo6Q3sGSVl7d6
0LfGeecn2WjbEyAof+3JvH2ScUcVYLg3PLKTVLiZYmhnP1ndaDih2jFr4icCsCfJWF8NtjpFGZld
YiI7onpZYX8FNgGUXZoqkL+RXwUAe+fD5ARNaPXb/zEDGPNhPctDiIQAQcrlM8mKH0KGLDuNAJW+
KG26Hhyo6ox0mLPMJn3u97ZtX7Fdx5Vf4JbpxUu1eyB0NLX3bnc2zgb6iQUIMT/4JxoyRA70qJFU
NRY1h6NORyKMO8Du/jZZg6NBNR9HqXvzC5J1oNOOEsTnO+j0Vbq9CLnXULdxLO/y4KM9qWseVWMY
IQkIGr+mHkgj8yF6EutHSuhkx0GVpbHbSk9YRtG29Y40UJmf7X+pa3ZvIrsQEKXb7ZZND2Ve27uV
aCzH0k2scybkKlecqxDD/inzRDDHkScEK46wDc3n7/9aGWUykDvMSSAJKWOFA7yZdQaEUg2iukll
+rZc9B/TNED+/qVF6aO3fa2yXe7xkUBt6QHpk612mt27QR0nwLqVZzVSL9jDNzEGHCLYADTZPATs
xseI4XxkzH0p2p0MleCqRVzEjOUJp+uTPinS53rNLlnUfEuRSPIymWSv/TR6e+VXEhDg8BOm3MkP
PyLLmNL09Wdxg03GJI7WjOqWW/e2SksU+wAipcTdXoZFe6f6xxbPzi/ddJbRbhY7ITLyoxzj6KWS
BOYypUH8luwySE+qP8STSoWC9/VRhhWoMmIf+Xz6WskMB/Z3khRGibMOWPHbbJxvfOonTTYXI7BO
iPw6DYl0gWgE0y0hEQmnKBSqtk8WjVgXGjO6Pcu0VqcbcVotB0zCeKdy/UILChEjPjDAfl2WyVN/
akWlDlfRIrI0jNtqx5y9+Z1YCIZd2lSl8yFXlQ/0eEPL0RPLyq90mzMlK9YxUy8C7Tnca9OuWl4v
iQARQ0bR4DqxDkoJa0GOAys63m0exvObgEvcvmIdGDH6yg1WJxIl4ioLrYZKLy9+JW/KU16xXYjz
K1+xcjmGoTAPBmTS+OQZKgcJF/tMtR3GD9wSwWKYvtDLL/nlq4krMD7zuJ3l7SQpm3vvv3F/t2ro
/cWQpOeBMJxFBniqGfIZ6WcC2Xd2JTMjjadvLNb5+1rS0r5KkAXRQimEtH+DUnoiBKOMUo5LEmCB
nox3xqDeWuoNwnY7hAVBDce9g3Wl4s9F95kqBmPDscALGfvRoWXedv7OaQy+jesMPWiLRaoZFYNM
ERTT3LfyIqlBzI5ITYjYudNZvR/bJ7cGsYxTPsRQWT9VkyE3zQMqtJoessugC/AcPdWjeZa00uDe
YgeFw2xXpC7GASsYLZv/tat6qwbSdRq1jFwsPJkKyWLDSN7DYhZv+jgjUif6xhTvS/XOFY3+FCQE
RrqDYY56jSjFO8aYqgssNtZ2/9AvHPym1u991wy4WNlq66ttLhPQWZtkvM3vcVmgggtg9ljgQgPL
XcKlpXyTLAviDTInYqunBEMs9nK2uPTKJDjTxyPqMUNBckcfgfWTmC0KH0MMncv3QvN2Hvd7dSrl
VZ4ycCfbaza+JoJ/ckK6IcwRWjMJKKyXo43SaorYwd9eKALrkAIeDm/OXaXB6+udDfivMDhNON9H
7OhHyTB3PL1FuhdHWVZwAW0cl/EseVbQVo8uW8opBAqCc6K/Bm89N++PWml3jyKLjI6W1Lp8tFU3
OGqMm5nGhp99Grc8PQ/mBi2FhnLxdJUYV5K/kGx7ckRA7/XhVEMxnRsF7qhdpvNEWSQQi7TxbFRu
LHTTRqlljSU/cszzY5NLrCu7di30nUqlOoqQMbb6WCA3R4v1g2cvM+M+KIbwnloNcuryN6yNprki
URkI5sXO9yT89XovIPBdjy/St6tICbgLPEZ/oPQ8BsH9vHYzThvy6/8I7p4bY9sP/O1iVm5wQRR3
mPva7Rjni+L1iP6ENsJpR3mS5nkJ7+mfz+m2Jc2vLIWuR54r7+88A2f3lklhxMWde5DGjMhwxcig
TrJ8jWVgVCCDGwrbF2l2zr5ictakJw5hniMjoH3YBOhVhToqomqpT2+llY+VmshuFLjGRWdkfgS8
tNik8Xd7NdAIhjRJoqoEe8bttLQTz+jzlbUmUyOWS8PKCfRwLEA0TznxnRk631rZeMJeqxT3JOJ8
SgXfGFwL0/ZWGthj0NmxAZ8W24I8GRmxzLdFQa39q2lwhDSg/Jf3WQmbpsqis+nbLRVGktxAmU2O
XxFX48v/jplPGEWGSlHxGag+p+NbJ5ahKD0QxoylWSFelRjjX/yLwzcWBHYHdD0MkjPwbiAC76iR
AaCb5cHmaOkf6/1tgXaPW9Ovu6lHCWf17tzI1ekvjN7eD2LisULQveBB6fnfIXr4uwJIsTF37k59
xnvqN7eCgMrBGnZCaZwMJ545grMkvKAGmOXX0zDdW/l5aTnCLXzdoV0iqQcG1Gg5Oze6c4MxoZZm
xpx20r4vktIP/GoMMkAK3CIv+jw4bEnNOFFY6thlCPbgj37gTwT3Y5l7K+qtHPNaSUbmNnur2Qzo
Cz3JOgVhc/53P8C6A+9n7UpT4zT6xBphUONV4qXs99S1ynz6ZWm8OS2BdsMBBh5KFr/2fa2GT6ws
AOIbCiJSdAA3lkyKkLm50pR3WlmH8bZW4mUubS14RcEaBRN0acPG+YvF/Ju7hrLF1bVaoMtihIp2
FPCyCprJDJr9jRQLcjm1eChS46Ooes04mD+HuI5Mvkq6RFNeut3Yzl013vbwb5SOnQndZLsZ27dQ
RvvfvJpzxrlOEyvN7wQzg5PGhcE6HGpOV29c96pwirxlo8wcLa8vcHMqo2IdSMjO5yGkC2WggRC5
plbBbzLlykx9Ak7KAJemmEyo6+pFDm3+OVynDz00Jt0ma75JFlOET9AevJORotaMxL7XOy4D4TRW
9lo73T7MDYQmAVeYqHbd6xXvUcj1Low/behoJ6vLhlhswUkkGrPASDPE4ks8PtIoSSkiYE9lngnb
vyEO19VUEvsZYjwgmR3kOQSql3680qbDNGMYayTm3nWAnh/5FS0MMCX7OcCcaq8bVc7JLLtkEU4r
A/lj7BfSh6n5yO4/WFqnSwkb4xc/0ysb13facTi0zjPSA8cVEuZryvZSlCgEjJkeozLfcL6edett
02yMKGeQ/aAlwy/SD1+b3ajbvngm0lqoab5ehPW6rRaopiKRW9jeJAu8y8TEtbQFgivMekM2yB+8
dtBOWSsLiSfsOxGx7+wT/8FwraKEkK9uMhiINImDtQOQ+GYT7MY5B/R/kX+dun2Exohrwz3p9NZ3
+Pg8G3ajSPrSlmfzzFF6QigoUaRQjmnA65gLroYaS2umFM+SnHFHgo7x87fBS79U/uQ4JO0PyC6D
9LiXWCDXFBoVifRJNaFXtBn5geflSX1CQvPDu/1GuZQsO+IT89Y7hJO3UdN1C+HR8g05EeVOHCjU
xfSHtW19fxaf2jzR98h1xJNKBWZIkS1Lh+EM0mU/Dz65v0NT8dAcPWi1bh5W9ialKFXRFfvRHjJT
8vNA3FIgw6sEo877gekqlsSd+d3Aeez/tTPCAu3jC1xeMYg3kEBmDnX4LPv3bJkRvGGHtT2Idtjc
JJdeJ3tSlmvZx4gDAeZ2NM13Rl3sLslq5bKrOdYs4PhE9HWEF6IJc3qAAuybIq7cu+Rhi9R7VkDd
a3KMQQxSUTXWx7i7W7xlSlZRVTOb5W4CurwNHQHfhLfqQsFDbbtyhW4SDKaLWXSvSpcrM/GOdT4M
JMJO4awI309eI8JwATYQp09la9nT0kR8qpL7nUp8ZokeLS5wpbST8NheWID6GKBqhlZRKqjZO+fX
w033Q2eZRL85GPJkGSXsP4Qo2YNDfLP0ViUfR7QfdM/QADhFMttY3zuqGo3R/svaBMoF6N7+y/90
lMLKPbgVIf7lnRrfPi6EJBZronWTffm7eICdOwzQDgt5EHYiSArEE/edp8F1HHG8+WOTvTMCCEzh
BIlwRwtdNEaqKv+d5ZSLw68q5apI6UfrrBZPxD9iTHm1PgsFyt68VC6oeh4s1siss6bOGnOwwNJj
mK4UBjLFXWdrwKbOPMx7kv8oGK26pjb9TCicUnUGBN/rxZdn5vMHpiy6bcaRuXHmEokfP770ElOA
ETqkuFHcejnPFjK06k5ymnoReJryUc9JrqLX5ahAmwVpe5Bl+KtjJuJfvOqHnEaTA3I0WR8foj4l
Sk92zdJMtD7QXw61i21u9xxXgsGR2jEn1luNPaR74jD3APbCODqvUzYuZ2yRowOpJNWr0EbVG1xk
p/AXnUmuO7fbayN4JrSXM5162wceAngOQMFQdc8gc8PeyqweZVuQWmxw+LFoFQOHKSrAOVaTS3q0
JnGUthw4Lc4nxCEcryIj9ln+fZw8GYZ9IzpQawUk2CIQQPCbVhz41Mw2Z2Drw11p5Ek95ZILSOkJ
k35hnxjfGCPse3HldPy/roMwkTZxV1yTW/YxnIxDNhRg//eSHmPuI4rPbPP38ld2ha2MEiy3Z62O
0C7qFTg/hUGmOeClD0ElcAWHpW/+aGa0CJOgLVFHv5mneO0pVDxAlr64i89zulSzw3Lv1S5SEy2M
n30Q3rnLazefdV8LyYTuduw9X+4IQ+g7B25VB10N/SmK1fSPpDlV68xSJOsAY/uMfLYk8z88IuH3
PPnw5Ertmn+UHX0pmQHB6d6IdjExDHR8eZiHEdQNtaHnCEOFsgO45ku/CXFhDNDAHtA+fDv4xRL7
psXqbmxG/EkJ2MFSBCspMqPnxWr3CoqmafQ70zhO113/u+KiAKXNO/PwHKWgGBf08iKIAnXPpgUX
oPoZ4S544fYTcN3dwrgOwCopjUlmfuc6lp2R0OQTUui1I2b4lkhFHUItFh53WCuYuXogzHG2DI/G
1b1KjyiaYn3oHMN3tWv35S0e8tU/6Wg4kGNA1h4r9E7+s6YO5XVt3dafGZJfNC0ed+N2Me4/q861
7WUCLc/1OWP4OXP7OysIx4XcxBSz+rQnrR+wxavHp62aqjFbamNLrKEaPIkChfxbTbUFG5nly/DV
V158gLXiB517AjW/V3PVQstiQrWrLzZrbK1vLD0VE1gluXEAbJP3qbf/ztXWBylrf4Jj4a5Z0/UE
onOMwTkkEzpc2w9u1XitAQ6acZUGPBTh3/v9AfIavz5u8eia/uCRh7rfo1qM4oa/Eucvyp90t/f5
NlwnoUUqI4Ri3tmFa8PJ/KZ8rG1iGwBKLINKvaUBTNU5oQKGLJhLiv5EikTgy/x74un6HCxQJeoB
aJe3eJNQ102Vn+cWXV5eMYTgmbx/A2LTUUXqLC+k9m31Ii9DqTi3+WbaC5wIsRCgsLrEiudWRhZX
kgBAAgWgYCuKylOxVUEqZ62a3Dh55n0hFtlywucX0fouNjcQzITb5JFvS8RB6elz4/feR1tQkjhA
EmLbQsggW5CObyhnzWsPAzL6oWmP5ouOFWE8bgLSiTg3JuAuIRbgs4HJ9RIvzEXgw9lk2p0HcYAT
8InROtYvY1qUhyQyq7qmf2KlTJRJRIR39yJUYNcf+LCeFWmhAJqGMOxaTFL/EyAW/6FH/556dxeQ
l4FIs3su5V/QTGl0Ugy9DniwnnvOu70fWT7Laz3VD07OyD4YSTPSBmmI5d/RYPzPvBIoZ35+Bw2z
sPU87U08QpKG2GTizhGFE0pg6VrMEG8iBTfKgdtYun6FJL6X32+XaLNDOzmQRJswQIFxmzlUyFSu
ZQiAf+Nt1LFuT+bPJkT04aJxrPHsay4QCn5VPq1ls3/wdI4o8aIy6RO71fZiaoTl2BpSbPFu0u/m
PhT+9NaRdgV08YWIZuRywkZebiwEkhiUYKp/8gvyTV3oAdwtiCzVVrEBLh9qZoVmNRghcDwlfHJV
rBXK1L6dAFwS4uedHzwxSb7ksFsFzEZoodNwAMspsPu3KfVyGc5j9cqJ/F4BKF7Pd0VpdP9HmW/t
KhyyjNTQ2mN6J75eAkI0jRhoYzYxsqAouokGWmV6N1izHXojXMWVYHwEKAoOXJ/kCca7WRao9497
mTggqZS4/iJ+9QyQ933ZCDeFBRe9VY1XbeMNIRMSByFQQx4u5STNw+/2DxXIAGVhvSPEmG/qtRBY
VU28GhFXVUJO/KVl/MABuMkGcxIQv8HBcfmizGBKtlZmkMRAE8uDfKdUZnMUHT8cbi+8MYseaDcp
agqVRpGWagqhOqzgY3yUz0nUK2C7UKLOVfK5E04MAWlP/aszP+cmR6ma9MGO4hyAuLOwvCMFQYE7
QrL8jeFaqsHogdTo0oSY3+NEGyB8LiXIJUYwGaZcJbT8Ge+9nq+8ZmWl4KJV3PmrOqbn9rl/1rUT
3hR6NSW1PKF+bgqkaqqAnLr2my9+ofZdtEP1QHxKbHLoXzRebH5aJ/zruSoOT9FlU7njhh3+CDAf
PYZ+iq+0iSKsKbdjkCpWZY6Ec9MOrSCn/EA4MIDAUlqPXtzhZy+PbwoVB++qoUQcOyM3BjcLfJiZ
/137snZjPK6iNCABv6topB9oU/l/BctnGnUzDBrO04Y8VEuOHmMmz8QZGt/sRyPX7G94BFjdY/LF
o/evk9Akoq+OWjXStqvXf0zEykC7JW8Vnud1tRKBmPwEHUnyrje7U+qOPvvtt59YDDmgC5bAyzM9
EBmdWIlxneq8EMXECGXESowj5g1PIwqvRFljzEJsKQoAVLDW3hqIVRqn8kqZDzWQ8ItKZgwJ6Bby
L95OMqWcyQVe/ulRrYHw/C1p05wzGibDnZBwRMcwKvNQJ9/5Lt/WvwPFLPjhuk8GrsFSp4edo+uv
BUstGTrxsxEroWQogs6LlR49u/f6MwY/Elary6RcVUQJg1UB/c64Ld//lZtmaNzGm4JX1yLDxEQR
+JTC7LiZB4LGme4cAuXd9MNtUmUi7JFhOg5CWGMfuGFN/S+jm41oLCT00QwDj9wlXwEv6NX5OkE3
44yJwV+FOB9yE8G3AazlCUNWhTh6P19klhkdmiJZuQyqxK+KEGXGVpgkFGdsVXCSKuWn+4skKsTc
h31BI5pRkD4eEQcIcPqU5OGE9UntOlPbghZR8+NLc1A/JU31gPHoOXk6mdam5v1ALAPLT27MjDt2
EYUX/CQ66SfMy+rUpmPu20fp1mQO2QUDEQhWPmEldX9ZsAfGomzX0jUDyn/LOI+68tk0weeKtwJJ
p2XNxGdQ4uhNqxmKIsKKyoUQS7P8O//qbzlbn+0awBd34MhcDPC6UT57e0HBF+0l9WhzqynSG4Dv
aUDBJw49/IALOxjaYq0ds+2xsRLapvjGYjdFL9n3BCj+wEt8Px6/T3KCi7yXAqryzG4SfNaWIVH+
YJ5m7mJv3bSkctYqFh79yylcsslOfB6IG528rfWT2Pr06Q2mBIiD6Pm3R5BkjysL8FjNQjqrAXhP
mmEJorH++dD3q7ofU1B58vvl248P2bV0LOrogEDrcpHFI+5idWkLGHqpdyWTxXXcXybE2tt96O8u
pDMJRBpqbbgya8VO2UFP61WJCkpAXVAo4cP+3+SFZJPT0uiU8tK0vMh8qOHrxFMl4tf5TEOBn7WG
fKRubluvKoOmO9x2SfQvkUL152Pp2WVX8QdqaEULlBexaFOD816gOtKryWwkhLSuk6tzrt7HgkGb
GwnDSnMqBs2CG+edciKu8CRfT+9/lFjouyGqwrZqybsETGflTB8Q1ZQacFRqrSg9Q3pQ5yVUxRD3
/RBz9AXEDyPjQOj5V/kmdvxyonqoNnklEJUU8jWKZbS4wsXkxIAICE/CHYigXgXVftAWwFR383lX
wEBRNBfawn9nTFmLMgVvToC5Kml2hbxQxQqEmll+DsJ9ln7XE69wvu2tFZMBZhIC1gJZxr+xwOFe
BUzja2PUIqzRBnk6wabT6CDH2A6oLGHarC05NyhsYDnUoLf9SuOYiYphMajtLHgxFuUT6a+mqs4I
UHM2InX+QERAS0Iq87uDCweyp8KRFwml8iM4Z0rNGMkRPJt8FafMdHjp8Ojh+ibeUlaFVeKDgbV8
jMJU3CKfLg23WmH3uZQLXAnz+WKhMfnSfB2kyp1BQS1ctdDUfeA2OSdr2X7VFEcQ4PP1ABjGOKAp
P68vFD31S5En5IsRp2qY0VanZo745mYzWRFqBaF5vdko7b7s67M9eJ/+fy3QS3cDLmYfaSQhEBLD
kng+ZQcefskwq7jnEHydKZbf1qHhvc+e2KaRP7ufO6bcIGbz9YRaihFWN2zAkZJ7+hveso11KDV/
bWpumvks5PN4vX23mnVEkktIKI5NO3GPdKkp/hfHERLG/KjS5UhZMDZBCvFr+qgwcfeMFTUN8v9z
5Yqkutw/JVJHNmNI1IZoxqLR0OhCirnCudtIZR3BO/YjvYAQ/4LqzILoocyJEuvlsBa913/1Mass
kpxR5omJ+wsNUaXJSGBO7Khs7ArWxMCv6+lvi5t7L3H7PGsCBTKCLmsMy6ZObsU93UdtjswC6ZnI
DPUu31+r971/pL7KIhFr3fKkLrwp+wVSy2sn5ktG+m5CEPqIZ3E3xgOKpYwnBtdbBxmC6ka/Tbzr
REThp+9XwLTvYYLmMpdm4LudvjC7q+o8GgkqHP3sPqKh9DZKrtM9oy0ZBavWU+tS6v44HaEBvW8e
fUyIw40Szq7uq1erDeT7uszDNJIQJw+33VGuww+oDh1FCvDU6CoxdQ0zAkZE0ghVJp1gfYoxF+QV
S9Xd2ouyVFCxZj/d2XwfgrqghGZmDmKjTTU2G4tucI5beMAeV6CQcuZqjaqF1/p1XmCjsqaZBXeL
RPWRDECbWaDgSQB4hY5FGRDpr8uXCcKnry1MJa0ILIFfVAa4gEpeZVlNqzAFjalLpVmk+VdDISxo
2HC16lTRWXlokyM4Y2A5LDq4Qf0/ZfHXP8+qpGBtkjx53G5cGqFgkDAgUOVJn4qzNx3AGRegN1vf
x2sF3QqFGplM4S24CaLMTA5Qf9/FYyX7SY+NQT1QKU/ZM9VZF1VeQL5Yp4QQsaA+f+oTsd2JD019
zC2w66P4wSbY96FevP/pW5MxgJy+eQ9KAGoHK7y0++LL6PWLqdhRKbk8vzeH8xQuoDq8zkY7Y7/p
GrtTZbmgyXAP6q8V/4aZ31uHS5nMrC8ZV3+Jq+5dXIkltP43OatmgslISTuFHbtb7mwx4jf6I8gA
l+qCH2mlUidxmklarI9UKG6D1ovAoiWrG+4ViaaH+20dcv+SgY+y7rVAA+rlwoRYD9O8H0bq3mLo
3FQXHrcP4ZF4GVb6EJfZwJZHTDnsqgSMItVLCkjsmsNVI+2VbK56et1TD5Kw5XU1I231Tx5D4Swl
1GbstKtysjQ/lvSHa/iU38v0uWDe08CeuDyZMbAKIWSQcKBrfQ4QPiv89zMh7Mn8msQESUcgB+9J
ulPq8MjpR+73K0FZih96sB2qjJCVISKE9XCnrEQwhbgaLwGNXVLVYs4+DokiNagtoFZf7R/PR/UQ
jGCtypdiU9j04DfUi3MeyUjyMoEufqLEkxE2gG1VLWjphyy8ACIn6Te0DvKhJOgcgZPFK7DhOIwk
qrDRYhStv1WqUtPeV7+NPIW+1bHRQO5yZuhsTvjGUU6+GcCaH5wwfgzbqO9VmeYNSYhl7le7ZqKN
D7lk7/Yi5u+WpeX8eTT+PoMhNdeK00NLEWsEz+1szZMMTN26ir4K7C80YnPItxYOFfe2CfnVWgfG
/1TMbYO9yc1KhSt3P+7WQSV1uG/FGxhw1i3zqr44a0PgvlpOdkO7UGJCfW7/W2DjJGkRLfFHr688
bhJreyd1Ia/zTVaI1Kde3L82CPB9cuzAFZdNJnf76L3OQ1NzmDo4wf30seLLWg+wu6e1gB/kiDYw
BatppJEiLd87TMhVxsdrA70eugRJk2KstuBtiYsd8cq5m/F4nVUMP6mNOaLYrwj6XPVgYjH5gu2f
UMjv97KvaZ/2YTNj27NJ46UBW2bCTOnD4TW3UxWnCLcrLvydgH1nYYiZPOt6YePUx/pbGNAH30VE
4Km1g8HPRBWmf3pb8r4452LshFExxQUm8FPaFp6vJPZs9U24SWqcCl4wN3f9V8cDyLxkYNjrwyCj
Fk6fy5x+ZkpcpKu4dDXBY9KLNUxXUaziogHQXGukLNYyNi6GAIyJWtUVw2t3IrSlKj0/J18nl05m
jec5sslaG0gkcw/Y33GLup9WETOAi0cxj/xdK3Mun8VVkL7L9Bzas2gJ+i6QTROoWpWNjQ+BwYeJ
GByuldda5x2640IAz1xxR9bmaA6KPawpiHTh5dQHOLM0SN5PcGTVEH+2ztxkVYObbsAPby+9o6Yl
i4L0JJVWcTTKWVF5Cymkxh9mmrgjzmUbP5W0xHQGwKAgiYkl2iieJIGqp3BgdexmBVliPcO2W/EQ
wZsEXmCrTedI6tWAMQR0tyfBRwlvTIojkRjKHnkWoG34dfSX2rPjB3AJiYZOjTydLXgKvUOB4vIb
yO39uMxDGBzLkIWOj64RMVxw86sUbe2p7HFY3rDq1T5lG+OTOzAHWCx1wOsrkgEerOtTSWXdpr0a
Zup0gngX6W1jOmVX9rQQW5RC1y5feFRG04v7fTfARarI39U4McJXq4zzQw1+m4yXiXbEN8XAOK5W
hkjzZGVsaB+7+yqOyLV5a5rIlEv4bFDDV06G5H107sM2E6RhH/TPgJGE2++zF54FLSaXTWPKJSxG
gfdHqgLNxWqVLUF2N/OC4oWH2FG/ch41C09YwuIFIJcMULp3L6loXBtjtm2eXw0zW1Q1EDKhe+3t
S2gvl+fJC10S6Bxqe/OjjmBcPWRZKzv5Ki3R/WpSyAD+uF/8AF+KUjeGQ3S6CDyQBo981thddAoX
vYTxEJf2Ru+3j9SREHA9tayTbXxzdvzjLyWHnPCCq6C19RE+mxzW4BMSL/tpHYsXm4NF90gyusJf
IJ2WL+d/ebM4KIQ4wocG5x4o9uYVwvywtBZYHoX0xFJXE5viclt4AhbTI8YbO/5tHHSBD9H6eXQK
Avvtj1ptrqaStwe3QWcZvqQWXiQhRHJWEuhDXr+IJwzY7o0qNUXwm3lVeY8BzuyaydHGKLJkIEjX
l5FkSyFIgAmETaR5DowdzgJAq7dw7a3pU7D/uUoQJK1dXVsc5S8h/X6kTOU1qsK0419OlVeGZ23Q
be0wI58xSuwsjdbuVyuOYOe4Bq7OqbiRZYG1AnqDkQvGYXqaGXGGYkBkJhWGEd56H4d93kBEk06M
QKNG5yTiJR7G9sIgYP5AaMHaN33p3LEpZUI0rHJTz9fJyqL2H1pboN9enW2xpMPulSQlOQWdTgPY
yj6JitlMV4e+w1eIOGUuB+ik4wh+NMqbIxtiR2Vk4vFjoJ0fcsR9SX2VwGQco7a30RNPuJv9Genh
M9CI8IS+lbFbfxAXqgigMB9fCII9aFYnJ2oylKwO2w7Vc28BDY+wyQx7h7VxhVH3W1jxGud4s+yj
E7AjZBSQO5CX/cKXvaxlFtpwxIrFnzBoau26NjY7hAcnhgDidCFsveJd7r4CJkGZ+qkCwhbGCcvP
egpZnNfhSMY+CdWO8Xkd/qeItJfYFSpfqUzAE0yCSWnd885vAvIgH0B+J0zRYaXWHnE+LZkmFny+
pB/cKppg1zReltwM0HJ1ZEebwkCj1YANViXJbov8ugbxSHGWFKEIT9F49PbwMB8JmbiIP2triVVW
74+Om4/odKzsOHlfGH6EmXD3txJ9KBBzsZDGzkFNpFv25Agzzg9m4T276o9XaO8viUff6Nmdk149
KW9qLelpuviWtn5O6r/sS2tju6M/HkXKMojbD+b+v+I9XtMS9HKCQtblKvRPavus748t6PqWQOAn
YEjmlK26GbUfZdvJwP5x+rT/Pbphj74sbzi5XAaOOklJeuo0FlbX3kdJYjwq4yGR3zuG+eWKO6PL
E8A64AoyrPAQyXawoOqOTijHCVnu40W+Ktot9B94nhcCWJKZ+6Oxfib5WnV7yhmpe8QfjLnd4yrr
kzwRF5siskWFwQnqykYA1zmjtZVsB1dAGhfyenXdqqOmTHneV+9ubOeQecPBRJsPR03VnOKu82cD
x2TwpJ9eq9yIZrgmdKnx9v1dDTWCsQIRhHITVXlsdCO/lzcezPy5+t10xCQojXWr2mbx5yaNEC4M
DhAFGy2Uo8dKxUpJpIYW9j5ivdmk8jW+8+KTiBTQuo93hCBr/xeIHyZ3ZC2/d0Uc7KyHU+dZVKYN
nGN7+gHEnODXdTHwvdXqCJjAB4Xndo3fixOxaIqVEQgVSWNnxF2enl4KGsfU+ylTso60CDuUn/rB
D5paZ0isBf9mQkmxwFhIsb7wmD24U0dmX+AE9RTaWWcutyasSQC0blF6hNNhQ+QBO99jr+clVlg1
Q1lcL4DnRMGudpMLjKiifuNgF99ZtCpnWnQKH3tRaz5Ny/wL+xw2wz+UcZxx8V0GS9WTQTLwEm92
Dfuy+J7J/5PDpWHeXq2JyrKq9MbukrT1Kf9rl9qyPkrV3fprLrR2BK7buUkaR4jgdbl6RM6ud0R+
4NBlqtBNL7QmzjnPXlaE2QZ9W61EhHOjs/IgPgL6vCOvjKeL+VdVbESyJRz1NXHEzqL0RgoPxd1L
YxIyOpcZXEpEn4cUi+oqFqRCE18sVjZF27YmA2kjvMCNP5JraywwVh1EglKiyXrK7RAYxhoDyV8H
nxxbzJSKzmjxioSAiiGdKG/wjzEQoGhc747UNiV89xhSXAMy/rBrLYqbnns74hXBsXzlZpvXVKWm
TPyQwLmrGCqvLrCDsrF5XxKOtuj1r/YmK3he1A8xBdbhaHeuyu/kAGR69xHzsiD4PyeEjINssmmV
OMpdgZjgnjxPBqhtZZ7l8eQqB0YYEMMWm73obXlL0fZlXzLj1NaEjpVNbQMPF/m5e6vw3IwCW+sm
3NGJPRgUXxhkuancwDpnho/bE7sJXRYYgKiNfQUo9lIX60rczHJ5GwF02+fsZrueMcpzmH/zutWs
G+v1Lxr0ARs86luwtv+pxkiRCw2nQQ5kA74V774GEAwj0iQqtmYiXUoY2el0tk9OqMs8WaDrLJtA
183yWJYDkoNsB1B4wG2IDjEYGzfKIqXLh48/3nExRk3G/W9yMmbDadurZRN+Ix5USFChkf62qGKe
rq4MTDh63eLEvwMNVkutjtY3r3DAmaEeSorrTDHe+SUhPiVyWb5d3fxEWayrJee7O4qeFAVziQv2
TVPxE5UvO0jZRYOsQPxxYVZILOEeUdRGe4ZA2lpxco5YMN60b/ucri7P8Rtuw4w5yQeZP/tLb3/G
eXqqUGApxsxYd0WNfW1QGveMfSuI7GKIznFmbk4ceo7LPP1W0lN9qvLiNiNRd3HakZj7VgvVxUpn
K7kGfS7VGCR3JbKv36VkZ08VlnRSpU/3b209M5k4ELmRb8HXnsz21Z0iUZoMp9DAJbPbab6DmnFp
PT+g/dbLwq05TxoDLrwy3I00G7Q2RUHkwU8Ddbf43NpJWuRbXbJmIYM9uIKrnW1idjzidpt8Le21
/ogLMrPQIE4RQEp59fRxDplAUQxQC+PYR9rXvKxVRMR4RCco8ASs4JpD9f89Fqj+m7FhyVJu6Tq+
Kc6LwrXVFXXHH1UscALXdrIMVxmB6EywO0O14df9cwsPfIN2Vlm2G0mlixh+/iH7B0XOJGZMFBnH
DsLUxE0fZrJQAdTWg23+G9HaJCM9y3+25eMs738bkH5yz5ZPLstIuim+yNV/Uq+GqivmsEXjbrii
wPleU6BTFlbk5PdEYGtFC3BrFovIg4KPJ5s9V5cplMiGHIXZFp2WeK6UKowzy/VBjYUQNGopOASv
x0Kp4nwGgONF6tdJnEVusqf+NbgU3HVOqxTQr82P5edeWAsUUgFwN3xa3EgdjU18VY1mbtDFDkWH
G9CH5/nQCUfswHkA/qWzrk6ydda7TpEWjzi1Nz0nIEhUg9dkL5RAxpOJeHCtKicRpit3OENEhZy6
gQNgTpbJcSeLJGq7rcp8IdaQ/8kix+HJc5OYMEfvum0fx5qiPDk8sSZmy/MOn2rZ81Yv7KHNCa+x
eglWn+Vll/cjQ9G8MLLEM+d2DwdO0gRQuOMBxsp/buzy0F82UsoCXGkeeXJturcwG61gJCHhw2Tq
0dgbwsf+AiMP+oHHWEpqVZnl6LQQ/i3rtZSzFVO1lRSKYIWVvePo84uQK2Ox6gNwykLvL1B9gcMT
mmgyYznipkLd3yGg+0vLtEAwy6E46lUlADGFvIHEEGrpgG/6KTkL/I3sskDJ8+gpjPoVX5IAUYjV
dYgnhB0m3cbWhEkjiyJXOONP3C+I04vwcDWDUvPRq7FtcYxFZtu6H0p7+ibdJ62Ogd85qzHl69Lf
b4zua/kNLrq7d7Lc/Ic3STzY/vd1Jl2Wf0K8hH484RmzdU5x2f/D3QY/LBm4qL9JLibt4atkyF1Z
po8dBvAia5G4246WwPRNDCTehxJdtZCD2y1d2+20SVJRD8y8+Mbux9TAmDHojLwR0NLI5tdnn/lx
wLzzTm9yhYJtHo72zuTV3Z6cUtf8z7LhJ0m1FgVx0ySuz1Zj7HNTlpRAtcaKAUWY5B8AU2t41wtl
XNTvVKsooHbaLVZ2Wss+ROUUfRCl589SIw0J8IBUshJSc9WOI+LwjZyh0KpwamwxKeUT0OOA1C98
PWo0MdBF/nqIMHXvom2NEzkflSuWA9dHwGRaNEMtyBU3aVz2eUclKQFxYzhU50DTnj7yAPG8sz9/
rlnMDodNnBMO+g2COvHq6YjDRYolv7oef0NZrB+7ibm0s6qs+dzYNgXqfn/q2zf22fHdMUwzWq0l
2reBia5e7Us6/+HI3VK3D5TuV2hFR4rMrWblyfqrGq6mgQ8MIWbb0dOy95LFAoWn2BbT5OrM4y5e
5UQcGxYNI2uN/nNTn73d2T+81Ijbqm3r/acM1ilX6yXjmHLN4Lu2jRQEPg88W5MNKEezfqdRu/Sm
8Lx38jz86qEhr/UDEhICCLJm/rGU9W4nprUJnNjlvG66DgR0YtBiGEvX9JO2MGHRKlWLfZoorkiH
5wAlwkd2BbWOBJAeFxb6f2V1OmI3XBoRdrxryEFfKHYcs/6q8CA89Qow0Uy7uoYqhopmUMxtuFoy
nzjOj/wRPp9pGCv51EMFscrkwyTFL7YJXehhJlOfqop77NVjbkUMElo6uFrvyVSIy1T/7YkFp+g5
+DjWm4M1Qho7RqWtPrrTiXnxrzcoUalD3HHpuVi8ri/mwEiiAC+0KbYA3fXbd5tEUJuKKlV2bv3L
ugr1lrgMZvN5qs9j0IDEeNq0nsQJdXuFAuZEvrx8XOWJBHLDQpwIBs5409KyskCm/gcBaZtcOt96
KNLqm33eXcdcSL0O9L9VTaTQ8yUixiolkklbMXPkvoJBdr26tua4ZfdF9neEc2uZAYE7kPo2QRwR
bu8E8dX7MjEL7qwTRMQ0ySrZTrF4aZ5fnnV36WgZ0JT3yVPU8lmUtxsBbeE3zKIm2xwzUWYEIOez
mzg5hJz7aORrjITiTMuMjjHYGiJmZErW2SoEj+Jmtnu0DR0Dkg06fN6eS3VU/vy2EBWa04wFaW8a
eCFJM9nIbpXEMMSkxAfxRLUvqAFgBNg0nLCsNnUEiSBACzkZPFqyQrMuO4ZO4zvirCTWiq45GaaV
qbusWPwMwKG9P+vwIM6AacYcSME/pkEhlOVEHIFpIwv4o+yxmqUFHUKL+ZEE9Mmwz6T8TQvzQ1qr
kTmUFcEkbmDudzalCDknDfICNBN6jRAe7UX/KYs5LuPseBZ+U2EBviexJJHLhWPoDXpUpOwHX/Fb
JUlEoNWW/ngTu/QGrYrfD8OQ1m/tUmQ3g+KEyBFAshl4VaQKSKn/JP+XGVCoPGMacK26Xf832u4S
pPGIl9jjy6tcOCUMwX9zrR9H0518YhDxOoAUdjn4Vs+YnNWV4iuwu67nXvoxwbKIIq03BEiCfm6T
4RrMEbQxeErB518iEmDHM3HFyvrx3MlJ18L3HOuRCGbvrA1BXL6u8tkuhNBvrAAwf7HLKURU5Pmn
0nCVV2v7dJuzdGqBtKvuI5dgo5BbcNjr3JHd2kQFH7xWgZUHYjWDxXatsKlBzhDe/B8tnROSfPP5
SDKO6JXK0uCzm1yrfNJUEKBkwVyAyg0SqXN5aiMqGVyhzTDi1RlT4juXn7KFxZXbwSQkDrqqj3zi
QO19BBYFRlToON4OOAXtZEYHG3AaJkd5KF2Qym1cvzS7HFkUBPuX8v5URH5qlZYN6vdPQ2vx0ppm
jJVO884zVzSPchz0oGpMCnM02wlucAl8Njvb6WMzNYOd1petd630FlupjbCdUfWQZuZOGWd4DyHm
+GlkQZZLZ95LcMhlUoxz2k2PMGzIpeSAMNUky5AMa3QbgG+MNM5W1S1ucx+96saYTgvhVgb7Mf0m
VDzRuVAvYdDopYQ3yaa358d8CPNo+G2QPcW5rXJ5AsJfGeRmlh64Wlw/dXCA5ebXN5ifc0T3Le23
WODC2nZ1zw6jNx+10hHt52NIRVTUigrhW+ocMXF0jeVEPLqBQEtvDsXRWc2RhbG15I7E8KEXMctQ
5ihetsWmy8/4phK8hmQVw8XNfGJCRaJ1fQiQGrm9oh3cEsxxMHVF2OsRFYw49268cS3xbXIU02yf
sGw79P/PYlcR92ZlsJY9ZOJAdLWXtahG24Rei7PzdEpDE98nVsBk7VC2u/gbb1Zr7M802hqlx8RV
CcunwXTi+7ohtIob7iWIT0WOc/Z0XTJ/Dbg9vpoo0MKAkIHbbOiDET+jeMX9IWEqXgGtksfcJVUS
CMSfx4p+UZ+Sz9vYCFUXTGB9+pBhET9ny4mS5QrPLBDROCjofO/NFjmD+mssixxGPf9RLR+Jg9jS
gQyvd8WfAHWVo7atBpR4ZLvNdysxl6+iQzWU8MyI76X+Spn0LO9CfSo1R94xmKElc/2XelxuYAsI
mFRPAHHni0gSZCFz1PB7aV6zLkoH2TkdfVHAAOuEZ8q1CipDx+tj56YjwNAkRc09IYgfKsnhbsD/
00wwdzQtvsWhmRzJAEyqQVTuRL3M+29DkslMW026jTB2VZk7wd3Q4A8ZQBS4FXaIqvfSYxlXnodF
jN/l4ZkTbgntYwE4NL4fS7M5nS3xBbD8i4/eo1IULLiCferVmkLTsutpVnV5tiaK2N9NYxLdxiRE
TkfYDJ8wh+yWOnj6NDV8O98Hzq1/bbm41ZI0NnEjgksYZ0/lvyXMfnGVtPEQN4jdREYvZm2/VAkC
7r9vBqWZ8lJeWctC3qnhCKdcxMSI+BtAx4o1RVTWvNxy5YCNTbkMLtOujdxxnq+4wqmDfDS3dtyb
UDU2pwzSfjDgflC1q5PBpM3/LH5EeUR/ScMb8zvr+xq/zkqGPGUvDTEYhCMbqGhji31c+dD6MmdI
jmRoTarhztlOkMKI8JJ2eIQ4KmZwrgUnMksjeljRWR7CuSzWx9HMkJ6L4UkXnD2aOrPuIclxk9Mc
xM9xxhKmYHMbMpfQJyuScx3TsPMG18+gOEOL1KvNpAcpeKdkgBP7gxj7xQlKTwsoOru/2VtXVby/
BWd8mpVCCjSAjk43NuDHfsM//CizYBZl+texd04ao5zBDZ4omSH3X9cAID9LbzvMUihzL/YGAvrS
PIsQNXZDbt2O1HUYq6QdH6yEJYzt94do/Hlg3HL4ZOWaBNTW/PW9A/V+7iJdSgKVL2xKiLFWZJLX
wU6ss7IjbjgULWXzUTMSTwE3xGpkDWTHpWnc5GaUq8KFJrCZ5HyjiHFNTQtWIKHBhg4y7biRgHGX
zgoV7hdkM7N0iED8HEdeFpoJTmrJmRq4GIOlOvFzWC9y5qVGvWnlmbjQJMEDkOgQvt1ysB38OSj3
m3GohRTvJyqXb5rb7/ng6uWP0zfhWQxC92CuoRe9tKIHiLPOsihZMWtVVBuTqrgUU3K8ecWAmo04
HiQ9vPhs9SgvFDjvhXUHM/TI43mcXl/72066PA4aplEgiMhQKbe1ZEeC5GW4Lq1yiNRN7+w2b11U
aCErkoCJ8T/A3kbQ8yEtOYwgGXiam8A7PPRA5h9znLG3s0VE7v2CW23J+OyyJ5euI2p+ZhegeiYT
wHl74aU9hG/esV6BAVCLjyzi5gbKzlXLvOzWVdf60VRTmGJAK4iEf1TdQJR56yVxhmdIV+E/umGv
eeQUHNStC+drS5T3qIN9rTBpGEShOe+R0PGEBYusyVOIoDhEqk9rBuL6EiNf0SisN8MRR87UlmBx
/gci/p6zXZ+Vgz1JpLRZIJfed8VbRb9ATOsgwmeOFR3GNSWXF5SHLp62hNHFfQPt7lZ0cHvqEv2Y
G88jcdDmxLRb3DKKz1AAXi1lPM717W4kD9f9p34ttpHJYwl1L0sZigXvo/RyMvrGCCJ2xsEzli8t
pR6CksBEW3MsRf7hmeTvCDxbE2qHjwbuli72I3NAgfyMY0y7+gAAgcGl7CekVTw7LXYC0bNaoqC7
mS5fON3dGE7YW67+JVz0FF3wChMUfBF2sHwBRRIQkdOdMZVOljCpHHsZGTh0A1EfOrHHwZRbXGFV
bsTYGr32k6yf1tJK/A/dJ7wsCDHLy/DKuB9YFuBBWrQnYevaBUUU5B05k2Elgr95DPx37QSvHpjU
pcl7cdG/q3fAO/JXxbRpvtMemj+yOcLzzj0AvUZF3teivGeEnwWa6OfRn+c+f1uj+8Jer6JwvH82
QC3f9WkDSi3dJtai4N3kQ1758N/pY7qS7FRXTBC8sXl2DjwNhZfEo2inRAdWXdPIDPlQn9+hdwvI
oPjYUXnTtrq09Bh6eYGyxviBBHxW+2yEFbd8fFxfr77CmI7wLb2YyIzULbk8LNI0YbOHWI0sFbnH
P4X9SXcYMbdSNC+sw1TLkgB2utP/RvCcXyQdxpI3ps/+4iEeaBBquulqiwtTz/SSuWQ8ii+Lh7DU
0ptlCT/5J7rDw3J/6ay/kHlf5T6W/KSB8elxFve09iXOZfPv2QNeMkZggj/ZoyWvfBibHNslP1+q
Dsa3sT4EsSG+1upM4tC7FJN7gsdhSCCGOtqdBxFHXrmKK0m7AMz77DN3jRaGzaCASyXcqtS2aPB4
YTrzi/u2J5awCdsC4SnlpycFWDM8Rs+mbQVU7xXdzvzhxc1YizRkXH6x/B8n2T2SeIOIpsBTwl+M
SMwNXM68EGEPm+c3riTuNq1EjId8h5P/fQ087rSrDeyAYnQXRQdNSrVLGshxYFVsIJEZpXFbqZaf
OYLAg3eePab7tGFSNQZEr7qe5mM03zNgn8MolW2Unrj+NfkhMXDIkyH8Ae66QCclAc/LlrfW66Bz
xIAPJgqqa6XyymbUryyfloB1RC6w3MrTy8nsRekQyN4HMuAQIWVE+BW4Wcg8HN6TjRTj4JzRhyuJ
kYSNTj56YRsyHuYyz3iZHw6tFG4eTPh1BdJ3yKNf3ihKPny+r3DJRyk/x7K06o4NLA9rq14/Kq+C
R3Pzm3IsW6P6yiNU9D+eIN8n0yDCREny2oqs0pMOnGILtAQhqjyWEILUDKkV5aJLSEfcCUSh+ZEb
OwKiBTpGkQBmk+bF9GrrOWiypbsDCuwAhTKvFzQ9fT08Mv8xXIHFs39rwZZ76X98MFGNva+A7oRU
bRkD/wl7TAjO/ULX2+GtK/DGOAvhx+GAbZtwyxGGDreUxOM0BVaolgtg7valiapJG2UdRuKZKa5F
9nGiVXN3m3FSaHs4kQ/HzBhn/ddpWR9A8BOaG3L+K3gmak9K8bo531zbKGnUiaKoTpGu3ExuASUl
8PnWjrJmxQzhDKZXQEC5H1AAYo8R4o+ReLAr4mpJ/37BZ475Ul0A8x9fmRP8ekTotoBAm2FAO7WM
W7IIHyuntx1mEsernf+3se9uls6xXeCKNr0GT2VvfiPQ5UZqv1UcFCstBj1X99bhv51utOfQG/43
cpx0DAErMEbCehU6l/nYnZJGIk4l66b8/zgaKy6fmvk1pe2WxCaMHssxiK62qhUfG9CU6v0Xcw7S
xe/0IP2HvUTdgW8KoaxtZCh1Wk3btQEy0rjCTUphb4WsoI//KADPLMG4mHv5qQpu62hj+1yzkxkm
Uc3+3VGhiUSvE7bmODFzskGE2H1lixWGVxEy62z/tPrQ/2w65BuzQYyfNnBzrlO2RJDigAsSRwt9
gbtTuYDGQgahGFo/9la8VXJhg5AIOSVpu0cxFh8D1FRPepAXNB+7aP9zRvvpgpeZMB701qrR9oTb
EeMXlqom6LRc4sA4r9Onou+alx3+aIxfFgy9nQG11ldXS0Y3iRjK+S4vn9Ll5EVA1oQTDKl52M4W
45CdoIPzFpuxBa+10Ax0DQB1NcC6eppFPAcjFnN1cAlyJiOPpj6ArMOjO2tvWopjiEqJuLv/fJBY
6erNHx5BglM5o4BwhwTeybf5XOcYfWQV5B0yJ7bKBknOnXAtIm0rF0l+5ZlFQVR3iDNecEB9FhVk
kBhmlr6GkxaVzRftpQuNDNs8VlzwGWUnNM6eEZfMI0unAG97kEopPrEsDix+e1VfC+tB41jQWeg2
slIlE5UOHZSO1CcuQBTxjYXptAsNemn3JL7Kzd8gvsH+/RSEkaWxhSgdBAD4R5Obp/YTxDwcZJ4b
ptprxdpugh/W/wLXL4PQIJ66DpwdZvl1DeXz7UJfTojExVn0DdlbhYIBGoGRjqLmbT32aiKFU7EA
BfkhsK6ERX1Iqk/lNl8KqGiboSHWVN2EtBun7jY1F7QX7tfNLJxloHhQ4FT+NmxRzvzz2LYlHl2v
gvUKaefDxd8SyWhaXUe6UlVe0fvGIl8vaaMf8H4iUChgcNOJ+zyNXwp2PeZcK65CDTKJ+LBUQm9X
a8A6Fr2C0q07W6W+/CBjTMm4ZpWPdr8e5auDTkiyjdYRvKXQaeLC95jD8NzJrROGavzWmtPWCrx9
h2xB4/VP/kStJxMPqnw6xyBjMqCSNIw02ro9y+iOGzs8098TBnj9Lw232DyyKIudxYobRcNXbxuN
iILjIg8dmyns1/RQTLki/6rQLOQjBsoPhjUVV91FEx0NM5AY1zS7xPXo7eu0very8li6qNngrWtY
ufMIM9ASaTK17wzL4p7k3vJF3CeuWGZAAnr+rejXZVQoL8N+k2rtuy9J8fk6lzsiky/GwNM4/enW
Xl9ZeFFnnN2V570zE/3wwwncQct5wRbUWG22HESUFhMoYoeTllNTTC0Ex63LwKcUR7xtnMNrk96v
mQ/j+GCTxVBZlLjWtEaWokmXAsx4r2c/oOBcq8O2rqQ6RDzhubQ0VZ4A+YWXqsQOeYeLlAFLZpr2
EXkPlTW2m3XGpnORft6b5Vg+jFXe9a2BzHwocx7a7u88EzsaYWigV4JbZgtXe/RUTSmdwY9bhwOi
XhhGdF6A0pzxZ4KOn1MtSfhBcx1FDC3EKBkRquEMdAuEoFqjt9OKeedUYQmJh+gX8geCicTX2CK+
srGvJDYIR5EUCOLzT3uCWpJdPwYoP98ftG0/RseitVmBiGqe/kPkLsIQQfszABN7FZQ9EMuB8N+0
DjQl24wmGChSQRWwAq58FLFPb6l4o5/7xtL2m65VBgcMnUxlUrGjTzrxgbgUVs2eyhu+ox8Y/nZf
RMHY+sJCRBxs1/D1CsIgMt6juR4yCNq9sZhNz8S5//GChjpxXXDerRdgUBdMvej+3mfYQ19xrhMs
ohtwMZg1+OI3WYFqcVW1YbfwqFrQqwQ28Dw3spfUqF/c0PThMHX7Tj1GrbUm/a3JBi6g3zzoMjLW
JKHg48KyJbUBSSIZmxKr8YIUmt5mtYIWVUI6BgjiRuo+ufgzTTpcjiLHUF624oEGD+c3NCa+PnML
tj/PgJK2MVgOaxllCQt7xd0qls7LpERF/2zxiSjrXN/EnK29R6duh7NFbXOgdDjRHTzcinedUaQc
m0WbaHj4M9zIyF+phHyZbY/BdFcBnLWqW9kZ9fiHjl+ofyOtCkjGr2LERqCuPiLRrm2uRU8wKjpo
CldXvdc1kUwS0gVWadfC/tlMhHruSwL0cO0us0X/xQXtDBV+3RaErEbzz8ebiZpocyAkjBL/9jrP
dXM4iKSp43N/kkj6EWkCWoDNEwpeNjIbDH9lnp/HRNgu3ooWsKAggLNdoTBImuwfU1IEIWojYIbG
errRSGf5ZZeuCwOIgJXmTPPcSurTKKze8XOhIBoXUDC8kUZYgh+gscns35PCoMySxD3KvN2/C+ab
T5l6ibMjHKFKTd/uovyJCdHtFUKB/AxHM2kqKQFn/ahEojqRgGLpC4o9NkRWA0INe0CA1I9ydH3e
IqMJEwjlTmSZCuasemyVvzq1/F8gzLI0v/s1y/3qS+4GcSDTLBHSO/WfJoM8NBOaDKzI3FD6Bruc
tTqSY6LnE6gsn6knvhjWC1qOy1VMOf7K4/H3Qjl0L7ThzPi8CBfHl88vkwhB1MBJtbIBeT0tT6hH
Inw0WsLCx3dLd7qHIWORv2u1/Q+lhoUOMgulZQke0N4/tMHKG3peJLziQ9udGAoE+mYABRlP1b81
mFkdf7sx6UGPC9YfCGQNLALEh0/z5tqZSAI4ERLfSZEf8sWux10z2zEQ63gf92nrGIORoYb6DnKU
XbcqeuTrJILOuGjLpCz/KEXKnbAk0u4/Y3WvBWbjL4wiGlzAPYFUxsV3HaBLZ6ycIPKu0sTteizr
SydjHUNLdelGLCa76awpfgLwTEn+crN1Sr2DH1Vs3OYCA3DyN/4tGR9igHo5150g9sn+25WI/wGE
a669sQ1TPz7cbPOlNmRv8IA+uuw5us9meOI3KglQdG3vdVuX6JD5usfTaktwYAXdjyuNA17XRUJK
/kdR93JCyCPpw0rsk71HEzWSvlDcAARCBKh6IxQJqcgrdmUdUhNuz15ymkbT2FclgDRox2gTO2Pv
boA+qq/RIO3VlhcG8vpVPUkFDEJtzTnezp+ecUmpKm249nnYClIq/wEqU8nnIcxZUVer80mV5QN3
hSQruLNsspwGO+Il7FiYBikYEqKOyMl0sZmuH+1ATZ4AOTKC10d/DAM4OH4bcT07IVxJO5yXEop3
f1Q/zNBQMKQTBh4Gfhq0TjXYjfOHzODiOlBqBeYjVN8xu5cv1il9oUmkUXUHjMANTqFfOi1swZWd
TlZ8D1MPaKCJ4rSikEyFGNGXyakAIZh1JvD9s/KWNlhyPYaPrKK/d80/Kv0Z037+cNwir3AU3qK8
j7UvvAEQ7GqdjQAHAxKN/mhGtCRFjQ3AjoUQ4agBBbshWygn2mIEvh4AfrDdPbKAuI6lDVytZop/
+g63YTpLbEr5/vsx4oF13i0SxLHMqwh1UJ594Eaq4SN7Mw/tM3b97prfq7ci0Bsn1MpoVcPPT0ON
rL02+NgRSl5Mw+rIb828xY9wDHoPtPDupM4AxRFyK+svjAf0wlxghaT7K05t1kzwa9Nb+vJsJse0
MyCcpNtSbtl4G38bGWFYZd31zYsu4ofTMo1vE86ko77PZKwaOMrhAQzUkdNbjfqG8LDuVkum+wss
gj8aqjtaA+jvtsi3hJmGnnZhRitZYN53cs2SBdP642MFt13M6vldLqcMc6sfJGC7sJHK6B2ztDU2
4lLnPTU0QfduVY+5ViQIjImsfOr5tRYC1ktaWOFb2RKQHuC5WasBTs3yDZB9CBy48rEl0IfkbRf1
z1riTKpjvENvMGLx1odjx1Lu4wXKyM1j1GEUr1pXuO5Mb7WcLg6jcv4IdBudPsLaGKy4QRscDYei
Et/ynkvNZx+aMyobQzVOjdEJr4xfiCzJzogjhMrlJiAn5rhdmoc4MW1OtRc1NTpW38L4sgFYWHgm
wInoYGgjLkEFTkuOu9314/pn6ZOM9CxwAvbVHUzSVPsWD90CorZgoJ8vyht433AsuChHtAXYYDF9
l7Lu0PEWzw7rom7OGxC+yTToDu/9SRbh5/tkAcB6pObyMkErI7K+MdeqeCZWX+pLKkcE4Sl74fjX
yquaUQKt36qbD2xMHCGntKvX4aRMqaNmRMgm/neDPpPfBu7xbvnpJ+tl5j54eUYmWJ5Q0AMk3J06
OskDZGlA/gYFRSdoQcrrw4+bKVzibqFj/8Q4HZt1GD2IOtV/HmLsK2dgxf4wqOF78B1+9KHNeKt8
LIFM5drfaw8szO9GjOTbqk1Jxt9fu725T+TPH62GigSJcc9s19zksYdEyIi+ZKAY+OyaZ3wzMRvJ
N3yID7egaKve6bcX+Ju//v/pQ2w1E1jHcEEH5ooG0lpaofMXca3JChWqDHW9dIR6sLpHDg9xCLRa
8UwyVC9GQDcH2f9BGBdNv3dxNb2A7Jr65ROvBQfOnCgKIkcn0O2abxCM6o/2dZZJlnr9NvTKD875
yfBJXMuVy5pTnwL2PqzwqWj5GHDLeEwL8Et1xcOV/90nVYJSWXtGwGxe33apsYj9ybSSVN2p6AJ4
gfx9HgxHgHICIxhAT5q5czheZvj7JQtlyU005wWUraUAjbz8NbWHeCAcVfe1/Lj1DOLdFoJX4R5z
gUu7aYO6j3q6DWazVG1F4ftWbiQR9wMChrOva5l/wXgm9ItraPUrqFnPeCMq1T1WlwoUSTu2fL8Z
uc+FHE1L3aHu09XYTSYJfojv6FgfiiBA0HHovtW7Qx5G0ZREpvFk5s0OWVA8fnHpbE9a7xdQ5yEy
lGPXH3sNT7cakliKTWc7VWXa854pJ6HkO2WaYW/1TDCP8udS0RoSOvoMTBzeoebeNvbVO3ljjBx6
H3NGjL+8YR9hDUI5h6NPxrveN8Bxz75Ee8cS4KMXi4RjtQTZeg8JfWqcthm/9+gso1ke3up2DeF3
YaiZO3+5b+zEupZvIesPwmqBakQVLlBcyzpd9hubbjN0aUUrju+4Jaql4OltLouYAVv4I2EcYe3K
58ObqtECfvskumZpip7mlq6Hib2yEB7Wrx/fqup79LdmWJYdCrrV3FECvWoeAVcTdufY2+YyCrZQ
31qtSUfcKgHmXnvu+Ht6XytiF7H34va1oDA5Gz5Miw00ONYAuW2P12CNUMRTUxYNQ3CbUKazsw9z
wUEXUNwtF5tteaRKG1Pd88SgchFHokNwpIp5lmExyU4xBpR+G4cweY3lY8WsfggNtuUTjnfq5IYF
MuLrk4/7yhaqJ5j9AooSaHEzZm7iHbR734dz7l4NUWSA3hyhjGOQyqZVHMhLzenZELyzaeT5L7Ol
oipKqb0wPuF10aCUYcXcp0lLcukuU4o17eATiPfno5r697UMhgNuPKcWUDHO0vYldhO4I/RpVegY
ZCmFTSFdVczhtr2qCraHbyXjGnV0/Y6e2gDPx+WrJWTKW0BXipPCp/FjMS7g1TqFjMVKXNV9Z8M7
OKDqn4qaIj4nOs/suZjVSXMWdbzxUTzne1UwWD/yuB2vFKucotWnWMpDJC5yWrMXikmvC694PQXv
iId1AhUPvMhsk+PhRxJt5rtcdqnaM22O//bfJgaDCbF0WQErFv9TxQrpFpuS4+zVd7oCZmqdOQQn
/BQiKGWOPBia83ekys1nPRQ0wj3zUztVtBcGbNFqQ408fLR2sGH9+Fw4wkPbG/Gcfx6L5US87GMH
WAkRP/sKPRNjuq+7Gk1jxeaGMZqoEv4SywFsjOY+nKAweCyofhDMYvN45nLiyRWsqNGSV7XalyRe
4asSaaQ6/VvKtDmILAcr8xsA4GO1XKnyTdq/Erv74q2JJTXG4ucoxyDdo2b0ksxl+h9JPPN8pwXg
uVJ7geRQERK8sbKjdw6XVHk8tKwKYwgAZn6VhtTTikg5wCzCK487tpSl1Qbj7tWYjXz4vuSgw1pR
2uQvkZQHtDEvQCJ0RG1DMK1h19FN5Cv93CoKioYHppN7595Pmwf9Rq1RpzOlVk84+F4rvyv/XW0L
YiYJ8d0t6sKkOGjSaBqyRbIaQnj4wIF3CW84u/uoWw6lIo9H9Oe87N7xY7qkpjWNZ1px1Njq5UIO
PoS3brKhYn4M6fVWbU6oHwGjiuEvWIBQc6TQfSqIeWCLjbmXmd413mBmBUxe2Ocynjz/8RLZGOqK
UNn+8Kf1w1M7IdDNDoYBbv37Sx/BVP1HEVg7yzTulHjP3asQz31T85+1TmrREmEyNdTfgIXYLf9v
879jFtNtn/gRgYbJrE2KHqG91f5b2938KznIdZVGVi3upZL3ZNR9yCQ4HkC+EQAjXbw39luG47UJ
gnfDuF+Nb/pc/GgLvgbFoHRkmd0Mw9+B7nl9/PuN7VaahkszDlduEHUMzdtg6IwLCu9db8eI6N8g
Cz5W22RM2dPwUA6Pn0gE9dWu/BKJXOj1nXfbUBP/Qk2RVnpmbxR8gz77+CZkuDEfQqZ1P5+BqyM3
9c1zC1rtcFMMweXWaPGB2mrRN5PSycgTd7vq+fPG7MaLUUEi7FCjmv3xyN5USvVu8ZKnPb4EJa90
ifuCHbl+4+dXyASDmgRzxMEwjcyzgOAjwMGcSLzOMuwr0AP5pITK6ZM5sxL5COULhifdUkL1QkqT
X8m0RDn8StonNDWhNz+5IO9EYPmou3X2Ec1+c78H01ym6dRorZRU0YgcOKuG0DGUjn9fOHUU2U5K
vawjP5RBSfrrNdLE9jQhV3DRQOE9KHxjtdBWfBKfnt5gC9ar8puEFc0nXohFlQYdPXlKNmyyyWHS
m/wIh3EPXpJEAPIu2RiZcS7kwQIjGxmaLYwCo9ePyBBdW104vGjwe0/bsUmUw/VSfpomH7C8AL1T
llwf2U6EFRjloSexV9mZQhI+bFTa11SvDkwvt7cunWZPJSGmKF4DSNMnfF6KjnVWrrKnF5nskNrz
MYaAiLlmr4kLVdw7HiQIEeymCiqNsnqw891BZOzjJqMiQRRfVI8o48yIUHj6FGBPCSWLfocYkMy2
VU5uXtroG+KWa5hugDR6glAZdLcEvNmeOOx6jcINSeFoLUMzs+vyQWH3i576n8O8pSWQxtUaBFDI
00B+btphucOpJw1gNh9ObUu0NZ6ucsi8FTfkaSad884YEO+k5xIiN0CLE0jr4Aq3vbwd99RCaREi
V39qwb4QfDcftgDqewpRGVAVqFYaJU79M7iPdXsNDPYMUVghscs8wFsM5oaHJOl7mK6uEY5jll1o
bn07Qd7krD2PXhq6AD4P+L35nrttSPXXtzh4GOqI1nmqv5R+5hLEsSTxP/LbEtf84kZ40YzANJe6
ZFYsLnBCcD+2V3FrKj8ZnueATEXbS9oksQi4cnBItuRdwgcoknC1U8s9FlfjYnOo3WamKiXdUAT0
CE6v/u3jROVUGJbLwO8enCPASChQiZXMYz37DZvWdQ/9bKPLklTdswNhPgaF7eYxY7RUmXSzyB8O
rK3UCj5SWIIV4Z8p4smbZ7kIQ0O5OK+qMigShrUcI6dzHnkC0k8C8AZLaq1KjkVkDYONUWsOTPlq
Mze1A/tB7dmusk4uOsgL+W7gEZmFcesEmQWunhXQ8yX8e85IQhVrQj07TS8uPmBX1E6DpCoVLeHi
RerVfUWBEwxR7LvendRJ3fVF1t/I710RJbHNXyET2rGRLDM0nGncnj9gb8wDB+OjLxQwp+WmP4jA
vgFf7XeJW0S1Lwizmo9S0lzMYothpdNqvcfXO9h+nqT2Ki9ZBrUKlcNmmEGXNeHemaA/x8WVnjie
WwojmzO1VcuXwB9ReQ01nNI3hJ4Cko5YoCCXmTfwiOOTWIFAfRPSTVPE2zGx3mc9k6H98B6AB9UG
V5iThVtA8SI9Hf9bXX0bXMY9r7AK9+oIOEBmXkaSpVxX8i774DTyiLBckGZcwSZjvuwQnycFkJer
l+DoECWbQUCJRHMzqfVynR5yUjdRWgSDaSQh6i8BI+ryoKfS1c8g1Efcdty3z3o8GBhgH/W8VD8h
GyBZ763T89WtnZfQwL+Y2gkrHyioSaAH8bLu9oTv/G3y/BEZAExLEW2SoO0sj5pfN+Z1IvC4+q8a
r6Wv8pwlOLrWyVuYUeLE4elDgA8zpMwMAw40Ejf6w6bp3Z3L5TkBxnDzRzpOvJ+c+CMKeYNSf/sY
y19/+upqRMv5xC0W4d0uHThSaG/w0hGeeyCFPTP3HZDsTc97YvjGmtSrYbfBL/Cc2p8IaARegn63
/T1YoO1pOhr6W0JZPGPIqS7LH43BrKVNeBPTzrhrPbx7Vw8QAX8NTEw4Wc20xohGVV1c1wAy0qZs
g8sk85HC1N0IHFIg+jjpqh3di9+qtGPz2ZOr9DQqQTtWjeRtdMgdW6nRngQlGKpr4NefthPBJ803
3h5U2yJi/vK1x+BBMM/6iTPwJt2VHWddTbwSVnsWgAfQcIXKP47vaEkmnRcfbb2vxgrkeqw8WKXq
nxX+fhMdmmkGy1c3dj2EkN9ZxHunxeRQ3Cbo7hu3I7wJZsWDBHjPZTLo2hzBwJDnjo4m0VmQu0TA
kYKSVJQLFl4ZYIvnY9iAMFSSzUFdX570VqwqAzGuqmTP6K/63KKk16atG15JMXIeSOk7glZONzFJ
k9hTs8qF9B48z7JW5I/kfpozGSzk3eyW47oaq/NyPLvA6cM4WFRN5NpaQoCX6YY9I3o7l2+YnN/M
5QLGcydeGgyLV5ldvrv4u+XxmixAr03hngC0DcTf7+kuks+XunU+t9Hhq5b04in0gzteg4QL++Yb
1a8EIzmt6zzTB8GZYhTTDNcopoif7RLoH4WEpHHrQ0dGjNDq6CF4/Mvj1xDkXp0H1XPsc1EMDdtf
TgwgddY17tgo38abJZz1oUHCtN8aYQ1gkUG8CkyLEEWKCIY8Mue3Wq5HeTrsV6K5PZGCHGVfoInZ
pviGn3o9myW50TWvM8ddd8+Gw6RzAvk0Fx4b7Gu3QLVGaMoFsOrgSp/dk3FK5Zl7NE8BGCzv0a4U
yzhKBU5nkCR5+8zu48eyhO8t5A3amzSCSrjJU9GJWbCGPoR/qhWSk7eg8aOAXfPSHZTppnceKLZy
0HiK2oj6Mb3KZrPgK4bMKZlAj4zUjxrPkYydX8DbVTsTg2kioJjPGhCvD2SpLAlhUk+pZ8BeXE8B
PFdianJZbdA6JRaT53UZpc64Oo023OvyBr2SL+muDS0LY2hPlOAcpbSlzCo4OtfFkSIu3mUc/exu
R5x9WeRF3Cc1wE/LPL7Y6zSN6Qvdjq1Npu24r6bwpBOcBuiXEO7zd8WID/Ld843oz/3q9pmYJJjZ
hKMTPP++x7mNWumfK7rtXX6CNmrujFMCcXRNeEd6pYaZhAvnApLKNrMXIKtIrAtdJJ1Ihs0376IU
+7GSUVpRWIF4OrlrKaE4YROCApwTaEroZNI2UsOhHVzOr6+qGYkFIVlQQehXu9puN/jRUmS2d7EC
hOy9SOMuIcLK4Yzu0Bpz2QTAAVO/KfvpnKD5x90Whdl3L63gMMRBbiAXH2k+I9Dg58SdfECx7DSt
N5VA6qivscmW3salLHBclgBz+mnvBwAiGdCSBFY5YdMWpK4x4zKeSLZ8+WQgDdtNH2psrvlsiWE2
nn5mqbCRuxioyrPmVE95k2hjylBcmKUecLvPRWSGyrEBf8BTUS0xfS1tLx5RPNYkjxyb0LOf+YGY
lIYvk8vHgvrJ06yHpnbJieacvRByfe5oZ3J6oZR493y7KC2oMThn6kqvC4QzFrquPcfj8jy3a7CE
H1Lgsgohf8LAIxkg5aQqub8vK4kYPWm60Ib0mZdogj4vCzEjeOohkfEjWgw9cwcOFg4omdLbNH+b
j1B1jpxat1j6lHbHZW4iitA6/2KFqQuNrWInRRJhmmvZb+hvgAtj6TBFsb8wSBj3AzGiDvSUv9NG
xWGnz+5K1lBytEPedehvoPCABtof2sGYBO29ZVK0uimdOvgR0sYU5ajq6zi6Jhy+KBuVCi3okMVI
FjmJN896pn1M9sY8PXISuNAx0E45o2OgvMDKV/7MIfI2RovG2bHzOvu8FUjKeWI5LxVbEEbMHqhb
dyFlLxI9G96MuCaBeFRHsb/vdhhGiwWQVA5aHyEImBnx+RikZc6yC7sYq+4y3E2v511lgT1A0EPF
EBjk7r//bX1rZ9k75PeYHGKMEwxtyVGDjRrQ3ccMoAu0r0TkyGoIrk+nssf8QUbrNtzHb/32wRQC
F3X4p2OVkvl/8ZGsuLwFKPbX2WvgjN+vGBHtS3qs/wOhodaDFVkjMfCJqIUEhEbHY+zs0+vG+AIw
jKootdCY1im2Yc/Jj8BbvCUhgja4tqH9vbeKfEi7AJq/ERz1pyzUnvufx+YmzmvNuY3PYmSiQoYf
bHssS/NMXDXrzpUuTBK6Ylz1VXEk7d3GZWd7EzBTSp3LAf/lMm5kD6M9w+ErwrnpNc8wwkDwBeW8
ougLK8DW10ip7c7B1JFLhhxE3SaU+OeNIql38R7Uf/GV2bL0ng0MREp5SL/6rbncNEw/x1yGPifv
EDPFGP+Wv3+GTD3tcnz+1+TlEmKYxCvaFEcNC3arN/cFylx9ZXOeJ5qnqVukPLD/1rzIs91IPMO2
4Ih0zYcAtvM8sF6NcUDOLOzgHn7O3SZkszG31qBbNk8ppecUPfVtU52tq3x5Oadt35jJF7ECGBsA
tVHABOUaBowUiSpZVQFKHeNkqbW/eSoS6hwkNrNOsTJZJhlQicgcgYrrPddNk5hwPYjQ4AZ/u6Nq
XYaikmQYjjvPOuXJQv5gNpKnUkrJh4ifkxAoqvN5jQGPfrFtdrzn9rO3520xcgUbF4PSOo0Mrbsg
JuFUJ4f2qSGl+3Qf6PUqAXvV3Rn1Om+/O6J01dvGuadIEeQkn4vuPiIhNQlboLg1NGkFCv/YVq8I
xmAVFHF30mRoO9h52PcZH8wwEDvV0b3hsv9nbxC3xp/IF1lt3oD8rlWcwAOFJGPCRK+ei1vW8JQ2
3/dSuhe8+jDJefao7FD97eQNKAz3fvkwJoZ4ZonUymWkKdzSfzIMXI3obLC0Kz0KVgmmrDwwNeLr
+EiYXOSCo94LEu0YV4d3i99tA337VyNQdl2gbMvlI3QUOb5QclW94KkBedsn8WOuQ+TWs/OVKrFV
NeW+2XhCQ2sk4zLLvtkMNzhxpahnZ0aiIJEQdBhF/pUw+sSSF/zk8ivut0zCtoBjNUVhJRPAvRaL
4YrzHeOIfJEkOuydOb9tEojQIxxZRi7w5Kw5m8osgHDqZQqbbnOAhIeEJOOAU9OMN95eO7iIRRCf
cNr3BWWMBmQL/TB8+Zk+jN8o3pHXz/lqWgv8qznqGL1bAHV9iZQueaHrH7qqJBkl8XlW+P0bXDpC
B098q/yOSnzfWNXcqcEJo5S6peoo4DK7hlqpbfBlFtqokJSn2R3Quz1hWlwEzl8ClVq3EDLma2c+
rbpGMMjIx2Wcl5afxe1z5j2ytAUEUCH2Ec8x4GDkogO2Ek/h56EQJ+K7vRXmxtceIJdELzWKmBRD
G3+xods2Pb1jLO6r2McGmeweRye63iWEj9JCTCqa9IHcT/sc+BPguQHtnhyoUsUoVnC4a49zSG5P
iHK+xDz87UGgrp2hpg4XmTEb80C+KeU0O4etAaoQ9LHaBXFr/58/M0rlMb3MogkssI03NjfJneTW
CIi07b3eeexsFpfoe/WR6ekKbZcoRysr0pZoESPlxvkicsBej5saIVVwmhxirt3dgH1HAXPAfgKi
Nlij3k3yuVaNsqJzWamIFIq+UL/P8qXaVvS5FTqCbaw7nlMtla6YfXpRxynPDGHrczq52shUrmyQ
90yIWkqYL8nL1TWC8Zg+6tbW6GslSw+tCpXgd1eBkPlqb6jMFPQzwgBSh98HVn8w8fHX3z2ncYnm
lHox/S9a9UGtbq5dzz1mo2W8+r8fUZfT3sU3wok/xzLV5Tz+O4JcwxMbe7IEn4vtlYn0shjJHFUX
QtnTlMDQMZbuI4wM9ki0EfZ4XdNQrp7eFuEjMjp4WnElGJvsn2YnukZOuA5OYuHJoqi0ClgVOsOT
abZMd8+8DESFBwTmjVlGRMT2QLjhPR/xu1kuCNMq8WD729T0ZSUIbk1NRLAHBRtZZ8BrMdfj0Sq9
8QB6JFn4SBbMpsTZR6SzBKABYOnMckMYINyJrXzJywcpFNA5fcFeM09WKd9Qm2dQgLc2owYhpTG2
kmkt0CsoQVDTF4clKpeKkA2qDXP6emdcWHEaBDy5UNDTKfbapuReFcPT2N7t+k3D/safUoE5Ndfz
zRB7QpGJcFEJNDWI+Eo/5ezSk25CqVscyWJo+Ms3mimjyF0KvcA22OIiXazhD1TLB9+lFnx7vFuh
HRbYD23KuPmXfBHoqyeF/lT3644xCccyjFdMSEakVVNMpE5+myFy3lNzIYzIvwgbbrkKEwzTjP4I
5SYRHMgBXoj+n+zsxkxweLPeP7r4IX6nbs7c0YwjMSS31I+rC9maKlZHF7g48uZgvZPTkae7TWDr
Lzhbnua3Ux1kdSRwfSO263lsMAUqIkRt7a7Bu0gcP3hmCjzF5JEnFQ5YDB12jPo2Oft5VQOkTC8k
Wnjq1yDF4+9LVndS80BqOSs43MwzGkPN3u4/+TC1ZieACpSFY8JQrO5q1KCDQGMaG7nkMDxnqbEn
hMStNEZ5zYQLc9zx0s2S9Zyn+I6/yaF/2x+Y6yeu9UZZIcBMVkaBGdUWygmRu89NI4/UxtR6oj+T
xrFEYTmm32cwrJoz8CH5IVMxLgQnGuaJ45zLzLuX8GogYOgLdhTTIxKFvg25iAK0XElprASbeiDP
LrNhKVLUCUIsET4/Lkgtu7ofKKRxRUUtpYtAJA++FNK6qTs0vSZHB7iXa8LD67aQCZ/4k/5uQ6LH
ZjQhBQ8qQZOT0d1bkV54kuKAX4VjMn/lJgsTgtTy9/7aBIcyRyVADG3WWaad9H9xjnRJ/MmccFDv
Ji3E1y9sQnqSYKKHAv8T9NiAplB6u6oThsm/EI0YekB133MKjoCUAyrWR5lV4JkrOnQrkFbCjqcz
PASKiA9bwb3U2H1uUaRc9FTfQhOG2+rZ4BbHjaAaU8uh6eeVz+mHy/ORS6y4nJ2f32dQPZpdnMKa
XG7LTzFM4aZpjIq9/4OWrnEd5x7UAlVzcy/mVq5bXUfw9SL1tN7c6LvPOsUzC5tgG+eNbTk5oCAt
i2Nj/GkIE9zlzcBuAtswd7NOXs7ohAkLwhL5RgAzeGTOS4eehs/uDHWlY9dfUmhZJtxjmXEQ8ODp
E0q1bl+akVS8mHVVaOdbjhZNN9PXyU4kHftDP/ARxZWqKB54UNyOpfIZ3Puwa3vwPfm/Du4lHc7r
9mjeTzD1exLtzzMz6mOfOfhyOgG+YzdTPcYtbPfaBfjP43xRtA5cR0koQeXYgcBejumyeCZqmZEk
0JU20sigaZPdtRYEnDOMeLlOvdpf3Sw8hvDYmOzhnrhrhoptXsmF6cTv6iN4M/YH4Tm1GN1W1Whi
soNvXkFPTY+pkJVPJhegXc00gTHOuKumY5h5XlVsxxgZQHIJwtV9N/XvhbA2V8eZewiL791d0CgM
dLfe0rxvGAjW5xw2GHOc5mmf6s9BU0gOhRiWNeyvyxGNok6HaoRN4HACWnYwjQbBi0j0dR/YYN7S
5oAAnNrnpizHCeM7va8g4NwgaQLds7z3ecvS3C/Aa5OOKtQu6LRdo5bBFA2nOzrVbeWRqmNhJuv3
THACGp2zJ2h5dxmfledJpax2CknamN3g1JmDZG4sUL9+f90jxi5W3KUcMMfGAJk56kSZDgQjh4+a
3s/znn6Qpn8DHeWSg8SCJntwU1VuoP1zhU3DwXananHkCEJtEDEsFfLGmZpIWRPUOk5z78cepsXF
pDknrJ5M/aF8LVxojtn/3RWG5Rsx7ZeoJM/EVY32q3GdKA/pAQ7B1Qb8YBXoAENNwAjwzOxxJSnT
VmlQPVhCZtxVG8Xby8DlL0zVsOllLzRu5RhgjnUrXecUDxio9ogvbZUPI3o2R5DhqAa/ueqvDF3l
dqjb/DNyd/KccsJMNRJL/FpDqHauhaIC7CBp1kJFh/9JE3YMzXM/H7qIDn5vAqpNy8RlxMZDOX4M
ExlP/Ar75OT0qQNintDsHb8+JylIGlKMXHmCqQDRdVDKtnzmXTUbFS/RVLYiewVi3Icirs43EvPL
0AAVjI+4/zMwi7zfp83xhhdcTSEgbajoKJhZiNYZb7Q5U/7Uy/tFDX4aOWYia2SZg+5JDunwijtB
tWP38QuuRMy7fIqECKwBrsHoEcHFVB1RzUPNJacXub7rEGIZcGNdvOHQjYqLPWuHW9r4nQcbolXJ
n9CAaIYU6LFKfak59ttDX8QHgHvR+/bE9fzceGWGElZJ7JuUZjo98YvwugJS4/ubpncn3r+t2in4
jujF6S60dajAyY5pVzx38CI9JLJH4sZKDvH+yoNnlcH+As0+xaR9He7PG0GeMU0gHG7NuMDgQdev
BLRg6xLnbaIiwg3rvtsK8ffq+xgi+8lZSojwB/nSvbS0mt1NZ0DkcXtyd/WW5WPm0rpGiieEAIqX
FP4qt3h1PRUn6Df/xxZjbOJo0UBhvT8RqGQ7jrscFIN+++zIgMbVXhdTFiQAki/aAFPRvvdfMAsS
WWkfWXRNn8B/m0xwCkjjZ9S+WDlIhH47yp0S1a5DZBFphgt7IAZeMbXuzZoNMXnM+FRUBruVKbLB
x+s5d8uAqH3xPuDkWbE8xi4t6yuFPMbBYPbUpadsF8I5WIvou0y+55j6heZ28VFeXIpmZ/HG7N4q
fHWlRVoBpFWtlnqE++OjGowTaUCU2p16O9LHuXLN/PDnz2667+mtFsgAvvAkV5gYBjAluiaYs/vI
o4CtLP4nXxzFkrdUbTYWGNHbARAsbokdVufVpUjf+ClDIuzgfVm/c8nxiV2iKIAgzAMa6okeICTj
fBjB8t4fTZV3r1GpHsRF/9sydJG5pR0YsjMmLRvw6bhskBuzehF9b2qzuHaQHQkALhY6V8p8EOYV
t94y4KLIMUq13mThImVZODZUdiE8zvAXSvAoCtxeAvEyuQ3XplgjvLHATNltnb93/TAequSJiZJk
oatBifkgY5QZi/0iOcVT+gI0iSlvQ7oAK6XxPVChApdbp1ZL0d6TYO3B2rOIZIuPb+7v+t2B2uqA
imW/mNx/KMvHVkDG4ay3b/S6LFcF5HMSnr4Pl9u1g9lbNiNFpHgDy9Vkph+/IuZ3qvSzarasWv/6
OARPYJrjKNZ0qBtMIdsejdJHzWbgO9WIiNCO+dP4F+9U+S5MWH2cHdliNkLSqBcOGoYjKkdt5/3r
tvqpIh3nu1j8a5wjPI7frr+dLd21QGLP7DARy/xeIyMc8CWSWU38QvMG8XvZELt1MJ3pga3Bk2zQ
iu8LOtq1Cj4ycoVFlz842PAt2C4Bdb8svyrIjtWiNyj2khG8Bf4Ee6kZ60phttTQE+9JxsoYnKN+
te3c02hMRTrmVPYpToUOnixuUBDfl3+1/cIwa+26vZODpQ3pxpdft9Fc2I/0F0jQmHmtUZb/KgN7
Yru9P5fVy2lwqjbkHH3iNMRqunrjjMmtWdwKM7im7rbNZvHOcE2ZCUeXQ/253Z5Wc79V3khjX8C0
/ba6//8ui22eMUnxX5PMLXiPseqY+T8UvETAUzqLmrcdnRs4HLh5dLM1HwIYfWLZOjyaCbW3gCo/
aZvfUUVbnSKxAEeSsz8uvLeHWKggcDzkBSA0S4mxG/yJzYjl3Rn3JY/KkwczUnHij2KvdYs35JJM
1/IXLIqwsWDGC8UZ62RtRg4z33d9lc36YYHx2vTk7ji5wtH8r36uiQgrb2EFPByjQ7+RAcmmENAi
afO9s2olhAfHoHjTewrbkjOFY1NTGBJpQuyWm1Iv/LGl+8cB4POmravDGz3zRtdPPjgVxEy2bQml
Vdtrcr+n/ufCSQMZFfbZgrVIRm6kBdYvwpsjFxpagCVTByS8wl/P7vYe1Plz5MRg0n2J42LgRGL5
xPXu+yOO/uaRXU09zvgLdh01Tl7uPVOCgUZquaGB0kSM5TEAetVSN11nYWvfVWeNxSeG8w0uADKY
TIrHnNmXfB6ytov6iDCvJP34qKkKBU6CY9DJtmQW5nJQWgFFAmffgPg956LtxbJWrXZ2n7d/x2a2
vm+c2BRxVaMmIqnUTaPu4sg1bATajPNPfcmv+Her6ePuDuseNPAb0Kjl0e7n6iRXQB9egE+QDd4D
kZoHgUsffIsJrzZruEXbzNhl6b3W5othcniDRQLe+AQumdfA+HjlTnYPWOhCWUJxC5JBmB3cmtaY
JxmyAiHICeLS5Tyh0+Xmp9lHu2xXqc3CnRjJF4Meq8LXpEp8/Uem0T7Dwfqb8tVxMyJ8e72Tltz0
iztDuO3M6ezcEtKmnzC7PKHnpWs6vgB7UgdPyJdt65UWPQ2XQazynphCc/8+97dMqzUdajRECWly
YeC76h6x5j+HexLBZVFrHaIHVfqc6+tm9XL7GzcwbRvTaLYimdS8E+ZW7w+ZwRCa+2yz5b5rtxE6
fxrA5pr6O/dY/NXgEsQc7ZAX6Ggv2K5zhQB0/BANZs7uWFtyMzus7qbn7AWN3KP5OpHwh6ovPgD+
1iIpXUeLxMJxLn+i1hQQbxYFpXdfO/wSXxpYAxKeiInNo5fCDkKH+hGKwLz40oCu8JfgssMMydIQ
cI/VVeim6SEeifuyd4wnpWnkQ1JjXW0yGPo2PM/YitdIeuySuSs/ZYy7yIkVdq60ORXfyrOxjvPR
UVl3uGsx9HS/7PIioZVRCGA/sW8Z5UV5Bc0LqvGBvjXVUfVcC4vnlyga+h8G+PHXB2wjgngRmOfg
nZd3ZPDLAoRZBdAX1nxUVf6SUlk+nvst0D1eEfcHOe2Jfkmiep5Ai8JEbIGe8qY+tP5DhUSEwqpy
J/6og4i4pinT+pPo/c74gsAUB9CBp/DcrFte4YvJiLGFy65fTbIqaENiW5+7bgusQN59VA+x5Ccd
8S9wunJB/JDCOt603fpssmLuppP0wNsWXVg8oa2AakvKXU6C0M8rj7Joet7CZ1CDY0IROMkTp0be
Ua6fFY9ul/Glsa7bI2VfjZxQ9y6fbUMZjEh+OJece4LUH+zDjzcDFpcZYbKF7/zVbzNNS4hEmGBq
EfAf/nxDqj8Qdo+rUswhtOA9Y8xCFOacpVyWt99cw+rzg5+38vx4uGmDmae7/i0+qxbkB5EVMJpc
bD+bmNZS9WtBxSzTqSJZX8gfe6E0zu+lcLb5rwR+9w4QXT23zRNglPz/B+I6YVvMluy3Q+lCNE5B
xK8cf5JUc558Z0zC3B/vB0rFB8BkaEP8kXldglXpKPpYhw7OnWnaIOBGfauM3zbQRrDGnb2+WqkW
w9mHm+9IwFU7nlPQIVa1Mc9/dayyVWIXXUQZBIFzftimN6srnoDcBmT9MNzDf2KOFerwOccR2XRY
vlgqii2qcwnVWssCuzcjf1yzMOdcnz0xwNvTZmO/jNlJn2pUOOfXAZdnnV1O295qSvsd6Bf/1cpT
N595oHS5MKGAutibeuGmvmI5TfR8RKk51tXtFDWNHUOwqFr7M2Cu7mc9Cq/DEzQ9yM5KjQWnRJ5n
emt8fNSL973PYkBGd89hqqTA7Wem6oPXFG3w5to+1fUoUwJzsgJeRXCSQ1xQWPXDKZjm2j47n2wU
DxtyMVmIpg1UYqFGC+kS4EfpcWotS93a/VBak93EFyTIqwiewjtLlyMNhbd3s5vp+wmag88/mxUt
RQIN6i0tq/9Uwtw9Oc64ENJHy33YETgXZ0AbZiBOMZYMeau3Q5g+1k1nf3Q0uO1yuFZnlT2TpOH7
1CHZL80FNZszW45CMpz3597QyhMi1/+cqlf+W6JSfbquDgO06ADs3e8jTe5Vo4bO8wtxTqIk5X7J
9nObSnL+6uD3iDbfzEZzpO1x9CtPMT2lo1pIFj0nfVhnQSJG6G3y+8DPV2I5F5MSkPmk0bwwE3W7
SNQsXyCQp4MoKGiTj+NCBVz7pMr7J+qfSceGDR+/WDvLRYiabcPHUTnMsQUxLdT7WelsaB1d2wlY
BvsaW5+apX9MxFJYhsgpGUWutpjlx9YZLvzBDH9HQGz7bHuRiUsqOq5iEz+eJ3hPXgTtGocrCelq
FDQj7roeuVBMG4tSL32nPkBLodvH/A9AKg74CCKHoYPiDNwvb4BYcIs9cLZ6TnZIl+aRDeYnlgYx
4qHzcV5IqXPYIQ9pf4PtspT/3wQHG4fCWxuGbRblYXI9oGcBdIOO2fURORm/P/4rdM/mCAgxSYbW
hX5HGK+IJgxkKGz1zKWsQe4+q9M6kobdLHan68ex1Jk+/f8+6DPveALZGS64RkN3zeVzqdttDMdp
Gsm7D+pS+xBTLpZ10swOdYwXnf4q0repGPDf3ZDgNohuDfgEDdNWVFGLn9Tgr8bbePkNk8Ki1rQo
sRdWM80tpJ4sH1u4rmPcGSRN+2h2Mi/s2VuglgPtEi1IRpzc/Ui/CjAOQYFEwuyDVEAM5PQIDNdc
yeIUYdXQ/THhP/BUpt6Eau8bmE5CbKb5vrVXK/xHU0weuoWqQWd1ufuKVRsKR3IttQNURBz6vDDx
AlZAiSVhOBLwa7Qc9dEmu99zsSdtXrhIk9TSbUGRpNAMqsDhf9SzD81NxamDzpEje/XrtJ3r/0vx
mqM0PPoeKfENQz59K15+vCFb3/ENPMNzrVq+eYWZoBNF+L6ZwuxSWXMktgqwE9bTEfZw0n/r1KAN
4ksYyI/ekViueoza9/529uvuUIrdSsN16nAgDMXzYB4Rs9Jhj1AMRsbEz9QgxNsrnokGNOy9D3e9
kOLrv0C93cOf98YiALRRjiCH6zoKqB8gmjg9hv92E1LW6MKwyEpqWidApbvpGJ4VigCBS9aGV9a2
d3v4Gjrdg7rXGRV+B08wCT+yeCyMbQtrb1Un38lcqqVD7z0b52FN54g/XihQrO/jqZEGnWVi71Fz
rj3AEvIyO7cBiXkV0QCTxXiPud6orElbR1N58IC+lsGKqPAhtTdw0k/+E4f3LPBE3zSDu3uQ60h2
hJ+ljZCI45OHUXM+2lluSM7z/QujBz8AXMHv9/bvPN1VRfXx/3YNMrkLyQgm1p6Tl38nqckeWqfD
0UA+aeyrMVaGGrg4ZkcWwZltWLdwKDxLB51S7gkg3WjT4jME2PZYF4x7MJ0B4QYb+pM9A1oTAE6/
aDLd/cE0cxvxyoeHNY1rdiJj1Fnw9brr9XZvVVWLDDbPlZ2ygHUQXV/LeSaD3aOLlRud9EhHaOOK
RoMir9uLlvuYzeJB5fuquqUgaXg8IAzU9rcGBt6P1tXXr0WMMYasv9TpjA30h+mOWWL9oxK7YFQF
0axnI8730cLWr/skCi2fh1oCJqvSDKF0bRZHm5lY3jI0ZfkVXP3DRbSihXZnzYXAXi/SAqkBFMXT
A3PtImktKCUZxBGd//xhsFpgL7E5PY1VuLfjXoq+dgv8fg3KMwkLTV74uZxHCGrq2tWrckYSNc1C
B4ij4mTWlif+pJUM+V+Uo6GIXT5whR6+l69EZ84ulX4f1dp1NrCj773WWKkbRf29NUpeHGUb8GPF
Apz/HFuJ3JdGy1SP7MTQsfDw4f/ut9JRkQ51r+Dmg54rV70KSubO2ySPi3p+giu22y5wBq3YQ7p8
geyjmh4M9ko7IlWHCvI2bfjUQwhKtWEvyw7ZSxsDwQw56B4Yu/oa3ORekA1s+s/83kjFQ1XXejj6
Gq7HHePTdQDB69qCwnZxQHjyXMsMBdoIMVUYcbNGG/S+W7QxvZswW4q+I94oSmAjZyB4UgMHr/4N
19UHbFYBirqTfDa8Nuq25d/lMGo88koXASPJ/d3yDWGx9bPAVjifFn2O55a0aKNJW6iUKGa7Tg/K
vQ9X8QLsEZSyuCTyoMKJDZky+ee/Chu0UXzH87sD5wLibpK9BEAY3J/KanBsMoJV/ntk94GlFk+P
1bRHalY1EsDhVBmcez5bEHgBmE3N/NMjkx8hVEp5SgsSsPwljyMhdpjoXJr3wT44HwWYDdXoyET+
YBMRQ2xtsREnsf1ayaZ2YvaW2+fkrl94GGpRL8hEPgk4Iqc6zB81gPth7CYAu7eOF+h0ZuOJpNwR
Nvm9axA53kYGnKWIPcPSdNrsa99+o650PlOzENU8yfyS6mQHbTrNZTvZxVVGhidjMVxQGolGSWL8
AqqICIijSb9zIAXXFese/ShWpHkDpMRiam1eFg3DlpTg64cw3XAjewIkqcXIeoSiIqjjjK/mdQyU
zykJtWx90a4YjcGw6i9OZREDDXhha903k+lYSPdGIPGZYnYA6H9L4SBYQ5l35cqusf8aIFVc85+R
vMzxxl/YX9Oyj7QoEL50rUbnmIW26B67FqDssS08bQ+EXGPwurfPrVGsgcc6hVxGrAlEAG28qQHk
t3pUSseq+NxSIu4k1uHBJYW4M/xy9GxUdUyjHYRj1JqGyjW3xtfLPkRtLNCRoe/ufK5UKzlSIPvO
ggryyO4mI9dtwgn10BJ5ITpMeAPf6bhqokBWekLMIUbWxNSXocNN+UrgYdprgSXVPnTS579cgBBr
4VyY8mhcbMVENs9DxUxI4P67GsqLdYa8lbfFoRFG9znaImrlg/TC6Wbv8qL+DHbXYDUStnWULWxI
i5We1ZRhhRlDKx5pnvnQoeA6blI3W/IsN7fwKW3/zHHiyBDf1Y3TOYT46wMGYWoywgGnCgoa0Vpp
uvzY3QS//cy8WEJn8WzSP6P3PRkSvkjLs7Z0Z8IlrAxA8T8l3oVfwr3cOYTOiHW/MSoYS9qz5k4g
1GqynEKJ8WKbKNdkMrhRZXy58jCNXJY2J7xGut8vBk0nlI8ywnIXboY9C556NjQ12vtWtPMckDSt
gjvmN1fwmHIcLs/QTlMJSZs3BpiSCAGkIEBWdOtuxzT0zURciOCxa4ijF8L+H81qqtan7NQr4HMY
9qoyJOjjYsXfPCSb+i7oTqivBKq+6lalpGNMceDPiLdq/becsGZhVGSpk924HMsW28ZDpZl4GhQY
khAvr7oEmby0EwEnfb/itmsWFBLS1uC5AjeHXZ9GCzKBniWMsR0kdT/4rSk8Pp/W5d7oyTP7dFEw
0lyY74LhD6js42oO4NWHzjK4ep9jLyM9xTxna4IxYA10MRnpxWZtV+xvrjTVnC3+ypZTx0oresba
leXiNiI3yTs2W/i8XX18nkIAfu4SC9vTw/5iPw5GrRrZfxqNpsE+DQxnriYFTYZJ85Q4BoIo0Zsf
m6CE3nz5O8vQn6t9DOY9QF6oQNQ5mZ3y70UqQTIfIt6myDXH8BUToSYsahF4LYfY3duHuzAQTuhu
mjj4TXYusOvNCtdqGGkhw38TgGicNK6SePoVxlhBbL8mkbIPsuZNPcPzpwmD00zPtnUincwcTzcV
2W1BS0QnbRlN2txLiCIeBPW37z6m9C+dckXsDJj8JeYLX0KMF/5m7YQN2+yVLdHR8kMrIEiLol8K
iI7/NpaovFrx4hX0uD06TKbnVaqDShhXmgWBwd9c18jCmyhBe5jQhnKW/zbg/H0yHqMzj4Sdrulf
jRYGAVGNK6GIRBl7wmY7tqoAW5TK8J6HH5YvxP7U0bVuXuHuioqE8slMvXJyUML6rbDE46T2gsLp
Ox+uJXdG9NQaMgMPVux9UhTdvTJMz4qWmlBsn4kuXUHiuhYffqyORtDli1oLafa+2PEOwSp9PIYk
LKGKbOJ5fLqWYwZ/7IgbBDL1d9zeo3rsNe9Rqby8hiGOmPh3luFGbvRnFn1MOYyoA/yMgubU2RGm
mycNs6D7O6BR1Yd9inbCe3di0dUd0QXlFBdNwTjjMnKIByYMIaqn8kbR7f+MpXLijO3a76l4L8YP
um+Q1s/VlHwi+9CxoPnsQJOk8QHzv0h1khAjLM9f2eJUlnRmT95ywfcrazl5UU/xjhQ3cS4BrjrK
Hv0n+LoZqD6CPnB9kllBbkJ5B15c1sV3c1+IzeDjZu3JkVYp7VyZlxDPJcybwME5wpOeHKf5r5Jq
amd7q6tPGaP57E2oxbfWnExVnatwc2cdo59YIWtdzCP3zUw+GS1kn8RH1dczHZ7eT4shQhPOPyce
iqwzBbkWLXo5zQW4z+OqUidMLAgB2koKi0vkYlP6zTkGgInG83wm6x/db3/bfjwWWPkO/d7Q9v+W
l+04nDmIb5hTjB9EkDSCw+83KC/gCkAQJUnE3KlIAGY/drJgnYrMuAFH0LzNBbzwvohw4YvRB6am
Z4ixf4LxdShuIoD5kzwb6F4Tfjuq2K7Uozv84Tz6OzY9R1Sqnml/FxF46qa2zI93++WLkbRbuH9k
8VfudFoX8VqdXX0qVaJNmazNdI/UFgCURM4ToPSOjMujQCM/3XoRxJWR5Px+/QrVRJ04Lv6sRSUz
eBli5d33rHSrsZHBMRaYVVy1FFrsu5TnkU3VzaVTqEbj/KBkw+WS0dyUfBAM088EDjHZ4cqHbDt+
c2ZL58PV/JsYc54QUmAs/tf2zSSZkc9YwjmOVgdOcT9VQV76LTw0bMSaxSdbPXt8aUqr8R362bmC
03iocPppxhRT8B46GQgiuVCJ/vImyJGm8CUQmm+DtZzM3gSWBmZbXHjU9VbnwwGwTTFsMhMZa27y
q3jF0W1JD+AJe9fU93E6YuarQMV1yLdbY/7jn6iY5qr6piUuFEgYkn4KDuDZ9bkUBovCuCmdlJzB
uWFhaO7H9lQBHtlXGM+O4SVErcQ7ln8qt083ALpn0g/5ZF0Oph/m2f0rffKErjtADYeEsWUs3v0C
6N+AJ57xk5TArVFePsvddNLuA2uiBG5xzTOZTzY+8i+6L2xGi71UcZ3ou0id4A4OOm4dpZ2INZB1
nGcbUScn6i4XIykPOzhf14Mi3hBoatF7EINCAu+9n4F6cQlpYgVpVZ4wQfyU7PtXytfW6+DSkgK4
Mf1bIo6H5GFRUHB4NhAazTOm9+Kq85O+jmBNTQ93jeJ9+OzQduLz/9ryH5o+Kpy2XIaY+rx301Zh
ARA9+pG/os6WJbnU6tmuBbqkyqiJyHe+lZw52ukgV+DCN1wjkyWWCuDSSIY/b4ApjrAysJbT2TD3
954w9QEJhzfMhGGh4NlBNuZrOkKN+Xu7ugRqXY3qckHdjgDBsD03pkN8oNuSynLEpTmh02rwAt9y
CgNuQ/xG/eU/0/w9SKUEQIdrNjiC2KjGElOHdRYOt59sd/M36rS5SomYsY2QH++CJxvBS/T5eAaK
mkWkArTDrojulot7xsfLfNeNtA7seZ68XeB1iR68jMV8Uor1f1CYa8QI3qL0gf1H4cIqxt3qTn10
3P/dxfrNMX1mPeNM6F1xLMsiSoazK2/sFk5MToitP1CA6JFTnQ5FuH8oNk/fKk2gtcGqT7UTDAnr
F8e618NRJlqB+/ZihrcSh9RlEfm/fX7aPiNklMedIR3WImP/0eIblTCgr+Oh0t5cLQVUBQm6e/aB
NlDoAlfMvvEMPjOkGw1bBFHfchVpVaJGWebXURtolZOkk08n8kJU1Mw2cZ5iVm1oIZhCVPRXpHBI
u13YMTuLo2S7VCLvsfMa3gqyJEX1UeTOhum1mHwEFXfjynnbsc3tUnPiSXB9qWhIOxTqfTR772Tw
dI6MTElptJddGlC8q9w0uB25AgH8tkDScoAIsPEEMFrIKQdf4zIPiJC9zzmD2fmMPUGShrDYps1i
EUdapJGDGNDT6njXSR2+HcFMO9Ju0DgVIb/T2yO0fIE+ctoqBzYOO/6NhgRkq1tqh7tmaB7+W7Jf
Lrir6qm3jqLCshWLSqCC45FdFChTuP9Gf+hGaatvmo48nNZSzf/PWNld7EcWZ4tV2fzCOTqHMTFG
NZvOD+9vH4igJ3B9HjtfNC7IUGmudRDnC7xjDHnq/2BkF9RACTKZstSkVFGuchQoLBqPTbF9lDo0
QP8ZnxW7VjDhWh3RXKAeakzj+ZjK/dAFvtJYMIRiCLrsYxxejdmExX3QHBEqfQYtaBXWcgymPZTj
ipH7nQMaIlYkVokhB8xKewSBN6SkhL66A4ozl2aDRuILmmuuwXHI2P2rvZuqOYzT3qyQzAABbUOc
I9bvIZtjJ60FsXdyw41ysFu9+x/cQY3wX58r7SwKnrt3QqbxzDj12E2IKJ663A3EWO/+f8yzpbqI
DOS+IP4a/qiop1+n1VJxyyS6mRjiRsmUfvfQBu+eSl/SK2fCWjU4mHH0qLNKaQ8zBtZXJB66bOF6
QAURQteI2D/9lZlBi2igJOmIg843dQIYc9f4x32JtIeRI86NOshOzlEecQm8XUL8IVHoYqOGZUsB
tAlv20w4r+SpSBk5bldrxRLD+nHzhovvtvvUGqHjmx69In8FkH/h/p6j1dVMV1od2SnAs8IwlBLR
LGDUuq81XbbdgTeQenpRkf/5Zy50p8N9EjuNx8etaKeUJTIlUkfA87KTjI6QjVaS2SBo1BzKa2IO
3GVtDkwYsSoM3zhKrjH6xgaCgwNUjkP2qcqP4rH2KV+UBQBBpCAYLr+FZAbOVFHVMnUt6AWl3DU8
5MgHJ8WsJTlBJxWfwZJVecFECQebVe6nVIDvenQOreGnGXAtOeBOMgfO7KO74lGAqe0b5RJSrF5C
fx9e5MrvwDb77lQzoFYnsRgruEyRCDTbybLoBgCorJiwPcfHdUHKcuIJf7UG9E4zGMbFnEBPMylf
mm94AP5S8/AlIqYBQ3+X+cg6MOc1MZ9xmRD+h8/rfsK3VAM0hyy0dkpXG7gKdFhEm/+BBCJVeUQa
w1uw6DIr1thW5DlfCgknWZMG1grDHvU0JT4sGHBDEOTVTbbNOtU02UGjG/KMJpF+nAEha77PSjUH
4UERZlbuoaWJ0a7g6GACIswOP7awPZdiv09Im/Wh8IcW6G0x0lmmAQr+zPtvanRIGDuPtzOBQbO/
3Dtou9H7xt770zoTqUpB2CSaOVsu8guljmFNh8k9Nq19j00Wgpyj3UYZZiFzAjc9Oxn1xoVy3Jq8
kl6+r4nwdZsQp6b6MeqG3ClFxiZXxofoM9BTRpPL0fk4HPDaX/y51aRYtAEc0k1hXVBSGYBhYnqI
Y2JTLpTPrspKnkdxWCpjUWvz3rEPCqqG+5F4ahOgC41zl/TELlh4FkXjuCi3mqtdtB6cOf2TzR3N
rABsq/RpNyyAc0FBH9au9Mc5WUBTsuV4PSKR1xnlRhsmLYi7torKZpQur0A5nVYO5nEz0pdBhmta
S025xEmedf3UKbQcTAZuACKkWUj6cfpE3Y8ujU5p6QwPet8/O42qUutUOArmshPb7XOELJQO1bdO
KkU5H1cKhD5AOzjm4S+7BZSOx26Q4yjnNOT3gBycCBbItU+pjJoQkzhnMDtzLtVnCST/tCO+A556
0HEV7n1cUQLQpsIObI7pMZQUr/13E4IqYQW+MiRHlhztmGA1NvP76NCNc3uoPe25v7qGTpZVV0oT
fo39pSONa27NiFGGhTKcD4KA71IYLcssqsNLzNTgkYkRtnUZb/i1VMe14LbaCexWkc5ce6tidjTl
Hvn4Jeu3TUdQgUdrd69pIMiNcSJeLWkejZ6d8dEAStD9TMXxQiFmLPFonrr0dwyJKH+zsQE2RGDV
Rjsghjbd+PoX8rHwYnXVb2akRflmYeBZQCoMC/9lWZp49/AGRIYwpRj+g3rxS45S50kMDjbOrp/Z
1f0/CKBERJCYht0qlw+pQU7SXpJLztNBlQfxDTWbtyhZ3bERQNeCFg5rpEgvr0s5dBsdm2dbRbPY
+0hKg5RY+UOl3pcdX1JSJWVUfFnXZgcSKTNCyD+uIT4sPbzan8YpfKL4lgqvOv7t2xHKdShBhZ7p
2Gb7CVOZlTSOrRUm4/6f+bCpzVDx2AJCfro7l3dDWMlEMkf0V4+T9RFhuPTt/zK8bW9pa9F01lZk
3FlOprjoOW7xp26wi9iluJlkALEbOfmr63FstPGQJD8unyTkQzKwWyuHuEmaZhC7J2zByQGdHIT8
/yP6Z2W8lZLvaX6UQw59Va09F/SbxWzJKYW6WrnsgCnVTa9K0SdKSZUCahMt4JTYPtU6JnPG4r6V
gYfX87CRqcQmACgyFk4mLgk5Jd3dGwF/DojHQLJoWs7H74Ykb1JUXkJ7pQOL3sUPoiQJvdq2Y5dJ
zmVks9HU2x/Vpmrn1GdwVWnJ+8PmjSHHvAXO0fo4W7VlJfPjR3GhydcigxvLkCQho4zpUZl/1Wac
zAj54wYVIvyUmVH5gVBIBQ4CVSS0j1T+aqpaZGUbXFwdJgl+XAHQk8KElJiHz392YD2UliK+vXmF
rVkPbSieGDK7Hyi2gU02M5rRdSXEfsQqZmEV+K9X71U/nUAOECmwSGGMDH/4/ffPgOBpUQDmIVWk
KEXsdgbfHCwQUD/ZRq6jJQXnyRn6pSN+AYbbRCJC+S4OdZv863WBq0i/VAWkh67XcK11Tjs7M5Tl
bUYluQrtRD+zgh2Hkmg7QtVSi9w0UYgi/J3Ez4kOG/HodwUl2rQ+w6+fdiZ3PxtQrUTmamJ6j+9b
8LAErRNha8GmAJXJL3V1dh9vA8gWG2JIC54Cjtnh4IyukkZvRiJLx7Weu4WKvqA5FDIs4eO9iyDQ
ZGN2V9s4nCoT5O3ZpLtoSng1cMyFVEuRFvra6rL9XhFbWhgEga2S3A1YTCC5Z9JNxnkdjk414IFY
oSDiPJHwe/PvA5vvG3+YX2ArJy7z67425EKofdvm9GcpSPR2gnXll2e7TuvWIvqBBS8XInxib62Q
ofjTK6bK6SWQ5aQAMHUi+t4hBir8nmoeXhuANh7gS3IV4QiCDRi5Dpr8OUZGbDikKMryNMlkKMZb
lRbEVX8MPs7+7gu9KRvpAe6gvK8DjBjZYU/wzm4GA2C5wQ+lEMlvjmkkw2y4mE35ywoeitw/M+nG
8KWsZx+GG5Sfhpb6DM0zGgwXAdH8ctrYttyo2yWoVFVDpviJYmX/p8XWKvOAjKuo+M9QuvfOl126
XDT8XSmkJbvXiITMCyajf6gwgNbWDi2NlrT2X6bCqJTjCF/LNxiiZKOdZC19f+oZJo788vAkyY2D
OMftZ9D4G++npynLhHPPb8fGsvlhn4HKjsju82qCjVIuvGUbTDUJodQvqc7rWyES7nlWLs5dure4
lbsf/08Zcgnc+aFsnKB+Ly8rd3djeTmZRwr8JJnDp3XjT52KIe1+LfQ92Cpf2o0W8UEAsd7Y2sDD
Pv568G976tbn3F/Y7vFmfOdpqd47okDItxFFKv4JfnCraaWsfFiUh21gpVwgT9Royhz94GubOBn4
c2EvFuk1JF1tVv1wQBxp8Q47QZGqFKo9yk9afeCEnCGESjoorI46sh+jlstb3vdtm9gzbFD2oJmg
MtMLWYu/2iSMixE+gpgSphYncHFcUoVIUKESCSpLfKmNlqZX62IIGAyN9lA4WTd9g3xY5Ru7cHyD
5af1aM5+vulSes41BJS1Wf+MLU+CuwTnj23Lq4H55uoWbUnrwR5sjVZXg8FKjTmhQZYIDV2io3oN
rLLuro3C4Vruw1xNj9DTqum2E+gGOWgMFkG3AcajrdqA2wZtNnAzOEKEv4aQ2/ZnQ7zU0Qd0rrP6
K/QrPaeTmPTuz85Z9yakPb7JZj0T0By9wWuHmqjFLZcY4mTK4EKJRG4ZhEpOPdYQwKqpwHNb+P7o
nwewsAcrAOXqzJIqDlgsmpdpZiPdvILP5Rtd6QhrmSwaIh5vP4AszeZjMXFUObM66tupSnzfTyVp
N6+wQ/aizJrhYsNFgCc/T1dTEcR9EpAVqGjj52TFuZT1gkrFsdgsricMTTPPew6pSLB9QVr2oKFk
DMbGCK+5+2ROShkTkqt92KPQRkuoA0MPBtTjKNz11pSAZhWaQfiF8Z+eSRX0jEdiImALMEjQyjfC
8992BBotebKRPWbhJbhHXx5KveL2DxQM5pM1vgMb1DekeKvLRtyna43Rh/+GdozVwkQC/mVZJD0G
3F6eAMi0o8Iesz9pWR1eXVBsD9iWcJVjJlcywWkQJON/wYVDrylMmyn5vXkEDH5ZqlVFd47VKADY
f605U1ccIq7X1qoY3X2LzBlgt9Sx1Vor8ijCwHm1DCee3IIU+iXEDQyPPKg+ixMaS2D2l0LfnP81
S6PBJexbV+vPtEr7noVper74XyWoNS6QzPax0aBY1bC0O30BVU/RZCXVwkkt57l/cmYgIgwKylxu
0NkrVgUYWs/gMySV79CVv99WDSIYAsW/PWjJHJmQIJVE3qZFHE5L9tkGlCE/ozBdQLqxV6H2aELq
aojvYH1DNjowRQVTsdGVWKY3PitmpFIMzRHGh/kaSWtWCiyuFnkO7AMMZFPHj3TmYuiePgVjcmbQ
EwNoXhQfukPEfqNxSkFUATSLH8idoTpJdWJtt+846EVvP3M79NrU4gPNMrT/k7exn3vg5eEiP5vG
zggtG42xNdGCt/AnRqd6F5l/ZssIzHZUkdyRswAt2PQzeFNahDVv75txa2tEZZFzKLyBZMG/qF3l
xhLWEtIqYteK5CT9ymaJFew7Kqk629irXqtsi8fblxa5h63z7SRpZkGVRaoiAwWHR15g/FnxnbI6
whr+/VnwGbZ+7dVnUjixjeJSQyAUpUDqJn3gqVCp0w/RSP6gYkZmHK88DFiDnkl7SbtQ12nYu0/H
kVIc214ild959OyVdNLtRJnv12dSgWkIFXhzE2Q9iDmXCPGFioFFZAq05v0uvXlRMUxQhnr9IYCB
ub+xu97T2CnLuJosePliGrNF66YpGJzsWHrFC0+/B6yJESX8O5ZjHjBoaglMg4NYeQpPpg1bNIC6
vt106jgv4eZ9+/5QJCrKXjgi/4j0DRkmxKbq752O0Q96hi+vOgFJT2W2G76DW1vEDhL5BdWSv/wT
7W/ahttZeSqj1u1V2gwt/hpvTJs6FnJfzeckpOQmBUrIQs186tMp1LGeTiy9GP9TcYJtY36NC3X4
r3BLq65oDk/ZtqDIhjdBx/GR57aIOKxX+zlq8RuiVdWpRlTrdYlcH8cICceJGa8ZzOa8TFI47UQ2
WWmmLaAIrmz1mb/fNMxT7sZ1hwz0v50aUpeO8vD39VQyoLzPt8l4MyAqlZI1m/cMiBZOL7R7eCGp
dyPEq6ELIJhopSmkVxRGdu8TAJ59tz3pgGL4eNiT6Zqhj9d2kRIu7CioIqBn2Sf8d3VLybWHi3tb
hHAjIaZIqZ8zYpxpwoFog8vJMN3h4GobOMUpGZSHa0DUd4dOgYQyTYik5O9XPvUAuZ4bSaIqVk3Z
5d+80IVtB5KJ/yRGHjHnj+AvTjofkb2s6UOtQmSYkIiVfu00m9y/TyzA6WKVg/MH1ohbWGnu4fxR
rTbl71N3n0LKUPQ1A6t99w9Kd2WSl6+ePG9QUXK8ILgKKTO0Ud5jx9psKdGbZKmP2oZF9pdgoJoD
us5poVH9BME08CPgh5S+4ZXM0HAIXnPBwsZtXxR2RirkZqyjGYbVPHmte+oGIXgopwsNJJA70JEF
Iq2KiC4u/iMJZHQFraG5rYv86U8GhYNX4/H5QjYWCZzULd6xyDHfPvN5FavSpIiTOpa8sx9EKpCR
Fhaoqh2zRBxyOsv32sEpLSJm3imWqfcYPsiFi27wloKT/fjdR8Lqty0TWPrr5wRxRPxgFGJskKa7
xrKT1Kl8TXsvsEstwUv5hqWPunscsRmZvOADs9Y4q3MofghlhdZg1izy0WrnFZH2DJqUvl5W0V8x
0zPjRtMYMX4tQNZMAbWE/rmHW63FOLSw/ErJUuq0UflJ0SgUstPnLASVvi5gQuqJjOLXhHQTINV2
K9h3NQEy9xkLBG3H8Btg11J9h4wFmUZ9D9lPoTnT1wkSfU/u8OnL1fDtvZUWNv62lcUDzAZgc5D9
HUkUmk5cScM8bqLRjGnrjZmzRAPa8rixOefklhfIkN592XVYHN/qPsz1SlD3e0STynfUUF1/rwbX
wcKXb6uPstYH4vixWOasgg8NrXNDLT8EphpT7OFkKjPu3ql1MC0NqcXLr72phiIVcikKE/uxxC1X
2YPUvrdgGFt1bmELU4C4zasdsEsTIBO2QDkBoZYDaH9aFBTVfhR5Jc5ebH9yD+cGktuVtuhaJo5t
LB6JbRrYgfVuXc2KhEESzrPBu0Uyto8OUqY8KM0zXQ1yqGtoABsb82CSidVrqMo5uZoTMXUXmUzm
CBNhJHFJ76GTnZ4lmjl76OjvBa1M+u6yzfPQg+isH/gY3kK4rvekjmy0gh2VgI7FZrxzi08C9S7T
jTI83NhRz2Hb84f3KQf9hAtt/9ucjkiyoUSDsPahEpK6kB7YQcu5ojMB3w8z9gdYzvLOOJv7gIqW
TBWYwxgs235lGjOLD0y8+YGtWYQUPFVPosE5E0u3H4OqbtFlJbUXbyIqULUUGAczKEz67wtlK1wd
tqFTmhjmN43FmkBy7ltsU0mKJHDOzDxrKVMnsq7Vccko/KYVzsjbZ395vvbPjJ88NdRjfbroH9ca
oAaNhWMiWdu//9H039Fe9iJatnYk8D0V4SBWFBStky0lgWyLWQsPI+jJ49M4KxP+w9Uvgl8dqmB+
L8NJWcUOEosFcKfW43vB0IBaaXV9m/8giTVdU68C0hb9Q8eQS2T3QygwZrP5HlBFnsaIPL9JG9+8
MyQ0YYa1FFH5upjqR/acHbQT5t40viiOApTHr9jKbvP+VQs8cmxD/VFgbqSzinRyNr3JIAyGxDye
Ik1QTfYKAdCpKe3Z6j4TqMgq5gywGU67gDitUmu+LVjfqqs1AubVUCuLcc8jDtrFWfZshcI5hRLk
XrHwElq2KVJw8DLGLzA7pdQ/oV7Rv2G3jZg24KgyhRSxZPAq3D8r3DPKIb9GbiWv1FM899pmJToT
RUGA4XPV9VH88yAwHJ7K48qCn79mzXOvwcRWitCZYMi/54pd2GF7Kg0zNKf3fPIFqogqmKvNClWk
9VqaG4dWFcFvqwT/4wwCiUg0ulD4MW+SMeRW40RAWqJVu4nk4DQeKPUhd3oXOAMc3USRwnjvABuN
z/FrgSllKQpHgU7ZA4jWlpw5hn6tlXr4XvgGgt9JVkVIikQLQZOmm51OEzJa67oRRvGhKUqqyTZ3
ouIRC1MZc1Mj0g6xvXmt57O3d1UFFeJ5Fg1FGwzYOKV3hZVRUJ4fjBll5DX0R12U6JNHA8f7p257
p92XwAn8kuQ0e5pb1GCv/djg7pA/7n7L+Vd3EMKq1HORhJzlXWF77jN/WDUhKfwjwKFZZn5oVSYD
zNVONX3gprIgJ2wIY7rBQJO7WVrP2yyIhxbqfdiXe08MrlofZcelL41kYN9JEdNKaLqZ/U8zoJJv
rkPC/UMhEdTroXN7HumTz0bATsPUUUUJOZj6vhKCp1rFvIlPPyrxGqDbCXudcZFaMVm5igtIufBB
UldEgGMXZx9eHjfAa7tnOq36+ArwFvnGrGXJricgiYC8yM41FjcddnLyKWVoACqO5qKNQwvMQwcE
f1LbPNS+HTjYD1Rkggr5bOW550QXb5JGyUGfKggvKmOAmF1XSKXLljGnBbxwwZmXoIuv17pWw4ea
TgpcEaVbjE9+B367RwM4f5CsA0tyI745S6ImpYHBtNYIPM2BWod/+bAxXceSnTI4vkn0q6xhHkCz
VEptYboXaL4UWZrCnZGPwNj6ZDdum9JMNUSryhCBHhQhm2PwfHmAFvtXG4jG9g48b90dA+p+oUh+
RRfw9plQtDHGWL4RuTPZW181ZRr4OTkaOhB5a4D3t6OirM/AiSiE86V0luMk0HEX4Kp2IfICJQtS
8KRvUT/D4EAFOAQvumvO3e+tmBy9t7WddLoov0cInxhmwMlCrM6LzGf4VHInEtwccBTRYTsXB+Js
dKBL/+fV7n8BJaopUPbBaI5gc9Bvr8ctMMqKwo9GNglpTHMMrvCYKE4f3iDv1DDXlkKKC0FNhyOh
9Za6H6+PlHL0bQyknoo0hNo7vUZqJF8SmIpKPGPPYWR1UwWCjpZXW6kXb5AONHO+w/8oRcTaba+m
qpm37i6KCcaTq/oNjyDxJUPhnqG+Do9xQhkdiv/YvR8ZdTtp+w2FQikME9oMmvPF8yLmshBmjkIM
wYirmUe8x2plwHJPEv/sh4zJuJ0MsLZwucyeZ3ODfQaqrJ4vN83jcjLdI17qiIuxEyb6pvQvjhIB
n/lOTc42pfafXm81zwSdRtdC2d9WbltaNvJq8qDsgY6+GSaRCH20Ih6y4GdxEub3ZUJQ+0lipUx9
pSBTB0hU1zduc2SpEnaHJYywJmYtTqUYTKM4pJnpErAy86qeKElyfB4sE1ag0+QZOUTTNkvQOOEt
5mlpemswCAO3/pzEM/FyfJxyIaG+vSdnv47cagea4rfcSVCgOULwW/pE9MPKzxo64zM5AigP2WVm
2KZKsVm14g2uInR8aux/x0Kvep7fujwSuQysVdHjHrb0J7T2LPsWBxd8JIQe6hdkd5ib4ozbXOqu
WXETLAgjqPiqXH6iVcTZBUa/EL17lZnpkx8UsfEXGFB40yHwPQOsado7EV6x8fraTtkhaB60G4dt
YKM8nYPMpstWcqbXqOoiJDxwGcIk4InJ5fJAKBS0y4xkiLA04sIzrvxGDsgI/db4JqpJLp8wIFGi
fuIanqmeSJHXfFLgYmSnyABAAITGJ/8DFzJkdy0CeVKO3j+ZgAfHsyf59a4/OPD+WqO6qVVh73Dl
JazXfPthgXWMdrpgjQveokDRXtnAOJ7zWpIvoRqQje3cre4KbVYGiUb8A0NC7GtdaGsmEn7P0YNk
6MFvLYr7VZC62c3xhrtIsL78f+67QvleOUCM/kYvS+uxOXAoB2CuyL4ZygvkinGOGxvcDrgI+/RS
wsioic3Rv/7fEAc61iTxD7Ysq2jxohDP1Guwtd9qONkyDK+N7Pey+y5zkDoaWPT9j4ewcNQy7VgX
IWLk2Ra8c8h73UvEbEmmfmdNRLuSuvjTBgDXKlBG/kjOm8+EVwMb+Ab6q2dJ8dDQrmHGpnDi/1fI
U7IDOlBlP8bac7XCNPTpUcquhImYjIwAC108YlaGnpCvxFq1Ck+goNYTV7AhTc1S7FJYubzmOWcr
15UY7+TEQJ26Ppy6xwlIGJV66+Ixe4PWBIWo4hxvb2gZGs0PIdljGG3KpLGAXt0M+03+EF1oki2B
550keV0yssxi6WnCs6gUyij/WHJSTTu/UYygcv/RE+jWgnUc1G6utLw5Po0eaaDWWTnLTqupupf6
iUAUK9Mvy1dXKuA1FJ41cHoV/kB+8f4FtsLjZOMbarAoj0+VVlTppb7QGnkCUKDbMd5JrbdknZKv
J0wRSXCkAFDEo6a1y5JXx6ZHomWFXrbbKU83suaMz/OsxyohSUFKkHnVWwCClNqEoOKNLEoh41+A
XcnPGoeR5EsHWRDmD9o/kdn3QfY5OXhqQZDimQ+6qLwBi7jLDubr/OhdLzakJwxkx5qSlmIj/pyC
eRWZsAgvXhB8DNcZB/q0MG0BZMhwIEB6ObLUIqq2BdEpJmD9RwR/nXTrBVh5B668ZQDTRQIuE1qS
hnltL7uWZyh3dLU3rM3f0olCS0oR77ICOLdR+zRp1np2kcpK/Y1dwgSQ+6Bkkrqe7wCtTH7QK75t
hkc+q1xTyYcKKlEA4a68Aej3DJB5hK85CVSQRac1FdXVNioleH1sJKrHTotPdC4JfLfHCMB4Tn12
W2CyfZYPmwtL8qw0U57nfDWVDdZylwjakTk5MuIzKpLQkHJGAUZuUfG5CiKIQxHV+nfo1Ozfc9WX
4JuAY/mOXbGsjSEhIUkOoePukBijIP0GRiJQyVocjIro8DSmC6P/lMlHH6UtmFxZ8EybPgweP6bp
DRZmDM/TKPpj9Gi+jPwHlmSSKKajBJA/jTwAxRLjukKj8YN5NhF9O05Qc34l2JMxP1ZKA0Y7yV6G
qr61tDFnlyEFRCdbo4Y9o4VSlv4YmNB4hUCGzHpGSaihBICDCaPXe1hpF+cmb8jK2zL7w+yzzmYz
3KS1bzEtUbTFOdnBqoh6c/MSXCohpxdiZZE4IqgI6I6x2t/zU0BzNAbDQ6T9p/IbgnMTSZJQRaNC
JTU2mWall6v3u+urTB5EPDBJbBeiQmV5yPp+zi82K/pooUUmgDQ+ujalqmpjkKKUx6JigpwNVJoI
R98MICP5N85+hb7UD77cYQNIEqIxGZswte1+PxoLAY4I1FfdJfkx0wbjpeYcy7rdQ+iMGeyb1xAP
azX/BLHe5Yf3mAvAfUwFlkTk0AJj4YhpxGuanVcvJGgDNTKz5yeZEHIiKEsacQrGtPy5vdDT2JlS
O+SzoStGGsmwruPmfuKUrQ6rzZGNz8PI+34UluAShdgdUyt5s2dA9qrocqqHemyHLhtQT6h2yt5F
3gl8lNEwarCjC/J7moQUZFh6UQtVoda+33BsOtl8V2CHUnBsKQ0SBd8UTDPRcQwPLkZ/cmJdjmZG
Bsv//S6uhUfGqJIewC38d0jadw3oK6qIZ1hEHglTP/TI7aOLunp/Vyy+GOmIu2zms8xDEDfapF+V
G7D0pQny0hBiTQnmeOFCW38Oh22FwnCtEEZt1DjnXTSUb5IPIWNnX99nbngL95m66MIJ7nkF/jM4
T2MIoixsZZ2NYzMD++mwVIGVPfcxRiLna8xDNUrEuJSyZXFusq6xYta1kPRDI0OIfR119NZFifqx
omhkP9NEEpdGIW5EigIAAAve6MGA8HzQZ9fUghum+2TDDGqzOW5UVAq80Vqq23buIVn+ENgG7vpF
ABgLfWa8PEXKHwh9mZyQsPr6cAncEAisYjl4kCVUyxg5+mnhlaV1kmzJ1jS7L1dRwdyMR3zMjhz7
aVvg9Kz0ilsY4xD776J6sypKBX4MExuxw6uKWWPkGpSVrCEbQvGocj7lMHKSZSv4ASuo4BQH/iTR
6OxG7YVswupDEBnEFM20C/PDdCLeAGqEM8PC1bHZH6ALAkD87FsEC5sHUJ//amYE2Re+fSXOviyp
Vy4y10U0EQ0umpAoFGW0ou+9esYaHe0TrQGxYIOXjCLhW5Lrh+wEL6RFlZOJSt18pjIg00lAbesF
JA2bxfJziqFIGZKE52wf00OPmDGIjwB8ZWn4/7m0WEtArgP60TduurOihPiH3va17f0eZSIr7Hjz
XXHQqcj17OVe4OjvBdFD6Lxdou1y1G5y2SGJ/6b+U9sWXnqvdemPV5AJ9cZQ51RRXlrliQz1rT97
VYOuwdiolqqP04tPMRcnXF0t3mrd3eJbwxFtrA31V9VhWRgoTInf05nPn8eUpMzzEG3JeOAiCIXn
PzM7lp/tJVosgygwIUFRdQ9ZOa0pBTmu17rpmS6OoOHVhSWo9YleJ0JxoPR1xiKqgoutj4oWJhLU
a4iJ8GGrzht5WdIidC0NHor79sxhf/zcFYYXKtZ9+mpZ+YNMvN6YRbVZz5+03dw8vBqLchVNyGK/
9n9vFdZuzF+TLLummy3NUtefYRR8r5ztRXgFhm9MDEApBOZSe62MC8Qalf0duemP13KBpINe/0cw
A3NNuVbzDi09BZ4Utff5FhbXaqhCMTQLSZ0D4TJ2NHdCND6E9LuSBo9G09BCvsOb/AhXDSOzXU2H
D0MHlXsHIXzsFgs1qMzo2LyZCwschzXbcvXrfBVMzBjDkdA/fdEjlW4RJFYozKmF0ExF5W+Jiq/W
RpTCK5aIFoXhNmDRh67FqE0w0wmnjDNXH8c0q1MuwZIk9AjC9+tJ0RjNRMQp0uQ3FVrfx09r2q0n
Pcvagtk2dB8144ZGVXckq2+agqXiD/rPALDsyXnHypZyQN2eBLDWosfQ20R4w6jD3R0ipMiNaEwL
FNdrflHrEViJln0c9IResfUQiAv1S4QfwsZHWlzorWInm92ISB/JSdw9I6u2p0u4yb0ad/tKVEaC
FFyRsC1zr5kEG6GFYsBpLgS3NGZgPNEGUkYlWLKkWSzNA67pXaBnJz5pVFrS/MrP4A4xiXpjnVX7
yWMFariLvjZvn7oDXToLNrITQcrFgQdqvUBFdfrwb3qJfDCEIFRk3vOkDXoNx8IS86ZNNr5yRacB
7IGomUbnuY0KF6y5H2bGT8zVRb2gTr1dIGs6+qbp1vdfTGxPwBHJhP1TxCJYW1cMuTErPr0EWlBl
QiHJ0mJjCJCn8wRPIeNGvASWUricQMevOCHqzriL6weXL4ZekVSVRQY4bdXdjAckEjUfJ59tURZV
8Vbu0/fBfIBR1mMEJwS381Yf+dE3dNCb/nNF8yooYgvREw+34Xl8Mk1JcymkS+sJRQGoSGiRldv1
yvHl+5f8IMfg+77VnW71wZz/JeG+szixeMxbiZ8+YV3WFm5y/NSEIvByUHWuBdg52dD7oTQfstA4
YEHd6QNYKFdHox6foxUuIYzZlkyoPomiFYwktkJMRAJHF0t0VwYMPaULtUuEdMAYDa4tscyIJNBz
j4VUqplg4v4DmQpf/1yrLq38ESfMam9naYHSDFVbtNfX5Lvnu8/8LiJF5C1d48uJF0o2YMQDJYg8
WGFmu5xX75fYC/2DMPWl/atKOh+0MVRbSM16HItLWmqozELuwxB0PxxavjTiGnP/pmeUJAt0MzhB
lYM6w8m1gPzpseraQVSU+nWXdXN9YmG/QwzawUS8XQlkeOQGBAqcL2YBWCpKr/S51kOuaWXjxRSv
ehq9/SjOqjMV/j/dGRhsygT1xj9VKKvLXRo9tD+wRYn8xPJ1A5rs1tjJSXWru97QAzoFlj1QPiVH
7Hshji0ZQiqBnD+tQbXMp+g4XZhD0/377QdKUcA8GXneTVc71Ffz7yP1W3LEGxCvOaowOegiNQsW
Y8nUEL/T7XIby72spCwMxPr3fcbaILG2f2/tgDCry6JNtgZT/f1OEWuhAiwwdMyx9yQXLQPTQCu1
bGb4URG1HBqLTt7ve9V+9iGILyFdThHkDnOi/eGHXg052GE6UD3s+Eaq4Xu8EF25WiMOxBkMiwJs
ZRBqQ+ZT19y9X47g2Oomuj4qWMMRWRjJqJEd7jip9aPx6zwqKdSTeFLGY8kiSJcO4v5WD+yC3tVN
sDfZVMVM68o4snlS/ChlQ+7L1o0o8GulsirhShU811C29g5GfMrcLqgNDe+LHw5K9I2uCuWpAF5Q
3jajo0maG0C/0lexTm+HeaPzkfMYtZHVr84r3TCQE2u3CBuGsBIl0Pt3c7kjxqep4lTEevLiF7WX
/X/gDgQb62kRvTaOZFxN17D7nVG0yf421KIwyehLWgn9XF1Ivtsj4tOEg+8kWyRNC0gJFFv9MiKE
WMrL6V4wbFzouAdpREiJY/PjrfVQTEwpWzyCJJFa8B20lShtcU16u1Uo5HaHhsclfzHemlu5kQNF
HWVVur4NWh3BrWeFLOeoKSfgsP/yBpEWSUyQqtpLHOpn3GDL8tPDpaHkqAhN553dtfowpI5rw67H
XM0UkiHV05QwtVW5FARbA3sX8tnUhx5TYWE27kF2pAXFuBN27wrbHb/l9SwcR7cxqj8qoTkE/q3Q
J4/uS2UhKPcKYvUszzvy4pD6gIqnZYiq0I2GlRbTK1srZ2TNTsfYfkznW+6lKkNrU/+f3aYfGXc9
VLoSge6QITxu884dxTw4fmFvk9ns4mnyUCd3XDRmEumQbOrKBIkbDE0XI0ul6S4PMow087xQVtDd
ucY0T/nHVvOPBPzrPE5SfHvXERVUfaeBbL9Q61a05pzYs8bSvX0jINtjeA8SVa2nragnUd1Q+xf1
+2UsiXqbQfR6I9Yy/fulxgWt0dTGIgjozsEy2VJasn7NASGodWPQpvDstBcYiGxwYwRtfE2139kq
zoh4u2tyywwfbICO2suNXStC9NmQcdObuYbc84vprf1FbAALsHqik4n6r6QW7O56Do+596F11KTV
vj4qf8eyX/pE7f9Rv2iNBBw+kjgvWrVLOGU0s6YR1PYxRZbHXkAnrTZRWu0SdWTqR5kg2XcVN9oc
Vu2/PWT2IRq2RpcHE2rPuWgCTvzeivTlIZHnFI8FgF0BS/+6sfuHkW1ZOeLzgGXWrY5T6gI2fjyn
x98sN0LorjJO5JPw1XzlZXLRMpqnYzr7RcM5KaCNtLDyi36MwzgfCGF4E4gqV3RB9icSeBHmdpr2
m1BAToS8ucNyRIxexyZGn9p8dRyuYE2W4hjGaZ4IM14aOOgtRRl4d9bwWB76uKVOiajWN5o94gyq
4ytYRLmRIMPqO7WovTgW9EL+AHMzRujSia/o+K3rbgMyzZpdi1Y/PoNHiJNX6RvXZk1Cs0a7w07i
ZAthppiyxYZxv2qB68vNqhjyO5nAXzOKrmFmIDhuiDQD/i0IZYinXZ/9Ob8x8hj0SCR5aUC8dvkF
OiRlpe8XC1Ht0R6FbKJYflgIJgzbZdtI48SuM+oLxo+S8tDvC0C7nMDW61igihUwTmACrfkmqdsb
oe+oCcsEVvfQuM95VdGTh6Uwe2mBu99NzvApnF8tKm+bZJBvH3vlPGHDHfEK1JaItgl3FoTWRPL1
6TdmwZ9wJ3vgFiAqu6drC+Qyr7ooPXiIpkUZ7jDKhz8wbM8jmTupMRDqBq4IDbgEhuzLUhEygy21
QFtul31r83MU32ynkKSdNQfXnJky0MyS1EBNthWRGgXCho6VODKyGnrKYXTcfnPZNuaEsrWHIrlv
adm/bDjb+4p59UubACw/irTKdAXHJlQmjuaK97u4lNQEYv11WxzgqDyHlxTn8nGyaT+bNCdTyTpp
2rLhO/gmiOHxKu2WXCESH9922XfXfPGNIDMqlNJwKlVyuLluEpuiXoknE5hrWgPIINHWsjeXyqax
uoaCH5iWF5xuwNMKuZhOP74aP+A9ijQ+hGRehWcZJUzbT4otBDZvlvUW50gbsl0msPxcwFISo7JY
NTGZVhGw/db9mAafr0nwhtoCVnOj4OSIlcYE5jvCIpqj9df10sxxiBCEqDs/3ejtQMKa8zpqURBB
DOV1hRXzAXNRLgm9rlzUqFTS6vqSTPOMXy/E4jlljcL8RkhpJAWYmuscBkpdnk6M+1LGxQYj+Irh
y/7bUZSXo0+8zhJ+C/mbFgyR+58ypx6xM764zvMTHGmmtJKPUqdI9ykKhSPak8A/GEomF5/nALnZ
ceWqFlDTzcLCkl1v3K4XOx3lme809qPNZgK4eugYvknZXlTJUN4YIiXm86ElG60J+6X7YAgBH9i0
E7Yg85/zA/qdOp43KIndr5JdkT7b01KTf52rVsAghIa3yNirEQwmrs34fGbzjUu8C4FNcYhmcbzP
vzMjhNCZXEh30Kr1b9wuObfBygHM8N58lxX8NjEj7z3f9u0r/Fwor3gpk3MtWWBtfNUNUxxLxM+E
ngh4+yZjQezA3FZpIxAqhkbnrtZCSNyOHt5KSUBgyQQgtelsW2W2lEX2WoyxUEcjxXuM8pHIji43
3UuEqUcOhaDFBNyQUBYwq3dG53fRNyd2T46OcuKEAY+SjLoPsDwHcPkgHv/dMU8pK+BmERXP38QG
4+harauBlUtFLhQDHxzH3u/s27AtAv0DFlAdMPEgR4Dn8coM6+tCd9BIxVlVZKh9JV3dE5zaphya
01gh8fVBCFbuYvuCZbPIdKA6X9fDkCYJdYC5Vv52ic4LiieOdc/VHss1R1wJdWjfuE4jcEX4RSsp
OmmbBWhEgpDO3MZvtvIhS19whKAzxlQsK7OSeOyDpRFzn3AxI06DkX3L8nvYqR3ecq3htNotmzF0
ycbs1KmMnDZ87FRYyhWy9Tt2zpkVOoi965BSVfsilZdtqEdfXxdVzvpsjCxVu4fWV8zFX9osducm
p0nERfB7PWkmJ7TI3oU+LXnjKBN/4f0VPGeso9aXr9Q1vBbUbffoEhZUuQdtjbH8pC/gtF/X2/5u
cGeFxnm1wDSWDpAXaJCUm126YvpISKOJ/dJOQ/MKT7zjkiSgbUHoJaKKvOw3sJld5JhUHiB0Q5YD
Rb3/pCcaTVuYm+e6bIW2H8LQ0hB+oGIN4RN2OWkMWRXEMWZiOHan4BaHsak+lW5gIQLhiEOWmRhZ
RED7cQvZl/eTpH+NlxTZ24WVlbJQ4CrXPfXUzMvi9h+B95xB08N0AM1Se9SVATzrFidOpFUu+1JC
Dni3hTAepUIe7FzXHfZML7YyWiV2ZRUUxZhb8mx/fsFcPOTbI412UAX+t8G1NKduoCAvvHEYoOk/
09iaOizozrWTJKXrMX368By67gVk1TBjHV2/RiXHHRUPCjRBTmO/f5Q2ZIv6zQtM8XyJt9aV5ow1
Nad6awBPluQdjAEqYBSc+z4yJy3d7Vr+qrumQm5Uebqkiw5/sHlij1/e20S0dfrSlIcsnriBzj32
H25c9yO0/B4ijAPNioulcxPWgnPz4ZhoHMVtWcdlp4w5ZaV+wwO4wDCLSfIl3GO4x927SJaQpFSc
bM7/q96758bd99uuJ152A3/tYp0ka+9FZtfmBlXoHOXtZ/DvzUhjzqRYwrLazzJYEzvahCBj2g7x
7dhpgvUNSV26YDbIam26x3CGA/YAyWndwsrCVQz/s9GLi8Jz5cYiwHJTFyCmuClNXa5BvHaK5R6m
b8k/n+bdn5P2MYXaBvUNMqBMXqi+pXbtbXd2J72LQ3rpqfAhCoEQyP5DrVzqABWSZtPKRUbUkLi9
47P/0U7TCyJ8ijYu6JJ6MdeECkLUxCz+3tTeWYZUGt9ukZHCepRCz/XUgt2s7ZV+kWhsi9sxgL5y
//E/uYWnwPxoxARB21oB3HTw3Sw87NM0OGmqHlsa9W+0u0rG2oIZtk5iSqsrUhHoQlRh31k+cRzx
HhrQsJeE+DEtSLtjdNyQSbZ3w54z+EMY7WL/CXPBpMloHbrvJIj8wateFVSdNtG6T8GloQJtr/Hi
zmLfrxRAiC2BmTNwlK/GUMiPeS+0CPSpZYjAM8Cz94AFWqdYjQepLeuaahL5vk0SlIS8yd4HcIcc
4r81cf6hWjB2fdTL6U4BfQrW3rugNlvrlIg6yGme8GNZQBiZOrR7Gh77MdLqb1++eALvcmwiLxuO
pFA1COpH7hJI4RM73AlKuv9Cv+pdbQpDMYtgvf6JFYqu8bCnsyCr+6Ez9rf6GWsnIXkrIXG1FmuA
zNJQ1WdEastI04EtNVkrsa4F0R+NsvD4gmIfaDgllOg48VhB770VHogUS9Hjt7Jbe/vqfeBLEHVy
C11aYBsVApB79HPZl2+Lt9FhitJmAo4g86DgwAtJwEy0GDbjSV6bmcIekBemeYKvib4spm+RTjsN
/2hJerIEDiouKH15phzsxUYlnj5Tw4+84uEiN/PdRpAatt47IUM5XmJmWoRqAlkfug8Uc7ppZmaM
SPauYt+hrTH5H2S5yPq01LlDKTmWNqP/kZlgrQZLQLbHSZrJNIhJdxnJ1/CGL1nmSOKp8xlGsY4g
GUldbR9SpFvb1Dso8/pz+sTQ9M/aG1xJzCcNw4KdcJFVapzODN79sGvvW/Hgdoi9ZiDoN3InDfwU
ZHq1XADkhCWStQ/RFjQV1U0/EHInLrS88kPXfNq1mvhKY4iuFDqiuT0r09E/LGtd+xqplBEbGJJl
zQiIzSleIqh3n5554HBjSHKBcU0fIxUkyq9aVDUyvXGzifJESgsbCgsUgbl+UxXguNzA4yIUfeGb
fwYhBFee7064069/jM7447WHCKvTf7uC6HKrXJFw1DuhhbCBy8C1SYGRTvQ5zvApazbuvRw56g7T
5A4l6izLh7luzOxtn05fBxqU9swjndfLerEFfMtiwPN6m987Y27E/Z2mVa8zno6XnOSM31eWqTF6
fpH3pDa+XLTIOPEWYRlQWJ/zTYrMwSTTlFKSxbcR6oF8OoUQv27nQb4w5V5MLxmczgfEDeayH1o0
KvJmq/MRZQNEdVo/xOmfJYZRbLOZkawk9p5zY1f6JoL9kNgCJYc7da5Vk5N63OJ0zLBSny6hDfgd
7MgmGrDDgXnALqtNdm4yvECROCwitiGGgxTH00utpY7k4ee1DhIS0Q7kYmjtI4w5UZp8bVAMvNYO
d0ln4h2ZRKKLIgIx+gj6QjADrIvlDGnNByFEEGPzzmqPt6hVjQRC19gmk2PjbBi0wjrhaVecW9fI
G36ePHk9RzOGyxzSwoZZQAfv3iW8MFsh1CnyisEJiV2b8M6xnJunJRTO8J/E9ITGUneRcMRgXwrN
wyPAn0u0Rcxan4qcv9OmF2BUMrDHOwRIGsyTY5v95dEBdINtYSHmcMk1kjSArsbwNEVjoE6Hwpjq
D83t7D3SITL0+mHb+zm8a5FJS+3jccO7ARU6jW2r1OkVAkNUYUHmKKMHfXevE7tv8t6Bp7xygmGW
lEauEwfFxvFvOc2bjwMczJnLkhkOHssy3LkWaH0xnpiU/grLGwuR/hBWUdcBWZQnR4CNwu5WDaQz
cPMKWf5CpILAmhLzK+ucgEsTqTARjrJetFVK0U5UgeiQmy0kUYmXU+6eBg0vfcdeDfBO4UJV1yMw
OMP3jkimn79kYrU563AGw9TPGiwy6PTVmUkRKcl9PvI17an0HGhOmA5JXgx93eZr6ZnYyDLkWOm0
MlI0KBhS/Z5jfYqFL6SQCqdPejzr/DEXBvqciBZwRc8z6VLX3rB7IqK3uod/KU5+qdc+hqQBI3/q
tHQ4X5bEVNDlZ8nk5ElqpHJ/X86R6sqT4713/fmHoGSJ1wQ5Y52QoUyfnXxW1ZJhegsGbwD5dHiS
eqotjC55qO3x2rlg8Q4CQQkVw4uoFWakw70wezNPpl78Nc8s/CAsvSlamvkJrJ+iK+Q1p5Fwb89L
0EZT5bQ0ZDvsVAlbVk6jiG6HtzAvl7L5sGvdvprrYVNwR2zKRJsmCLBnYGDvjO2y1malP4tT57Wm
1OUi+RR1nEKDRqRiVV1grqBfkvoZb2nulUy/pY6gLpZT+q1qgJ3MiS58jtmeQr3WIgGfBsKcgtPy
+2p1eWgp2nn9ptlEFFq1don3qH5yS1zTOmD3nNjItMY8pubIOt+Nt5RMyC/N8W8BPGvIf21IJ1r9
UgBbage8+S+UtS84wACSoYt2pwchveZ+f8HPf4QvVX5ufb5LnnJvzBbsahswSPKQFGjdpGdz7IRg
rbXczZPvkxKZsfKHTNDfOwYq++O/A4Rid0qknnR0reM4B89ycO5wXXl7wO7uHA1OnEyJNWFoykEF
uCZHfAEEGFpRNHQPZyz4Rlkn9Xr0Uf0udS6OBhrN0Y8V0H95ehbPR+JsgQBzNWH5Dwlbtlg6sZWW
DlqlS9pqpwCc1gOrmJH0eYznO3WXaDYs9DV/R5/If+PX+y4oxZeiT3XukORcFwtm/I5KosWCoq7x
vVO9qr/2NxX3tzY5ohO2Xtu1OBgklbV/TInBN+HVz5Ub6zUuDLv+EMxr7+PCZlQWS3Mesa44EEn9
2rGHak0lRhNI9qymPDPyVElsFeY8cYw+7YHmL1IOE+Fzon9ixxnZOINNRan99EGOUbrjhTsPByx3
4uzCOnk/TJm9O4+mHHVbmUlrCY6XYXtADttry9mMsyXd2JCZ/W2QWYvfimNIdTyqmS/5HpfysrQ8
XSBF0vKry2zoDgT4Pebx9U+o6lxPdRrFQaMbPqhueCRl0LNNdeUgRYB8b8uXeJQrJe3aT4681/It
TWcjHAhehjygz2LlIZkJU+qqsYGckSHExg6bZL4pH5kLuI24t7WzPFgCv/rmGuskYPSz2HR7fptm
SM+aGJaVazkgv53RCmtVr2LzV1JTbNZgYfDF64gLlelXZ8CLUCVV3iMlTVt/fqu8XD872xzCMrDZ
laYx/HqEHs4+dgTttSYJnql590XT5Dd9Vwumyo8BSbkqXm2AHB5RdF2TSp+2ufcOme4c08jT42Pl
lLE+HMOZ120BFAHZXOCRwO8eCUXTFX1dvPMLydXQc4Irdn9XyITdLcHMrZy6iVpVh/ejh3/tIasL
afQSkfULk+cIE13296Kh2Izul8jLcplaIPsjGhQBfji2DtsIeQLW8pfKWBD0ZB3Vl+UVthcA9DHU
oE2oJ39EQOJuzCbbkK5Qq9liFjdDn2DlSBQjbHoaBjMa9S5LHG9ZtQGu8dLz1OkiCmTGfBQoKfEV
oLtlvy7l3kaQFR/6vqqfhZR2ocN9DTqgnwTXa3JiOva8iDsTv4ky4XI0QunSkBtF4sn7Rhqv6+ZL
mzRYNssUlnV9pEpDVs3CJq388ZbDtS1e1OK3Bxb8OZWaQll2Cx98t5yULIYxb8iZw5W0RHf4znA3
HhgKgtQ1OW3BWUVTgOVBgVnlTYSdueGno928rzNUJgprC48YX4+J0aDy+s8KZpwozBmN2tmFtWhc
zXVVBnFrAj5ZYP1w/oj/0LH5VagZrZ6W5YcVN53xjjYN40AapDEW/koNwKtFBjb34iobvTRipajp
6w1p+OCUEG5NiPfsdQTH2dnN76evVDgx3yWoYV1Z/NpTsFGM0zS41I+7Hn6EIwwzc4CVPTPTe+ZD
lQsrlkz9BftZ3u4bCTSrDseaBzB+qB+7fFxU3YSJEwg34fkbzUWkZ7Yf0KtNIShWgVrEKmaj0raV
ot4TZL+UW9zy1mCJ8ciBPGMSpL8rixKneXx0lTRe6taxrtzT7aoHXheKSVcpJ58Dgiw1Jd85WWhH
GQcqyAhAJNcmkHjou6V3optJCTAviDVR5DoWoH26PXaenU5W65GoK1UxKVWHTKIAfmRd0X+AD3Ix
H/1HPPXYcJT5N18qBngxy57SrF0ynr8R97u+DjsGuCramyFPpGgiDf1VSGcG51USQSgvJQUBUf3s
bH3jKqq8HHe30qdfF95YoxuCtLmUAld05AUvxCs/0sd6Yu9VbiFOS+I5bg6Ddg9NlxriMhO80qdS
XOYgl3mGdmRl3reD3ANfcrZcvmfVjXsIHVvV57h8AXNTQKxxyTbwWzcejoZF8XLyc4ZzKaCb0uaY
Tlc3q/PID7YxGmHz5VHSKcd89LxhPDp5Z8i1jUhj5VfLZ0Kjx8YCCbxfUYndkaaYPrZWxLXdAhMo
TR/pnpVlYbIlnaXk3vvjbxV8gFAAKnsnpcP4773zO48faJu9LOjA+wpAtCKv7/IurIt7rkMCrzQ9
3VdL2bZx5NkZfPTeYsk+MT24WAN8idTQ4pf2jEQVu6Z8gwFyNEEN68Q62ALqtSMyAiQyFjvUFiqn
/2iqKVV6tw22vGrxcK4uIfr5HXOxvcmA4pIuy9zOjly7qDQJg69rLQAzlDUTUYevZyr2acSEMOC8
mnYhGZzLbp+s9SkVYQtF7bi6pZilT4hFHA3H1a1DTMDQ6G+YpOO7m9oTl45ikU92fgpWj22hnbq+
eRNbvgwGk5EUakW+OddKJCNatxhbXrbvMo2AnhVNbn/Y3pQbfu2kNJ4XGZPUzkGAx0EPr/DQO8/G
oHgfRHu8JQ9wtipfuhJsQ8S2rJXwtgF09MudAjNpoqcWjhghGpJcpyyYJE3qpKf110gW3Ynfg4bx
up7kmQpKe2Pls7tMReP85nM/MScjtuVHt1cFTxXZvNcZDcNGcSN6Pa1LEaIa1OJ7EeKgg2y8oMDE
Y6iFOTCLH51tJjd3ejkBgiwCAgbVVRMY8KBqx+5pxSZxW/Zzicnb7Ht3yuRoEHkNSQXKHPX5hCpL
CedjP0cn34I4HcFhUD0/nSK7WVcbVIr07LUeY5z55OIksAp2m5EOdpBAdq2Cl5Z3llIq8We9CqbM
ieM126t57vUROHsTT+nYVZdJdjDq5gRReMCvZfK0aiEnpx01qYgI+W1i6KJVekaWdGMSS2knF+gX
Ymj0UKi/N6FNzt8Zg3qL6pw1THAi1iwcVdvsATBEvHTy2+V8OWWXAgnsWIbCERD0m794xVsnCmqq
ad3Ohe/CNuUM9KxXlaNLhAQOo6YbNaRw0Ou0NmXOjiiwX1dOgGSVDG9tj07w1ks0pA6PmvHlrFRa
MWNUQdNL2q8OWx3KXer1ZRIkvfFpD9+5/kja1WWw6mUorl8hkzSApTBca/cgYMaRoXJYmOhhXmnU
PrpjD4y2BlURZB0u+aQ+p8bfg9oKy6fEJh3yL2GgFknSVzXD92gXpKoWNaSSQv+K5HpEXUTVrgMD
KQ2YaMXHYtbGiptGJCshRdBuHvB2FcSRacIo6GcoH0vkliP1HDwt77mRBTBVw6Ft8Juhc6xlBEpP
TAbyLmhK10v5YozvkZ6pdMgdo2ny0XlrjUQYciUKI99RmXTByLOGw3sPxoja3phlfpYSZtnM0jqp
fMlce5qduAPan4tZiDWOH8bChX/p7F8xEh2a+bCcZX3iFHH6mi9FmRF6o2iSLEUJ6cLgOtRCLz6P
io+whjH+9LdygvPxLlOC6JOqGXMSdSqHWfRUoQbZC71VJbN08AtBjXhvLjpT7023+S1ZOlfSlzdY
vg3SloqAsVd3n7DWP/BRBDanwVaw4p02suBNBzLmncZSX2ZCTK4BG5tf2KKGJvQpFyp5ycMH3jgL
u/KFjDtji+aJdYoivpfkbrZ+mlVl/2FIQQKWQKl/hu9u0duuFJTnYfxXPVjPZPvimavN8FDpemJY
rg4mEqalpD011UTvZviIOcq0h1MFgYIpRysdkbnlZ9LD/lm3G3LojRUdVte6PClBHcJRAFV9T19y
OMaKyGkOiX/ResbimbZb9wT+GS/Y8U4lYD9RxrH71MV0uV67JVKEMEgYHt/9VNydJSrN6F8eq+Ri
P1dAWvZU+bYDuR6I/cRo8XbfwnxYRZa7C4h138T6e/RWft+LDh/fVnLVG0qD2ci5kcIms1Ly+OIq
EV96RKuOpMzbBLqXNnMx0HCLZgaLciIW6kvCdbsTFCH01N/dYThNhgUJf3WwzP0xfvRPtjsj+cHJ
/G4QD9yWOirg8aj+xdg1FkeSfXXKDifBAeQzVnI9RnBiQrY9mld0MzFvCedINAIGKmz/gD3sNjCZ
Xbq9vEdrgx9Ui8ksyMMJL2PVh5D2mnWhyEd9kJ5i5pTqZ2dcbf9O1Y9Uj4bpY5cZnP316WtpSJMc
m3pVe93wJIVzoehdjpKF3egd1c9mPz++dd2y/SICNIl4lQQaJYYkPUs2dFWpKTqtpKGYQGlK9nPb
+CXD0T2EViVaSjuJAzC7wkEuhtdaR0ON5RXDJxPvh22fdFuC9JEx+2rm6YuOb9dIFpn7YocCqLCJ
WYPnGqybugIMqAE9xEsgZvdXbez2kgde+40RMLBgaLuXI5DcBtUlDb43NCdxEguRRXlsv7LIF8CT
vxoBo3V5Yq5uG1OShH9bUhcbDSLc2IGyNXjB84H+XC4OnV1+By1hflGgPpdmn0psmnK8x811tgBY
Fj/X+fHPUby+gZfURk+JKI+yqdcnZt4nAI+dcQ9wNG95me/ZvEqhJ2fnb6g/r12gRtrwEkiH7kWs
zUfrJcPIEyV5+pYHWSzNrrpaQwMV55Aymob9BoKUXsOrG6Pid/1Y2CwMmXPYUU//1Fw+WNYJT2Jr
aHZptoM4No/I9Qnyt+9Nki8u8Bm2fb0dv9SBQgi3El6NmC8XyUkkoTGNb5bgKr6vfWhAo11N0jbE
DRsXzS4YKqKjH+akrzTApF12yhak0YZmV8wcT+G65uVPXsmPtYJDKTq10LJPBpUZTPjH0ujOC4Mb
piOccLimg7WwGMw1ZaGfli9r9lxbOJyOjLWgYPwx9wtqWcvSn4PsQoYriwUZJyZPbC8SVtGK6clW
WyjTfG5dYUPrVdcb7R0AJ2ln2WLRFp/NuvG9kRd9nbP9rGFKq+lBg9IWRBAlgLeRXdwNrniETgW8
8V3a/Va8NYBuI4/iTcO4j/qXiAaVTOqm4EN1RIkCab/eFnENwZo0/pzprj4w2qkTj4eQCrFsQSK6
vGSmjPPxHJpBdiZ7AuCYgj3eolpm+qOO7ncHm7PMoiqXNq7KbFpCkpjtHqiPMRE8gP2xZ2/8+0Yo
rUsbHQRJm+qQlIe4R+kUmrNnNUMPioD/VsksjQ0LqL9RqEhzmpgLsV+8PKs0L7iaMbSUPCba/M0J
ezalZDIyXc1GhJGyfi0D/dB4O6B5aKXcvEfzBE1vL0dAoF0u/4ibVxqERMT6J1dXwrH6OLof+hbL
yo2JA02Qe3F8ge8MI0imQnVW512uGjrMuA/KcdLCQxgHeNdjh7B6Prmj5Z/UXza0VWLGvBfX3n9K
7vIBRrR4Q+9Q/cGVdnq79SUMn9gXb5reyr50t90Av9231fVMldoG1z1GMaNlYBTMhnwc+HZqdawL
ypMpH/vLqA5NJQzaIX/MJAjlBr5yqwgYC9DuIorg4kOG6thQFwbjzTMJeJXKz2QZvnjJhc/6q/Eq
mWr/bx4TUSZTwmDv2xrYG0RWSLoCLOwz6H8J9RI2vGTyCRHWi5VSXyvfYq4GXtG4JDO8e8j52fcs
KJ8SQOfnz8u8cTOnq0j1Vfe0+T3c3hh0r1jMHybagCR5L7X1AzBStThSlAAPO/BnKCqlA5k0jUD+
iKDuvz45gz0wtYn/5KgI2YV6TlpnZyrI6TIfjFGw+jEgewuejrHTbn0/i846GXrsB/cc/ce2HjlX
l3fEabq8J+wb8p+ndcNGesDGaJNvvj+4lHXlGqWqJMAz7OyyWtCISYjwRPPKkKPJIKaGCkU6HTvk
SuuCgkIwRQeQH0x3LWBf+S75Nh/MpIFrp3caqeCblOlbdcMXPaSizdj8mN0XGldbSfvV1L0VUMcN
AVgQOrswyTvO2x4OUauc67WDCZ+2Mvu0F1MbbBGbWCvaHST6nZxioA2l7I0Vb5DN8wozOs8WurMB
D6y+mCatxXw45HtgMj+LWrIIb+9yt3vbeN4pTGFTuHFBvNMJid0dQlI19KBgu3x7W4j41lT+SkXW
T+LULObnlNa+PtvS3coIpdpI736YAD10+2JOYkVTECK31oV8PGmJzrIVIa1NAz/VcezQQ7GJyYN4
IBgSXpWcm0M0qXnxTOkvL379YVKJ+QdaiBAUcAgHf26vQsjFk7XZIQOHo20nWSO13AW/YIP4ztDH
CuULVZYHhEnonbXspgkUAvSVgLn1UuopO0OIBdiZgprPJgpM8coK2OzAVPMzC56LY3Hwpy89G8Zf
LTvvE6KG7yIFwfzd8aP3uFpINgn+R8oj8sP/1YfccryLEBKkxv50cRlmYVSIfwcUPEhlzNjN4CuF
1ccpn9SggkVLGtTejFueJ+90b45fIEXq9URqbQ6dEc3Ofivu++cQ+T9N/zuZGHgppp/SxUKuEpjT
lBYaRNXDxb4zLp0LlHwdAXFQL1IkP+1be+Y9qGsJAL+t5IRjRhZz2v34r4rSAmcs7ASQ9a4WrfIE
j5ix6dmXs7Mz7rP+aI+F88+hofKTRl+NWVRMEj21Sw+z1h9Ga6+2EPj5rF3nU1+O/O5tF8+gR+3a
nWU0WVIc405yWLOHooQtBuWIs2safnVM6jZ7a79g4L5ZZqmiKlcmccNKE44NCy06khD1+e2VD4TY
FVk1+5XuLKNqwmHfVZOPhF0f6A+Gs+E+B/SGME7CythRgyHEllCY/j49x4XxmiGguZIO/8/NVYZp
ZY929K/ZLieCXQJ3R8JQiuKbUY3ok5zJmTT7BbGuGxfUpd4Q0D7zMO9zT/adzUq5OOJA802vsq3A
EP8wF/dd/IdfsYlsCLca5bQxBrwI40lvRfgWnzQNXlIJkTYjNwtWcVm+lP6x6OYqo3Imz9CgR0SC
eVo2nCjPpdtWu8PsBurJ+axU54o8VVQcH1aiHuPfbpuJzE7zAlKf8OKyw9MDI5mKNb/kE54agcLO
NcU3acyALatuBsACArEoyh6kdzhrzzTYwMgptoyeHbEAnlnvwlNfcWWH7I7/eEWI7c+R5lZ5t0nt
kt8p6lQujxBbgVIDUg6p14/kzfGAYcOeeu6jUDLokuDU8/iwUv/Qf+4ehjWuyehdNKxFE9YXAJue
Zlq8i6p0s1Icvi0EvLIEEe26I5xEPOW+N7nV5z601n5lpUxrXWRUM5aSz4ksWQXnmcNUCJ91YMzj
2IEfhH9lnEwC7kZd20rr5XsnVBk640e57KFi8w4ttbA5PJtBR608AALm0AHnrOeFasibNFy+WQ4u
7vUu8yZiTHtIDTHeCWpmDVXc+DH2hZ0qzqJWA6DoIAOu++IzNR8w2ukhzTzyonwviwFVY5DygT9J
z+5VqRcRzNWR7Hxh0e2QoGLMD1k87dA9fIqQqt6jICetNzHEtsgjdNu6Xj72krhBhk64FthnYcAf
zLp5dILvHE4e+SoFmQkFV/2T4N/FBh+ypaezg8FVz8VzbFzH3oVqCQvYoyE0BtttRynIl7ZOt45e
JxKrugKeEUnqKT0C96ejDmUe3psdFJZqbvLhvSVAjLp+L82+KAvwKkclu04aQ8erBT/wN7Wth0o3
qyksl+tIBvolOYmq57KA8ArY5TdgGi0EljmaIxmmLAj2B9Mlae1b7Pt/zqOmU0fRySQ3Qq2GVVP3
m/u1L0GyYM1aPZdQegp5RCGiyDiPftDpZ+OQSLBHpqWfZ3UTReGHDxb4gdA2fWxR2DiMgBhLmyIZ
fjtwjh9MKTsv60J8xREWFSSJ3rAP3Z6l8jQxu9Fa8od58H4cEhP8xEjETJqteKNl7DZbtHwL1KlW
OdZeKlWCzOPyo17Eg8PqqK547FCMAf+yGdamF7HNaawHKxLsjIgF+bKPdCnrfb+qm06N78TovbmA
yqgeo+iUtERYR5zlCAEMT7WQpyVusuHYU86Fa/x6msmybfwjEUITzikI6ChPrSD32AJqCUeNwrhv
2gADbIj6hSC6jTtJYNzeYy/TnOoae1SPAZ3OcvNN/m4Un8MHAuq/EJWvjPzM3FRt43KU4eJITP0T
mn76MMlavLO7m0Q0yPShOdDUZI4b/TxgJwcksUGZrqwctlOz0Hk4NYeszeJTJextxBBo5u+RVvuT
hyVW9+rXbvPp6oHk30kpFSxMPMvK+IfJLVFFGYvbXPuajvRyrmkcxk2cGhib61F9bL6GJnulqfCY
4bAWqoeOZilgb3iic51qnxxgJzdsDameqmpyapbb3Qbwg3MehWTylVo5KvLUuqsadE1q9gZNGY9x
SdQqAo8OZW7bqTexny+bK7LYndHaAL5ymxbe7hXwAIAUDq8ar9OiL6ygxJWYKWNzeaXh+HKP5Q/H
b5OxY35/RvwjdGpmw9tGC6ai2M5faxKOAWt4Vkgu0GIGO9nyIKavLYei5O+dVka17wcuiTKTA99z
2gxsuR+QS02INucE2UQnz3PXUDTDBGRIPTc5/qB7N3DfxyabhHR47YO9+3PDxD8f6OShUKanHZOJ
pglJ6Kja6BofEPu4Byg4RXlPMClNhAXr1/27vZNrZqV9GcT0E34RjbGdZPKyGfGZJbbdDW78lMcq
BStS6u7NjNGEdgizo/dpLyUVDXztvIw63JF4iAC1tpo6XCXrrAijQk/79WJYIUNLut/a0eT8bLoI
XLm/l0tNtkn1SJ+sc8npJy7Z+b3caQU/iUcBquCVxnD66jhmv+mfJIh9h8l8/oaCOOLw4iIiYjNl
a3UbYht4ISZM+r4JH0+Cna3lTJi+87CeSlKaLVjix8Yn0AZLnftrY2dKckNqXk1KRsXRiOgsQEEX
OGg29MB3oVLfA8rCtcpwiKKjr7b476D9gK+JZeRIorf4rxXdqLk7LidEwsxvrZ+A0AU7hqBn1mES
iOnneV74n/eypkrQBneTKmb4xHfYIZZYEnRUFDKpo6HPBxQBWqyZ5l4B08xP/u68OYXWkZ5CfCox
50Gn1qn8gkfiGMhcqpI79QvTh52aOa8bNubuUpMqHMLTkQc+UgYNnLnFWHLpJ8RRu1H7OvY885IJ
6QayjOjf7LvyRlUtSKBJMmGBXtVct1BtmGC141fhZ9AqwgT/eVlngb0gaHfV1CEggrYs8q1QYZHw
0PW3+7hkYh8jyjnFMrCpvJV6vNnexoGSmIEz0AgrNjw+hSHkQU8NiVoT/e9ZlyZqYdl6bI94jQ+S
dP/7Mo2z83zNYfzKpL66c5GjUbS4in1GlrxUpF2vn4R6h67Gi7SU6EDExuIKYIIhQ2/38RlXIvUq
NbJcFzigm5ad2Ee7oJHMU/vdZgDTffOSmDMJektEFebS7YbSuEueRqp2SmJz4zJclrzUT/rRTyUz
KrxByPmsPM036vEhrwLZHJ3lqo9lqTa+e4RHEZLYUPk7kFbT7iU4ruZdsB7lIVizDb83NP/7At9t
V5zoc8CF1W9qqm+SOUetuWndNyNRgT9Iljk+qySWQ/1YEDhRQJed+GHQP0igdJMG05PQZBWJxdYs
tqoBu8HWFNBv2DxtaqAjRRSY3F5WQban82RxfCLxb1W/uk+DlJoTT3VoSvFGQA4B/Mu3BXiYYtSk
DcE4JI+cXp3K9E9HSKxjGMBzofJXf/3Z1vEr3kM8Hg4Ceq1W9MYD4EmwwjGToqYEUSlbC/SFlV8M
Hd7X1FSzH+8InYh4kxLiPFAwGnCLCy7IjeRnVMy42ftMgVTy26utbWdaBxcrAxMs6tml05ZA2c+M
9oaCbyzFD9KDLHdw3FUFnfSYGgivalLeAs/1qcTrwOA5nwgsb+vRTC1mVxoppek3pmFfUpE0VihI
9am9RtUyP7P4sfJcWwniuzZY8UurhC2N4kBfZxU4HgSF7txchcwwxcM3IVJxscDI8f59rYr+ddcK
zVCn9conoiX8/00nJyldWsJ7R1u8+1IDCzAtYzYYQDfmWRrB3aWlkVWATLvXPshJTrmqLZ6mdTwx
d3cOVeL+femqEma0RxwFZ47EZO8J1x679+4/49PGFUjnUQxZ3iXdj94xQTthXNTM260Mit/rGtl+
C0oIsFU/iHighDTvu7QdopMGct5SHruC85YArMUGwsk//e/M5qBSV9FhkDVDrhcSG/z4mT+bUEFT
XMJX9d2RDzJQ16xEtkcFtQk5ZWFIzqVJNvO7Y8I9LNwok/4ZFuN4UD40n3Xn6fvQRGKz9PVpF+J3
QXptLMmnyYlB8KptwDQffHu3Z+7lOaTyW6dFZbNKAR+rGC/Z6D+wQfBhScCrAayRtFZX3QCv6ne9
50hEzTuCrFfDHCY83FI7WnWx/ZYha8Dl6pQJomhCeo/R+G9jrmK1z7HJQmBCQCDym6A9Mdv2pFrh
sCe12YgFV1s4xk//TZD855rZIMp840fHAFKTsHq/A4GnoMuhf82dzwVn3aDnLhF12jmKsbAdzA7B
zSAOIFHenJEKZ/TbmwMpkXoMy1XV3m0Ewwzm5O5MnCRHDAKvCYI+KzjO/z10W6Ba/6c1RlrULYbR
5lIzPcoNWDP6Ga+6DbCQ7XXlON0dzfcrejTGkLs2p8WWSODc/61oYbquRtI0eZfy92PXY2sawE7V
UXNYpBuDKWVc94YSRnncFDCdp/mllyzkntRIM6igB/qlsoJaX3JBwzCo0pVLtMNJgu98ev8ei5wb
Y73qQeYuxr6g53ZbNXusNBy8i+zCP/n3id2EC2WAAlMx6jDF2cbAADfhfELUxOwK0Kmhdzllccbw
LyD6bN3kkRa5/5BrHoSSQvnBZlHEHC5kEfk/pBzrgdtbhqSDLPOra3Qz5JLAZNBSxRhk0+i37k5x
g7jctMY1j4rr8cMCD7tNithKl9yY4yJZAagrfV22u4fmkt/qJUfpB1lf3Hxu3SuGhlLNH5nuffl7
q5thT2FSLRpLM7UDyflk+vN8WoqA3qhEvn2MnXQqwIXJlV9ffejBEckfECKKKB7bYx78FU9moANQ
4NDnbT8CkLSv69mbQNQUba77eLur+uBCRHgW1J+ue9S/IpB0rIXukzG3QMqrDC0P19RTN1yxq/Iv
90ZlJU8CTeOHrIMhJ51AIBUUBx9nO15Zo0PhQYBezySl9tN+7APPj7rGOZPsMZo1UoNW8EB0i9Gq
XxWXoycvh3GvF5wtDe8xcBVixT9ohnQPa8eAQMuWqGbzy4XbzHD9mkwpbxNtFSiVUBLioiAX/EsF
Ef1QZkO8fGRRTDr085ZY/2DnNvw3LPcgTNDDlI0FyVUZMA/DWkZh0qtNawOFsTgeaiAc4538QQPf
V3DqK782Tl0Lrhk9PWFZiOAG4IYtnpwwG9M5ObKyvkfoN42MFZB6K+sJca2YCBoIJZwfRW19zeI+
HDpx594ZsLYqLMHUtQ3ot5SH5Zwi0Aq8NE0gvlvu3wfaJI5MR5fHP5om5WfLdDiuRG+mWNjvz8Hy
71NsOk+1yfpz5JK6N6fKfaYVkmuSklTJRwr0Wrokr350tktyGQa9a0E80Zr6+EvqlJS7qDfnTZE5
z53GQHd9C/bi1Z3ONmN0z7ae0TIQQia1m3L49zH06ubc5hO334D5bNH8KqiGs+QoHOdzLtC+xYLS
8b+xGV2+RNg2+LDpQZK+AYCTW5eV4eDKDPjEyFydViANTp9UCuCt/sjJ2ykHlsys0FIFu9qXZCc2
XomNTMnSW+inFefJc8e7/SIsknBvo1zzu34XwEiZsFsBg117611TWvuqSujk3l0qTPyfWhXuF626
75kpVgmTWuACZFYomKPu8BpA65zhKYdGacAEsEEF8Sunjhk5mq+RO9+WqdMtKDF/LTnVRoEyAD1o
p/gyJMPa12xLVyUVhmadGYlMR+e50V67zACZHZubAtCpRDNr306psv/LXyhrLOhncG/n5nAuipbW
O3TuiqkRugvtbVrIiMVkDWvLIhDK8Ij+ego7ab3dspOptCkNRRUOpZCW6fla1s8kQOIJeEvQNnWO
w3IFGgSMV/OFZtQHlejvsmjdks4NoOycMlIeYXKzrjVFe29ybBvv+UN38StlzxsJ06IJHduh2bug
dkndpXD8uGRSVFod8n3XYnl6PQi+qrY0IiDybBTtdNslpJQ0FllLus9Q2JxseSgPaQ0xmRzpr6OY
qjH8najDcayRuFmPSzSaqFeUg/fBQTfl6fza3CKUALWWyc3Enhz+QKa9xIreKQIlTzs04IIee2D1
1oLxtyQgfeYnMCFhfO5rztJdQez2XTrzdP9G3xLZobaoQ0rZvQ8ZGweDh4mHsPbMLLwvkf94irxZ
UIDp2Q4SqTYAAMEKTncR+3+QwnvGjaK7Hrr5XThWKedshCghdQCDL8RcV5VuXaRuNgSCR4D55Ncw
FqD5xDqT/tbKnElI8Y5sTRjA9rF4gSayrOR7AwqvA06dX6ciLMCHWKYiGSvPljQxiPduhIp9pY+P
kOCU8432sVWtZdLEfqm5k1+uhHgAOec+yc0VsSSBU1L4qBfJSEmNCTQJNe8KKugU8wign3TAf9kG
tVO84TxNYzqTOlPXFtPrZe2sNr1G3aKzAuiF6jRESC1e1DxCL0ZG5LHM7eHCOtNEOTPeHxJBplJ0
9noiyF1Qhc4uMirYwLm2KALyuNCRUue28pk/rN6r2L0QtX2NK5zooSrlSkHdiRleft56xhivqQBr
RBXpKoUgQg6wgJO99EhsmiXmN8tJrjM0Wo/rEHwqfLrwO0+6M8742X6pQ35QTcEwTcNTouCqlgIm
IgBa3AORKumcgmgpLg+Ne8oV9+Ht1mSPG6vs48zqYzZhGPfccp1Mtvr58Je+xkw/KVk+Me+EZfNO
lwCeZLA2q+eevCZWhE3udDAo1wTX3AoqwB3jtju80Y7XixZer1lwEq8g8ojlvmaRceJ9qtaT2A19
HustakUe/o9hYCHwuBlTHGrfdDCUj+m3uPayqZPfhLKyWGafkM9RtuIQl8Kb4dzcOXfBSWYt7bHR
NcKGvumNnjhmGZ+BE8HOEMxhpfVY8yMM+RrlcY7phIfNxko2ymRBzJTD5LHE7H25xFCqVE/9Gmz2
o5nHn4bYtPU0onhID4qS8BchPDJ4F+UCqDgmdssCieqinUf0GPTe1TxKk13/7jF+2Glxq1UjfIoa
HJ84FPecPBU2aQUo84ybiwmqWu2MAtaie8XEMXfgDoWFS4fD6Tf2Dq63AOA+cql40FMNuQKH543/
WiJKZW0tjU/q5flb26CCofibHvvXbh8NJBQS0rWp+LsCzDAGT5EYFwY0uyV1lIiyATIzWxy0MeDO
M/1juh0JIBEZP6QEdApEPEu4SZ2oKkOvbeAwWaUz25Z2QJMCWy0LLOeOul3vHp/R2zgsOk7lGcug
hFHGuQLGgzP1K3X+KaOcl/sc+4/SBE5GZ3TG+gay+79rbvppjAHDpnVLdFh+v1fBbHRiukQScZo+
wd/wR8eSF0Lb6rbmLWoFt4zsOJ9+is6JFLyjNjAjdEW6NcBtj7eI1sSq3ODGxhl87G9PWvRGDI3o
IBoWyS5M3aZHz3A17GJWPtZFYmxJpwNLzZgLgY/fQhVkyhJvAW0MolJzwCRIcUCwPhaM8G+RzPHV
lTgzk7Ru69rc4NdndRILQNrlpwD6cGAvQqfVm0QTUaFCriKwhCCWBltronriWqipMb0ARAGnP89Z
Tb57EBDbcZgCbQatNkCITH/5eSOIN6vKAucNAYx33+6uen5NwqmIZJoWwpdWYZcPrY9Ubi/iim2b
sA5R4Bm+V+dY5CS79iQz5diG9VN/8tIATFS6Etq/MIK/kwYvmomYyL3K3/1LbvdOSgJX6WuqmvmF
ggDgYL4OjrvzTzr7nyXX3OrlzEbRsIcJjbm1ZFHEtP5pUJ+2zRtTkSBsYO9cFwN9W82B8Gcjsrae
ont8hdVubncJaA4O51YSmB/Wqja09TQ/QH360FDkQ2qU0gAqUVLSJDFM7KCl1frOuJTUDPVhM7uL
EUT3mfv4hS+UB0YNOrLB33eHYk7cain/SZTfGzgZ+nmKi4xqsfLhtgBtsG4IVchwnbdDE6JhIeMW
j3dCFGQlnMNAF3p3YAtyArO2XxjXj+zXSRJ7YHG1uE338q4PvBnYXZoTkFAXpBOmSzHOGi24TIs8
je4ldPXv0GwxD3+QzYX4TFq5J+9c238on8eX5VBbAbAcmYSHRcPg+hJPLvReC1YF1Rfn6QZsvidn
4Ziu0h+pOEMehKahvMlNAN4HoBQOdgu1n/R6oMJZKOdi2TPIY8NHfq1SBCZFA+08PRD5n9YbkA2h
jWDqu8AP4W4YKlbSugzh3BXRplYrkO42oqGfZkiGkfN5zVKUcKur7yBRXqT2FjJapLgpf2+CoRF/
cyOMgl3vcijjaWqvc86ZLPEtdnlvLymm0vJGHjfszbaGZhJzcTLjFnK2/b+AiX8VTPlOK2PsIAqJ
bLII3jZS6d5bFgbXiJv4vXRBGS/Ps0ZtPQpTtLWg3ehWetsvYNnc6LPHMF7JMdoEI+WqdxNVAfbk
DvG65Mty3Na6IzjGdY2imvllYX8NxzTFuGZuvuCsEn87STnQ75cd8IyRBLxuIl9Bv9XzJBCGJMkP
XDtmD3d7amgPKr9loc/jnY2sZFucfDpjsa1W4GVcfgIBGE1CzsKYC+1mL/DhBgaim15RaA/7GOoU
PvUB835Z2b6Br5JXlOWRqfNLAK2ajiZB/86TKdGh4PiJUy7DglTN1B66AGO7sc0NHiPQfKfHJhLF
tBD+pjsj0cJyvCa2+hotlRp+5y5xR1nSyZiHfLghzqAMSqh7hCbBbH4BTQ0Iqc+wzkQca9nQVa8L
WuBkHjzmJxFf2LFIsX31ceiOBrCSaKEFjxc4UkxDFP2M6qdtQ90jPq+U9YzcTQFoRpxmwWIVPKh6
I4g1bT92nTKW/fCN+EQ0fSFnlyFhbmZLJVfW8gIJvsQtwzOb6OJp67AZSAC4jAaxCHuGHeTl/Js7
4mSHrGq6JXwLy4A2ObFzZDo7VxaBkU+6ZNwMpHtvE/9uxi8bUexwaEBEZZaLqaRCGa782x4EcPfq
E3HpgE0nI/GLVCwtvyw+So6P4UrToQG5RawIQq4mfyqTDXkbfrtplsVQCk93psqO0Y2GqQCQ0R2W
B5DP2gmu88VZTxyGZc9iQGZL1H9dd7sm7OkJ6KpQLycr/3u1P8kcPVQHhLpCezLhX5V4UtzYq6Eh
fBiQ5IfN8GZJ9Nd4R5pFG1KaFuPDAryZBR5KQzYSEcWIOpmSA69yKoySAYVddeRXNrEFI9VQuR27
dxaIUmajQNoa37TkPmyZNq8EYNiFoF9XRSKFWoReN6WYAqqrjP27glH3IBAxMfeV4SkPVDzaf5fY
6LtrA9zK17PhMujHSltLxviNGbUeFyAKJq0F2eu1gwMOdEZ+QVpJLPUjA40en10sb1MVBPcNy9aP
hzJ3UdgVuO7g4KEBa6j5qIpcKCNDsmqEPYLJ+5vIXcWSj7Xvbrwrldv1iUs2N1NQmqjuLdBNeAWS
NMIyE7I0hEj+QXvG8/GimLHWiuBHYaV1N1EM0t/+x3QLMmB3b97vgVigeP1QU87WekzFssvuc/Ph
8TQmrL5UOFFPTHzms4naHGmmEYFu3GIuI6Em4pPSgsP/Ynb9MUnAOP/1bmhcwtrmQDzp5UpBTs4i
j6DLdSkPLXYJipFKqBtu2YA3LrewSq0BLnA/8wtvA8qqoXN35K5cybk4QVbexGqDFnqWlmmN5k3b
2wZR5FGjHlQUAVqXRZwIdEP90d1q/5Krl6BKdCaQEo/aNCUvdN3/Fitu+EYB/eNBPA5wF5d4Q1AO
rKBz/FzY6Aj7Na1fVvITBKaJAPV3MNWJuLhztdpCKVvIMOROl3pOQChWpNJxUTC6M9Qkv3Sfl2NJ
qdKkkgXPKE9jDaqRkHMBRB1LoVb8wKRdypCjMD3MtGxVj9/rtrImDBkeTtPWnPImZ/bDBZ2lcu8C
me/3xBzHsba14Zvy7mzhrLB0CmofVzdKtte/0mdfhaxdHCk4BQRPp9Sn8ipEgNfAmozN0S18rCXT
W7sS5fsqom1zSGsOVVIJHKZJg+XdfUjgd4+IM2LEuKQHwOLoTVOfnbAegfs7xSlmSvRhtb8TZl85
5b2QDMuy9/uJkSx6t/+SNWBcCaVGbL2PJuYuJmqpByCgiGpgk33tnC5H5T7uElI0mK1czVlzMZXF
QPSWO4oeh7Pjhv/0qXhloRdeYrILlBlqqeJPnSy77JGV3jRTTso6+PTt8INgT2CwjHyCMGWd6Dgi
ZuLsarMp0h2HJkaux5bJgefyUFBOJ3iqU4x2rB72D9z6PFg6fRGnIiknda8KdSUxzaIYaKO9X6X/
yjh2ytwDIVafx0P6/ZTAmoM8WmIiS4PP4/unwrsHjYeY5f68T0Y3y8k40t3x3XZdWJR06brjcXth
+wWE1dBeQhe1AQvPGUJuGTNcMYHoj0EItSJE/a2Qakg0ttA/NEOtfp9gJG+eqT/k8AHVJesgkrCo
i95Tgf2aFQjU2NXURe6841wt4SJoTvWpoPpSbFNFcIkylaFUP8CNnuimeOhcg9EkDaGMahK0gvAm
RI3ueP2GahouV5x+2bA44pNmWowwVHJAAZnCYmhUCwAa43sffG6u1XV+gVKbT5Jqz2CKRHHXe9Qj
5dTdZToi1jGORY3RYBrZ+zXrxAA65La8ibQEAK5vLQ0pLbah1vAwW5Zn6/QHJwLqTXMcrITABQU9
eiYygmDbeImT1r0FRDOd6SEVegLCP4UL0a5TaKDOe41Q+R5FSBF1CibwUcQ2am/izy3/o6U8TAIZ
45ZIEyZBo94+R1XMynqEUu/3zDLxRXddBj7yZsg6h7EOqeRU8FS+04pmH/dGEZpz01dVNcF8QHwG
HCCFU48QOHNvXTdqTfXHDhNF1kTsP5u1nj0FxbkZm3RZd6EgWLPn00BgCTNde1lwsZkmLa3UjyRb
XeN9ZbtXaO4x+zsnDxzHuym+DHvO3mH/BdRC4IX/kSEaKyMaVjKJ2bt/j1/OUrpewLs2vgi2tgqF
OhIZpF75yaEIhs1GY4T+yCtO5Q4HhqK6Cz2NKdvVb++pXLGQXrfyQdn8wlL3IBCaVbXSHrVv6ulO
7qcbQr6fR6oRBvbU7kw3X5Q3Q6Po2x7IXaCmcH5t+g9ZHAIbvX9DjcuwFWlEsK2tX8WbIXFa6Aal
8Z5oHs4IioVixm/1JndeHvS1LAxrk07B+yGDUWPELXh6QN2nJcDx/QfQvPGV/gmUsP9rvPSYDPv6
AtISx7WVukmpXQIUWDZTSqWGRe7jKXes1C3+6rvf29nbjtq1VwSJOtjz6d2ZjV2Ap2//1yyYv/YL
RbLCv/hzarIIkcU6A5SGqCS9l97l9PZwEzPqbTdaKUTu51tHx7OfZ9cK2uo9RV3xPYOCkAz92WFH
pWd4BEjGkIO6XRohO/HFdEiRweNOA015IPlhEcEMz6SxN30ca9dabUk7vB/LJrXQtqD+RlAe4sE/
JgeFKz4feTSeG02P3nFiar4SlT1cO3qETo7fM+aJ3bOewJtecRSp1C8lwEQFrqT/hIYSSvAKvBHr
sSKeJNcUt5b0etUiqoXqpoi2h6O6PTKGBfFyJ657mALwfYTGxIeZ0MhfuKuk0edpTlTNq9sIFDlF
87o3M6vIFEIFvKZ93MiUpJm9fBlggeUu1OPFP/rTFNeOdfUkzdtxNq+Zce9j/AtQlWwvDBtNHqM7
si4cptYlFNi+oJsX+cP0Q057A7PYT0jdxm0orOQsDwE5UZZbg74ILRRQIUAilAbvsAFcBNbMp2+k
CFK3XjgYYNWNlzgrtx9pHHQB3xTjPifd0Z9/CAJRBThDvsgAbZ+GO1EBMuIPAsyO54llccoi4biH
g5Q0mbFw7wj7xZqTQ9wkqeNao6f5pOyAD3nsVajLc0PgAhzKy2DRm41zRVGHvFrdKipFh1bDQvdU
zOdpPp4h1eHAFWmLCyNbQBCQ3tNtAXLld3Aab5bSqAO/l7LtEPTkMs3t5YAYZupPldVaOjt5QM3s
jbwekuMogC5q/U/KGTMOt7Gp3p3V2Dr33bEgGNOxPVm+fxPKR5HVWTgax90zh2W9bGl6YcrVirIs
Luwucp/gf8jlCXesWNo5Z/JZLN1mwP+IvLzbGeF1bitxE9pbdRFakRhK/6vobdj4BmiZ53ZUwAXg
AtbKKS/oawGhhgKQUzscXGRkbYyBLn2pkVP54evU5YXhEZ6trTdlwe58Vsts9wPchGG1f+vOlnIc
XYOwFTHf1NaesR6NY4kwRMEegqcHfITYudwKdKzlouxGxkjyAUZf6R4KzshIZ9UUh9ElozXic3MM
O1ECcofS+X63YYWPFl6n1Vw/sTPMzKRWCQlalE0kTBODJvnwPzoDtnS6/vpmBHTzgGqKWXxseMzE
DDGfU9UKxow5Im+nbUhvgO1E7xjNp+VNBf0RbYC4Gmd1UHeJCF0cNRRmeyGvXXFi7zHRVQqVgO8D
iW4fxU4wWWCxHSmw4uOK7PhcdeejfgtI79/yNeWBuobLd7oPuNktOS5NC9hD8ErMYpodrszTQ1H2
fEOJKr7kqL/vEQIQYKemQmq9IyCY3Tr2xmUvnwg4lW8kjnknKmJBjuVoagUqeW6pYk8fVQCoQCh2
NhvnvQumM5DBGdPCJBOb1CB90V9HMB6/mefUloHMDD3HVLi6uR9focYNJD+LlYQ9UCwfSbk7vmMh
sRqlu1Co6z0K/qBrIwfmctcYrY666of1/3pAvEMwq53cX4nhvJh4EqpGjLzcxI8OC92UUYQ5Yh3W
cBCkfNTOVF6nzKoZk+wDUCBCuiVC4VJcZINWJuJ6wwrgy9+YNOImbSZjFtrj+JDy5YNQ8i+Y8BbP
VmHpwxczdojCbz7BPJoZQjevLP2epK2Vt3H3JRHf1XwjxvppMZL/Fo7EUChAzwGnJsKAp4Yclwr8
HTvzuFh9Jw2cRccM9tQ2d8qgBhKBWCmnuBCRB766zw2MM0j1zMYhJW+JW0u2LA6IQTc5qzjE22Nt
7IDPRp13ClRVHdSd0HfOVANENlXIcw97nmWa3RD/qE9QOwBnzdrQpSAcSVM/guOLGcBUNiLXUPXn
HX+evLRRhQ/dDvqh2lNvJ1s5dvTq4CgeIvjSlNlbJrgypUJH/St0vLlw2juGkPtTSMu/wkrMQpTU
wBR/LFll/wGxOSvWjP7danSP0CJUF/ztud+ayW2cUeufFtlvPdrNt1vnCt3HsGP35wwVgOzKdaFn
xc4gD8O2us7tBFUsXvKZfgYTIZFyHdqqQsJTcMpilLAcifvaNcvZw2K5Gc3lKcdfXPwBJtsJSUQv
oK+t9HTm8tcTHU9prjY0Cmm9Mc7uj3AIeSpICBhFOdezGm+sI2EtB291jVFk1TzPTxUFjSqJsgVT
XXX2nWOUoulRW/K2OcEWTdwKljYh5NtoxyY8kfqW+2ZUJk0XKvViLbnS1mxfaMjr3CqaLdrrEwz4
nt57HPZYAX7Oieb8kuJeSvitOpmW+5qXhcSiXATQbpT8yqjflQI9FqIXlYaUhBF5/6tBxexZ3lKZ
GFdU214/fMdXWa7ICuurLJjiyP8D2sYHjxRO2xXTF+WVVGBYy7F6i1a6OzX5fiWyPgeYugbLNyhB
MCraYOPC881LHob6meX+qSFn24SG9srOToDBWtgJuwH06PQ6znTFdJvg5IQg+FMF55mUcwMwbaos
i0ehAyX8H5QmIDIuzYSYTQ3s0Ivw1+0P5UjQOVuAQZhDov4gdQmsMIBngDmmE8DaoSmHwmwPWJZ3
tnoO282BTUUZsvJcTFE9VIPChHhpbFazev+r+WeqtKhwrhfdonltEkLeFigGTAWZ6lfqcCvDWCL+
hAV6L+USI/Ah+570LG0BUCXzb4VgqIva70TRRu1UAsdE3HjnHSL5B1HRg6jvzbhI+dk5hCk4qEOn
xbKhZgib233KDS8wtGQJssk31M23fDEfVTnGPEeN/k4HQZiewa2o40JGgPA/50W0VY87erOGnLZq
3rBMBKSwbozSZy3Y7jECgpYwDcxLRokGrj/+jfa0B/yLeNdT/wIbmg06zLvveYsmTBQJcFgaFt2w
7wwP2nYZKHzFD7w2cUkVZdg7+slj5tUL0qSIW3O+lgs+yOgzDvpRhNJ13Lg6fEgAoU+5jfZuqjXV
6hWnYm2ZLV5t1jq9ozPZxWB5IzjGVkNSAz0ei/XaaKUMe9oXX5GXbIp43nRT9rWOPjsyfZ1m7t+F
lMll2nAWWg50KERxiCzsD6ynK0N9ZKcb8wPe+ohl+UskowIEVLlpLJLLSUlTAZzq0abVCrm8RaN1
tOE1UweAsbmEqVO9VE8FMMhRtbM0bH5mxPfBARIo8eqkT2b2ecxwIQ39CwIG+wX+arzdxkuIT2z7
Gv8D5M5vgpfgrXPtudc66YYRTb3qkQD/Z+OjDHwpOZ6e3BjcukbC0Uyhsq6GQR8XxapOF1Ng/7X1
E2Spsbw4tB31BaNhnwNiwh2dD2v3JPdJlpyO1LuReoH7t2Ksp3iHuTShKBVgxk9TveC1HYJSp1ms
oVFvccUrq+zlFZFQZ2jis24c8hbUcPOqa3VqthkVA+i8I+pr0dezlRuMKSDjKa63vZGUcLQOYIQ7
2cEFrjaszoyHmf2uHIejhMGmdYL9w7xBTU3qglr7le6eB8rDjyz/0pvmlQuQLSAB+y+Pu7m/pagO
SqL2Ghb8oJr/GmVdOcpmSW8XbAyWfOIuNjF8LrVi7V7in6LINunuNUhj5ybJg9Jtupp4/XIS2xmv
TTPqYTczdbz/ejqsHjjzsr7H6iGfiS6a9EAJgtNdJ87gjW2D7gJaynykNSk1N1IVkOQqD045gNwY
hCG0kk/zux1zJgRj+GxUO+1M1bKoDDKUoRSTaq13lMVDtNQHzWVJiP46wGUrqd48fEJa2E4JeA4H
ZQtJNzjzhWyQBkp/AO5iCmQSGH1Pfo81aRrp3Ztf33Voh09Vd4L9TPy/EcCVDh2hrFkJjJtd8uPN
Wyj1cy59MEoFTEwNzv9ehqRCArXWD/A1+pQeF43f7uUfJVM9M7IWXSRC3z1gxLU+HuEYFd7KLpvv
aGhwKMdYvnKIbxtwsIx+rdnxXnskTZoKV6ZklgGV/py+I5oWWl5qj+OUi9F5p0ats+lWU7pzQOpC
ubhXOsQSqYiWVhY6Xo1O4EepiQqRMDfAgmOSUMftIj5sK2nzZ8Qfy5lV0pMwkZN4R26ZsbPSBT9n
+OiiHG5Y4Qf6YBqN9/2KgGSiuRwJ9yw5ealboEL7KpMmvXl7oFKbCtfX7a42XZTOv762G36R6qTV
KQQC94wnyYDUCnmX02sJcHBrzhRW17KFLT5R2if4KE/v+gb+Gq2d4RXYn4R/pEQhgquhtFBz2lJU
KIaqe/0eIXDQwI1IrhjTrYPleq5FdLOnXeqtTPT5owdAHxXHeSGIgX9dYvvzZp+fenEJYALIth6l
HBlBd/ZOzbWu641J8qPEZRCYBeCmH+eW8nK5aXPCONTHIEdW4cjAWMvt+BcPa93CTr6PLccgpVub
fDMBTB3jnVnkKl0aWjMKuyZF1AzU4u0JscM7jivAAMt6Exv2nrooB/7rku4+05s/Tbk2o454Z+Gj
DD4yot5lTc+38bKSjGMVvJ+RfNk6JstS+NZshQw09UkZ0AtzuvegB74LULuA44d1M2veVGkwKgE6
oFI8zcgDJHn2u7W1KDDA7UHUa5IbuYn5jBy/xrxNO5egi2uMcU5cEaTjWcaeajNwuK22kt1gR9IP
2kJ2rQAFJkI/ZlrApOYGUBnGS3jadNKZE7JkLtfGEfXrCPGt1pB+MhYxmLAXy/3HMh4/n5TE/y0l
Y3xfZ9ZpPPWQs//No9Uin/m082hHvWWScCa5fpHkn1djyz+hA1gF0LvGqtU4KzaI0OHhpBpSYNqE
mX5tZlPqUbDDVH1H9ooVOwBg/6kBkFD+j6MJN3RRU03AKdrm+AU9fFtbFbX/ByX11JGhFi5IuPEV
sp5Z0yJNa8nvS86r4hQHLMfopqz2/Sj1zw302FTyYNXH53cXIUSDHdy5f+ixM4t9ycbkj+ca6l5c
b/wZTIt50IwN7EhAisWXpvDgoyr5lCHw9WpFbnBX4ykOB99vFOhaoO8xa43EyEKrPvhs8uVkvRUS
vIMJYEYr5W4cr0VHbN/ncKJLcF/ruHeVo77mXJzpMNSUNvxOnvOF+m8oWmP6ZBQ1Gw9KI9GVFv54
BZJuCdHiLPJo6nJvZH+RodjuFFMPMOwx1HiYvXrFG9oVNa08/3ZHZp5yw51+/KzEFzW24VNLrZuE
WGf6yHUEAFaVBi2Dy5ru9MrVnowtlbKgGxVqC4o5PDRbfztHqfUobadDe7biC2I9z2U/R08pZILd
k2RPxu05QCTRkj6dZAdt9hvizquGqh9d3L+9zXbzBVjZKAgsWlXAiFnZB6vLmYxFRxWIijthard5
r7dRcyVXPAxJyuw03SXXzb8oLFAcfwDPevip7Lqw0FiAJGvN9xmtwGNOVvbTL4prmAFK68DJIgVB
t6yyJrXz3EBlDklE/zjHHOEXYMn2CKsAK4J6uuOHsKO+87nMe63TLOy2ngVSBqUvf/19ipHSG6Ga
DY5pW7kkVEeDyOStF5+fojMGFjpYen7dUC8Fx8HloVurGmYWL4BTBD/JS/nxypDLvpJHWxkZ3Wmq
4bkiSEoZGDvPUWlQwves/nk57ymSGJYVgI54FavI5jjlazlRDav+DOxQZUkLVMXZ8vDFx+K33Ibf
lA9oem4QOsL5+VBevVXterdk2pDPjFViwlYKaGrIOlsBJ+ETqNFua1+gX3V94YgWWGZK750Y3Tls
yPAR4psR+EzBNZ8ky2/0SBnN7W7P1kWqbf1vJ8CEzKgc0YCBEfRuI1ZdAwm73PW70+hRQdrpITq9
wA+ouu3lqbxuz8LNp2LeaR9AXvWRe+kwvZtHBHCcHTtzCPREhrPFbyBq//ZcqiVlQAfsnHsXWfMN
7/HtQ7nmnpQEe1DB8SJm9OrCmVfMYwWN7uPEjJmStJkAzKxWTmvtR3jCb3W4zc/rCpks7MRw2K/V
BlxRBRh5fZPtHJ99ndRmneOdZZhYIo0b7bEMwOmd4t/INu57A0kmfEMnK6sM05EkRiWl7GVdZcoz
QABLd22VnJ2cuCbszhhZ7fLEnjdXzWtykwqx1/y7nLm0o7Bx6xXTl1MnqZdFXObHPWcaVvdcESDG
Bk3eNKmuK/d3fuj8hw+TDxUIBmgzsTVTY4hIjyrnIjjnqqf+pDEUxXszLW3PkFFJS+0o0eBscNC1
2zEhPChdPsFWS6k8SlynZCA05oPfOW0+M2N5wPJF/bdl/lfogm66/58nSc+hWUuhRWrhTwznmgFn
WF2vO1eT9TcPzIOtw4InD2Mw44RzrqaaujQpv/CfLRmKdX5jqLL091OUIEgk6ClmTGSpRZhidfKZ
PcV0g/jItDxU9Rju1LDQHQqoXfa4hOHWEx2Gnj0sa6NsiylU2yNrAmx2GNvti93NQtHw1ne5oYEa
5KyDZYKRQ/at7hS6aF2yOMH41/zJA3JRIAZAhQifVfNTwor6/cLe7DCxQfeWEOk2TiwYdqJdCheT
Qyy9tqmvlkimgWXdCeWTBNsWmr6Z8tcR3CCqNLTcMsPeN+49F6mHy7XuwWXl+Frkuqo72Dtn02TI
mV0SGx1aD413eKppgCNO3LOEBHgXkSsb+x6WPifWIRHl2zb70iUMgOEOmsbRFp7GKdGEJ91mdw29
DTv8jbWCOvgQ74WTYMt4j+CqwdCbACQwJUCxcjyk3qD7zTP3nYyqB0VLIwFQu149OTumvu8evr5W
wyXmuRJG0gDi04bZvGRjXxLX6BxKH0pAzYU4U351FKc6Nls0QK2FW4Xr8vopzp9Oqn4Ia0uzPrdS
NjkGrBAN/APKJlvzv/J4UzzKIQz0PVAVL7h2MAjbSBkGyKmeB+n0L55IA199CHR2OU0CQ/BRN9L4
rE9gEPDUXKQ4J7fTsIB+diEnmWiMRxi3qvBkhDjvcJMC8MVkDDJwE5oO0RtkRjc8l/kBUGrJyc88
xDjs2G0cXIRVRW+K8bEvLOI47GBp6+qAFFpvgcdW6S2G9YjE1DRKzRpKp7IvW0NGMWLOQQrV9emt
niZNFXb+yWxSO4li1bWgQHm5nMr1nk1sEaPC0QxDPZ8iWwok6bYilGtTIji0mY7N0+wRkCWJE8zd
QDcf44j0VQWYfBug/XhMqw0=
`protect end_protected
