-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YqjMu8zyfMcKVNxn11aqz+BEJxXLJy4XhLA0XpjTXYMAeKpFiwDUUWdarW+eWXt29KUAKMh0hoY7
wBAsIrLpPRE1qzW982cCuqUrtiOKlFJQ5Jf7VLqE7S8Bc3feV/UAhtM/R/7LsIo/+llowD42a6al
LRqBxBLmjwxsWybL6glV+rnscTXAaMwMsAQ9eTQQxdZEiTBEKilJZRQUCGmdRLIDoaLGYzzKoyX5
QrO0PCy7SIlzUBfgDaqE9fHfbywmCxCl+pEs5CzwYeQnIjtsDcVW+IO2PtH14WHNGaJw2Sx8wVQD
xYvIZP22yPRo+lW3T24ToueirfwxiVaEQtXnUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
dO2TJpZs4lCiujwy5AScBfPPVuf2x2MpMY9Dfu772xyYSebZeIqcZ9Gi4jwsmofNMoDgJp2PPQLS
lrAuNiwYRSkFH0uuQ5BGSOyHva4QlE/tVMW6Rladiyn2mRtpS/Q8wLSauOHd+tX5lInb7Q1FAfrG
q1nSQw8t1jAkSpx/vCwljv//kQ+oX4C8xVNYPm6w861yC+fouXN1ALaQvVtkYC04wi3ivmrAhBAg
sPggfO+BPs+c3+qyIZapsaafIE5KjqF8CsbCWFlCEHS7WvuviXjx4QID/W71I5duzcKkcBtPvTlj
E9E4nPRVfd3vb9pRV177FjqE5MjVi4D/fpUgnkM0SEIF8oNm+lplFsdj1q+CoMOWDE76FAhNP/XD
YZ4GQwrKrXZD3Vb3J2krVK1l5b7WvH5pwlLUvycqdhEwBsmTpIATexiPj/kXNZHoAIbBUfAcQ/ts
WAF6naVu1Je4U9ZvC8rndwWFlxqiqJaDA9E+En4LBqvJncKT3hRuIOmfWbY1EMx+5e/ANKD3kRLF
AJF9OJg+FPPOTsP/kLeagY0fRAqSiTOFS+qBnDC15CLbCOyYzP7ae3tMT39toW81lN9VI/KirDGd
jTJoHr9oK7Xa7B8QZKBGuiBxIs7keFDf2T7FjsQ1Qb7PWygBMbhm1eyVQ4wEsUvLzFA1Fy+hCcoU
fS2ZePl7pNme8gVveEW1Q/1Zrpd5aFFZvYof1OyVXeKkbOieLbaoX2prRgDm2Fw9P2S79pbt13Rh
3MHhLUD16PSuLFg/VythA8Skg++F1XtwysK2vN5WhlwQ2VFkDEqLUr67QXGKB+SAo1ruh+oUN8xp
ZQfsOG81pTQeEuyhSb/j/Q6L137nHSHsBR9zMQot3umkaklcQ3X/NpAwk2W0y8zbRI3/NV0SL1h0
7NJBXb+K87KSAaRCev0reml7QwQGfpYcz86CBGaFST6c/cxhMOCUbWHZMDmO7huIUHFsS/FJCvGC
o6sYBCPS2377SAFAV+aRvohz5bie56xyCvvzMa/sFPQKJicwEUStgOq/w+q/r/WC5EP1lJQWo6GG
6d6Niz9qD6L4kIROoasaT6RfSQxKOBImsPzsuolmU/T1uaKruccV87Drmmgd1il0oZy/mcogT095
+Fl+YRmNWYVg/XJfMoIWJ2vebX5gzYE+sjVpR1ssOUTCx/clZsmCBkujTRkX/fAzqOsKRx2TOI5i
aAmXoiGLwy0YO+1QF/ZY4CGB/4GzXXurU29OqZr3DaBd4nv6bAxhc4B9qGPGkyUGsXOkLLCVWeGq
PA2QrJW7hcYJrtxNwzc3rhocc1xeech/U5WepMpBGfa7DxZpa5olJdJnkKJ9DvHV+z/5+mbCta+/
MM9mMV+mqKFYp6VKoYLKC7BWjm3ISlmI7eJw09yp6mfZTn7PNn/e9tpyrNrotqIEkU/jK+a18TbO
GPa4aEg8rj9OQ1F5WT3T1I6G1H14s0aDPQuNORH/DdmJ1XzEkgxlZCZ3RLNXcVtT+l+OJDC6mchb
lvEjx/asjB+dUD1P8B0K5ERsLZ8Drh29fZtBQvKm3EtFqV2fJptdch84Ff+0D0PST/7hMyefiuIl
axRp2xEl0zYwj88SECbphy6c3zTjo1jpNx3ciAyVFsOXTYzMXhWs7ka/V857gWIwsO4klM7BNbbl
AYh0vZes7OTXa+yrJduIURwjPu9Ewcl6THPCWSYySb02vfAQJZOassZ9dMY8n4vjs/z3elbAu0Ue
gN0sLtkzt5lLww7z0h6BYFYzZ4LGBHxTXOYcD4X2HlQnv2Lwui47AWjkpOAJgY70VPMou95lrFX7
SieJC3lMFqiiIdlFSI5ENl6HmiEBFdEAwVlVqqMtjmmcwJjqtfbGAFji8OXnrBCgysvCByNZgz1E
Q1tFwr4wmht+8k/krhCYYgPTt7QOxAIlVeiKOiZkGrL9782PNh7Yh1Umv9yYJHUspcfcIesCoQBp
dEZjqvZmb4CyllCGCuglT2hTDBp1ZAm4HELbfuWY1nr2tmxED9SQLSYAMxj0Zdk9qc6DbBgW3uYI
Ha7XE17nmBIp7gfIEoCZ/73MMPPDtnBtK4bZqMB9Jp0GEb7pzUgLkrXDxQHJFeWU3fQOvk5K/cX6
OAIMUUhkS5CkdR/C9O6nUvquewsV3Wi2NTvyMxmwIG/ULdszmrFWkB0M+CGwv6ktL+1rNgYTzArG
SLTWyQl4skJH/4ST7pT8s7Qs1NGhU5WPHh6ShAFPzaIJNzEbI0Uko1Jb2r7SQuV4m/YxfIbWorTm
eIM7abFD6dVJiIUTeFrchXh0lmZlfJu8xlDVIMdxbXcFai63rvkEpqObCNA3m7TxtC6z6/JTJ64j
SKdcl4FnmtFcgC9Xf3XVL8VolL7pR+FTeZGG2gel7dHFPj27tYxTdxnvOEmN1/ijUVB2k0Sbd6lS
NNarQlxmEL/4gHrR60R4LoRLsNGpqJUl3LQmicKeV8dMTFUOcVJhR96KGGac2xjWTBDBNZMx+prB
UHdCgNdhqvtVUJb4gwzYk3Bz2Yaawu0Qt30eWqT3GRqdnw779P2+SZwLKpXX4xG5TzGlBYja6QMe
sGtTAEWLdb46JEmHGPKul+hD1ZwSxdDaZ1ICbkgU6vgiKHV9ubPFeDKvypU03akn0cAeZdoqeLCi
yo5c+x+uRlr9ewTJ5zXcdmh7Mr9ZXxT+gTTuDehZNUk+KetXsytdO+vFr91etvyifwYTZqzWmZs4
45+YHBY8Vdq3TBi8DvHaUthHAudGtOWBjyUxNbVWRwk6OjK0qFgCrAyXzjRXj+v+a8nfOzvj3Du/
RkStJOQmuGTUQhrrPmV+r8g1/PRmBFTbVdi19ZAEaZYiJbDQV19GM5pvE6Vx1P+tFBLmAg37Bgvc
Iop8yH47czU9b9MInHDmDGHnrfND7klgrjAJS72Id8sjRTvgJpkbWzdrZfgQjvXbqgkgT+NJLykR
yaieAxiFy0DPHmD6SO8lPHYTOT4VFQl9RPEq7oMBJWSjBuMJKS13SbaGM4l3lHb2keEWqH5FGy4D
tDcAdGRqMN3jRb7ixjarukN7WFP8TIHJvuzKDnvBE0bkAB6hEFw1JmNN6jXoGWhDjrpACHiGgMOv
1+Lr5yPdbwqceVVJtAAFrznWRsnxC80GQCg4ZdfEisTu3etKn4X/+utrOYCj1LBfwnPzZ8Xl7aT4
RLmUZBGOLHwn8q9ip03Da9TeB4U5FF21BfOoMS66Cis7erCZ+1qXFZ747IqJyl5/TEA8qbmCItBo
lPLsyRtOVp7HdqHXqvKrtBHUHbRDVN/9sIXcREIyf23FhJJ0Ntoko7d/Bu4h9cnmR3MQNr/f5OZg
sCmOwJzptJOVh9EVnQEqk8fYH7RLiW2CyY71OjE3N9Wlu5xOdvw9v7ACTQUahudLpWPYIpNHeVWK
uBbcL7sYFXT2vq5RwwyGp4cFHXj5R6r7NzzmPqPmtpvn7VYBaV2nlcEcNlu7+aB+K5538h3G0Rru
l1ZLhgGKb27X53UJukQShaY2ziiFkFeBNOKWb0XMciETE3HX9GCfb5beEc0PLnXIPv+avCTz1rln
EEOPJGmY8Lgp60uEbjbD4q5ZfBXWGEIKDNpXW9PaROXOxuH0E66SAK+a9sYjYZI5Hw0SErI4mLz3
W+caAONwEpbnzVsBUTONMRy9f6nF3mI80opeeoKf/KlWF4evBmAi7DwXJoCw+Oi9EnZ2zyqhWoNS
zBjvsNJZ2hrHKXQSK3oc7fVOuFeYGlGEGAvIEaT1Jxt7g9hJWcLrG/6HtRUstiLGJHiFJlVmLNzF
sQ4rlsr3rqQhnxyTGXm5elnMBzMmTaGJpIQT/L8r0Jw1ml29yAKhQ8FSGNWhiZKlZRFrqHSYcpYR
F8VWYEmI70f1UIe8TWGzUPCVPPHN2sjpWlifJ2BkOPp5GF+MJFq7loxJBasXAmFVWVK9pveEs58T
RMRoWbOSc0JDTO/i3HCs66izQxfcVkD3DpmRY1bFMDIomF0jpJtQV/KJQOIttibl/gwK4Uqzzkn9
8RtmqZl0FpyQwZ/RHb+yLQPBCujetA8jdWxxs4koBmd/+0J6Bp+K+Fi8B/sUGM+4LI+4ZRL/isSb
0YKrY7JuIXCHEK7pA/8hRit5A2vbl3Dhu7oN44d3nzV+5YxX4QQ84n7BcefvG7sMoOiVqUKlBIHM
+3vxqkrrTkvBS3FzfVv8c1P4fbGYCgX494d1Qmsa4iEivTa5pAE0mjE5pNFkKYHiy1/sFnWRSL2l
My2r49p3iSVe6XgenzG3Q6jLMH37tsPwgApfPy/mDFr9YLyblKPD5G1SaOVm7ZEDA2eaGzYZH243
QuUhGpmoACVoye0kDNh5mBybP0UbOd5aHVZYQbqxBe7aHkWW1pnE+y4ZuS8/Z/8wNr/GvuO0ZSXg
9eCNRNHnTSPkQOmkkFLqjBvDUC8s7h251RovQssTRhBUGehs0rT+eNHVVXiDfIiBtyZIWD0FoF2l
/JUS188bnHT5PN5lidbTvlp0bhtVRY0boo60QLBbgTIn5+1+uiAeSrXJIanYtbJRVZf5M7+CsTVm
0C6PiQe7sVi9V8z7nFdzU4fiumLw/QVW0MgAgG6l7uagbiiQMa1AYScTkK4ZpB/3zfP3yjzejyW3
XzODrFfQw8TZizaWaaEagGaaxX6Y8yTt890EpMGszV4W/60/rFI1sJDP7phif2NUlJBKRAz9O/Z2
0CVvqhWE9f+cdrwo4mX/ZF07mMincL/W41EMY01xoGZhXOJwlM+A7qk2CA/HvjJBufm4tjz1A59V
1Bkway5TMpDwjLzG/bio5QJNnkKnxpKFm0uM/6kvpQa0hY9kXr886GWouynWxYyn6Q9kUfajDMkT
8vkZlv8WDVtg1pJSXIfaH1euA7erAbW9maOz+mMrTlJ8RQuqUunyLFPnWIwebBNjT6J5Cc9fbkD9
/DSuaDyYdPAIYpgNTUPaW58FPczdJh2R3JcC8DXTO4zqkYR91CgPyT4wLa8dH0AH8WjkYKS8JGpC
IyY+9djpFXDdItsXESOvRB2WRRn8i0juYeDxQo4ua0/qnQQikUPffo8FX+iwQ7ei/49QmcDFoyPZ
rcqOiL/DBLeMG+Hxd6IAZ8sYd3bYlvoZZSuUKDoENKemkcVTu0MbK32Gf+Od4sj9xIGjVjYw0HJo
zGb7SrC5DqNz1hd+MSMeDoJKzItIGfn+s1KjFT3w0KmwE06d9jd+Ml+pg6PVrfVWNN58oN7DhljQ
Nv1jNf5ehYFzQYpWI+YgwYal4U/stw3zemfShNlLkkRA8drrcT0bVZW2+ZatXdmWQ39GLFphU0Xv
7JKUTUzA5XwdTgz/EyWKinpf7rz3LS5Stl4FnsHgoLJjun8xuMJaY7y/DUBY0Nkt/SFCh58i6P6J
hac5vY1LExwifRtNBp2kT4TimiCKOpZst44oKqdVX7buXAmK/mImRdWRo/pTrc6BRnMWkRNHmaoe
f9nkL9v7HAbRUYOR6G/ybVDu7UZ8E2cNrRur4csapz0hEnbSmv0hZc60lWSjJXz3j+HgndO8CsTr
lmzHwQtMe4z9sRlmZolz6h/+LT5ZP4h/LgJmqfzqUgqxuvlyazuyohkDZbixjr9Upycyn8Ej2utL
iKa2SH+vIIYfU9IPQTs7OE1SYtmfAgNqlVZDO4908mJeH5g8ksXl+OAcxiAkMP14CuEIOrankt43
xld0G72o9uWGy5gA2jxI0Q4L8bDDpqKviRKtszb0aKnv/4lGJqXv3n41r2Sim+GHYYLfSh9Q8Idb
l3q9sj+gF0U0f0Ziblo4AcWDQIOeV+v88MlnG3cFzK0qc65nShAe+RFGCCNmYYaEM0yIMbH72/e7
Gq1p814cujuHdSYlMQfwLWYpdwiTA+pfTDNUwzglGR4lnOmpW1+k2ndASfQuiXhjuykbUuhlNo7J
wKVb8Hyd9HZ4iotlXVt3yatR+omun3NxzoUHtlNzvEWzXG5xgau315ovJtnm6DlHA9FFv3q3zK0s
XjN+0CzrozSwXIwmGeJPJQhgOJCzX8ylrs98sZw8p50A9jESEHziPmR0ZY3mKE7ZNBu1ZFelUIX9
Ww7hSOD/PYKqqBoEbp/ZuxWojmxIn+hUBLRAyTaRTxyVt3X6y+48wYJhgJLCKlZ5IG4wQyNDIEBN
s5MRsak/AM4T6LNHqMJwieqsdW5+HVFEPeu1K1E+qxYVZKTmUdGIaIEJXcHIbTWEuG3MUmCmUSJf
PKjdWLEXQAhznzooRbM0O7XvdUDI5yTeRnyuYEtIX9O7xQ7kWXohetZSmu7J/QBIinxxLwqlMGcf
1sIC371y4cAtyZgmNFa1KEdgvM+qornyPFJtQKPJWERu9puqNdy7jnAHlyyol81/gRE04ck3Cdg5
8h7dou7Eh6ZJcMzUXxLMZZi+eoERX7W1B+HmJPjYFz+S7f+PdswiHTQVfF/MX8FD2ureMUuU+oc0
yK1egbSLD2vsLz6xiCaqeR80cSBJND/rQ6w+415aeU31mmbiLoUJ12fGEmbIaDGGk14AP6lQIOBO
SYbDwi8kvcN83Kthas5+6UvTvf4OCp/ddSEo3svy4GMROj5XKX9hbaD+v0dy3ahVTYhcavTEPU0S
jDRw0mMrvxeBIflIYHLIrkyNIRoRe4NuvWJDccQvEwD40liRzMduKDTOzi/N6vTQVX4eAv6nukBe
d8BwR4PcUGW7G7jx4jQuJZ7kmZO/gc+UIH/cktJ82Dzz5a0mwnohHYHqhdfkMa0ujhihtWl04CtB
59B7Uv8z9oG9vJ4k/4YB4DCSaozTANaNMl8/StsAksSlgRZusrvutAq1QicUu4CLZsegp8QX9xyq
t71v3cYM4lgAdI2Y+gfTbjBkMMK1s4nNJDfzkgHyruWFaIpWm/x06mvpx76GaByoP7dIYyRwbdhU
Vlhqnvvtr4ohEZDn2hDICjgyYEn188Eb+hA+r75OpTW0SQ18hmr5wt0NigVJsXaNSB/AqP4zGXKX
jcNq1MneXLi46HwJwfqBnd1R+vZikIUERKoHAE8pnqG0t595KbHSTT1MK3xJM+aoE5aBq3WA//sw
7UpP08adkI37xcyhmXnGXxZ1fh6SXjtiQ6mhs23s9sSPJ0eM6lDX1Q1q4gPvOgTZvSLUG1UrSfGy
fpZ9GvY1EX5seJN3isjK2AvJbvK6gKbhp05p7jQfpXnprARsuKTNzSc66P6VJltQqDYRmZO7vyUB
FDwzpUH70oFiLUZ5UDiEoHgxLADmcObuIe1Xok4ASUAvCxO75HCMfRpCU/7uuDEcLVwzmseyCQCD
8LG+qcDb/r3ovxBKIDAxJoZjYt8vLcW8/1eCQ7IRt0R1eM9nvtF7XL0bP9El8WinfChILMSCgWoE
81QoP5hb3zNIY0n1asc7ZOnsh4NgDLoczl0WHhn+8tLx7Xnh4M5NfElqkSUEf9W1GOfhe3MPgFWl
6yi6tJ2lwjtYESxmQ1fx2AM9a2WRi0ukInJ45AERU2/bAZqIlEo1vhkHu7EZp0eTB2usn2n2AAy3
EwMxKCoen5Uyuy4pyQsM4tDhM9kVHKGP+YmZFe8uFeXOPQ7UaLx4V0t7Ppm+COsvgSrCPB8vcLVT
/LVn4K93WnXO4ju4txSfU5XxsyeIF1quIXigp2tpLuFl4Wsjk4ke3LPTwkzmf2oV2UuZGagW5Gsw
/6b21V0G4N6iIBcwVvQdwQwXYe2WzI5iq+yek7JIvW0F9Aie+0lmgcGTeetAqbxiMIrUi+GXGS4Z
niHUyS7vyfSsnWvgqlBdYwuZjrwahmEffjLats5+purRlHVL99EXhAyqhCaXGrkAzZQoifRTeDoC
3tTq4DNQJEmV1QqJZDBosd9Kq5R7S2OgJmyfeXCAeTIbba7+zLdX6GZy6ySXthqgVsa4CNR8kMah
HOITwI7LqFY76wi/jwlb9snHsDwrdJ4gNkn3crcyCL0iUohASpelyOuO1vOc+aWVDvxiD4vB2f6y
zVoprd0Bml7QDBOQVp298xc6XkIxcasWWNNuFTUhqlVWTGwa34/JxBW/Hz3VD+U5yqqnrj5v+I0A
NgMwomGu9GSPjhTDqMT1/NJucounTmEBZaQh74ZCNZqkTVZFVzAGDx11/c5sC4QfKu5aMA7C/3EX
+IWZG0zs1W+OY8MiolSMH7baoDJMVydbe/LIMVtIa/uIG6j9yV9eZEV9I1jvsqSBit3ymFex6I0F
E4Q8QIzZpEM6GezwV/6fKyQouakjkJRYdiTFfGlxpnkSP6XkYLcRMe6vxXmZqI9m9Ry4Su++vV3V
MjJNUqneFmO9enDCGxhs1UJxlGLdl6wSBgv7YjAf5lbEYh16qstfxUc9MosrNmFWGTbWlIPKDEeL
j3gwQ5aIENHetufHxS/1HUeQF4jPM6h+pc0NsJthyli+rCBMbK0KYzhxzzDHNOpj8d/r3dI+kNAV
ymPnwhk30uQ9Yebw7aZMNDSl42fY9JGc/Nl6d3OF2C1BUN1LuaVUGob+4rrUKgfk4np5HAM3vKqo
MuY+kPD3O7LWfr8VRaAm+/7l3SHJsXv9oN05UWi63qIBqY80MJWkS/wk69bVRXZrEQHJKLmPBJdj
0WIQ6w4hnjAeTBIA+Rcp3zIrP7tBidokGeZbsTgpSHWsUGeD/p46OqzHoT0smQyyiNcTefl5THBJ
yoGwfdw3S+ezLXrJSwjB2AbntWFQSqywtboFlkUm+4U0/4LyIk3tGMG3nw1Y37AUNawv+IniFWCs
z79w3GB+2jqOEYP5Wtg6q9c1qQqGdj5SHECVQ38pQUcQHNcsQ8qBOtVDA6kpPMc0E9HUKL1PfijW
U7iDlOCj3rFhYZbAEGZypQlMNIpuJdvDwVomurcOcd1rOeS4gQxfLbSlbwnaK4K/ysJWFnkbN/G1
85qFpQlBe4OU8jelJF65wab+OIXMaV9h/0NgKAk4bKh0unAy/aixHWq5A3aGIeSC8mprzLReVheh
5dxUP0zGz219Tyj9hppD7Nz4Y3FQIsLKlJRlWgOAawleF5ZLrHWwAl7AEZQPiayUwOGZijtL9JsA
VoarvvFhm/7qgHdUHloE6wrCEWgHnK6IKJYnGEFfEbCKCe2Gv4pUdFw7VgHgFUOPxrgiPCZiVvtt
JGax8S6YNPpIjOb2Dq8sMNPH0gNBZqx7Yr+DLaKgz9Xs0ca1vR/2SUxBTq9GRjWYPFU5IpP0sw5H
XkyVomuuKDc8jmu7GruqnLqEzifru0j8k3DwsAXnKh8SuHezlL3qSxX1FaVnA2awWjJL38znJlLq
p4f2EbzWkxQJxnJQnGuErE8p9+o5w7ciHyeL25/KKWQr2GzFn3jRTrF0HdVVFMiWE8D7J7TjG9ON
1cBKR3vZsy8K6PRyYYrkr1yZ6AR8hMKr4O5RxOMi/VKxVpXVUoBi7oucvjVHZYoZx8rtlzQbxHn7
S7HTsKVD63UvvOlfg5SeuokjoEwd2cUAtpO+NCYBnd/MrNIHOMrBFvyj+zBL/XmOauQ35D2gH1JC
tk9lJnVuaEWS3Gg3M2m6H6muz7F+aM4ed0mIXENTjjGUj8s0Iig/PXXQbldgfsBmZNaeq10mBj03
5Kpyb+dnLpJVhn5hsWw8BaI7mVlmSbyZh3UGHSopBqa9GBruxRqLZaK+gXi4qSHDwIDD+X5P4Meh
7Ano91SRBVJFPcyfP48fG8y+CV/bIzXotFpcQvRmvXLK2IQFgSzHrOfRUJ7R5RWYixE7UbGSBBum
Z5cbsaevirur0cEAHPEadGQN5DVpfZe0NeyLl8CABY++LLYCm4r1llYCuAiJynMGbP8j3C3FtrJ/
Zv0zuz27D2eCRzuJ1HJmUNzgWzXjqpcs1feof19HuylbxXrD2i8YAD9Af95iAwHKP5UV4pgATSJT
ENP8toT5GtXIVBuJlOzQXXgfy75p1EPvtMptnje8eKkvCcyq3Gsw2eJivoQFE5K/CHTC2QYVF4Er
WBRrXQ4j11y0L4S+R993oCYMA4RlkrZKAW7a73KIvQOyxyWfKsUUYExZPUVPNJTGQGjFbnwI9Tzp
L4avD62q4k/+ovRDmKXi2FEnT5RJUDujTmTy4WfnzQPnXd4/+aPCACibQyAuylvJA9qCGRn2A0SX
jUldpm1d/FUp8GnVAjs0+XL2+rqEg17mxxT6pOavKN6mbSrYkGwUpxPWlimAe+VTM2JGkk2HJu7w
/9DDWKedtup0IzuJKA/yWlxtRNrkN4tY/fSBpZ2leSgfWVhuNsKccb5DRE0HvjtGFjrKaISJ7jsb
9b2Lc1PgxepD6lTPfw6EP2iCrzgg7Z1GEofLTDTVszNp49Yd7HAQhX70Eu4f2NTg/Q9RSHxV9p4P
6Zj78hq+e8jTonLA3BccJ12bkWXzR2iTpXkgQNZRV83PI1Gm6x3Couyi+yF9KbyXXMv71Ng6RDbM
AK6UNe3dH9omh/kF2L3LGFs8cwAVgRqFOPzIVhRpxCzxtdUEmNUWFuKiRhtxuvWMLGzU9kcEf62q
j0Otbllp5tX3eMbBze8cGXLx+3hFIWjNqCl+STbVtp0qHk6TcVfx6qCcXnwlA9zWpwmXCymSD68z
8gJGvp1CDOK5jxBRFOuipqM49u5q+j4mYubbXPAqz/V/FTMa3xXfLNK55ovLNIWiFlD0uSJiMUJr
H8jP/Q7dI6z9qZyasf7t414R+p9Nn0RsApKNqMyfuIagyy7YpAcs8e6DTgjRGqHrNcme/e/QF8EP
XyvivrvthkyL3Owx634ubKpK6GozBYsP4S1pjyntnj7yjHniSGhjGeDHMfPdP03SGDRicZVFdtNl
/62Sea3jVkRZMLfN/AJewnz7MH0QOJeqt0houK8b7sB7LkxDYPOv8NiivjwQZJRNS1hT+iFa6wb0
pFyLVl1e+0cojXVzjzhBp4catQGo7P9Gb3y/nOWwcZkV6fOBMlKQAE91c0Fln7XCbXxAaZZ1y5WE
8boi/e4c63NjpxkjEHTZOGkvMzbyi8QygM509SV197lvBCECMbe7ZxC9CbmokVut+xy/Ko/5O+rV
QMHk4+XVNP3ewn9mw05dAD0Hr77tiQYxHVSyHtJHuIe4LGkwL4Rr4onfuZ593otoSC50nhxEVPrw
PfyYUPLKus5QRt52mejeEMxB8rtbLE8J1hsf87BKq2Gdxs5YYm4xaomIDAZ/zoSmGSsujSzoFLID
o8FbqP4OUgcAFNld+67yv4MgR4b6l8ZmFkGur68h5BG8M/uVFGM8JzZHB6H66g8onYeswao1sWMm
GnZd2gII7ixNyWB0QF/cCqjUGYC907QWd69fFGK1xhWx/HEVLaZh4Bo+UZnAB0qo5g86Nyy6nWlw
KNGRSdXQmoAgIloOdjE1rDT4z57crEuJAHEJEsLLypQJRmRhL8u4MBwDa72etdhTkwYa3mvHoXYZ
Y1JZPZChEw97bk+B0fZ83Heb8OjLAEM3PD0ScpdPLuI4HoQfbodsmEIcEuO299F5313262phVIEx
djf5GPuj2YD9LkvC0laCCB9L745GvzY9BBf5OHWoJTgj6DpbeCY8u3h9xoRT9CzGsL9HhV7nElIy
FuJfKoLjagrz/2poUerB2yWapltcramFLIfAtGa/aY5wa3pK1h9IufI6QY3gsJ7ZYWGU+jJUYZ/p
7RTeHosbVgzdnCVWEq9Y3COeRF/zcc3v60iDw6GVO5ChiA+ooXfRjGAzHsU2UBn0S0D7E42V9ECZ
QCsQnWVIDPpCApZkWm+ubJa8wKe5ByglkF6SYsfrHkuX0wLqBDK1Torx9xcax4zu2ZfMCLtzbYxF
LxrmfX02LZj49eXUTSNKizu93ZpXbO8lrAz+KmLRy2175p+9UgTy272sHzxuZ7545/W5Qk0Ry/4s
lDj/VclFgjHdXwVMPqI8YYZI5FodSzy2/219g323Ro1ReRaaYK+B/jaEA6GRhXADWw99ZLlS+62A
X9Zy7SroUrzv05O5WFIvb67wbIqunl2TQHi8RR4fiii/zgs+qpBoHGouRf3UChFX1hXee3TLCT2X
pMd0HjVyFasNI0FTgCsbOzDDKFHax6/+Pc3hzHWqjulIc45HPymAbsMq0ceCNEHikaTRfcM00IWe
6e7BZ6fZx+yBeRCDpmrK2xNekPwqQnpKzUZJ/RiZW79iY+7So6scY1I/SR9SVYVuAa+o+I9I8YtB
neAI3huXwHTiK7fwcga1UeL3CXOFq7p3NpW9Gqq3PaZEcjpT8MQdrmZamLLiF8jL5M6m/ZcRjIbk
BADFdDpV5z5otBGuj+5BKmXpvasJwZ5FY6v5G+aholoY7SlAkKpirNUWoQu3sSge1bsyXvuvSuJx
+VCVXqHyqwPXy32XByEpJ5tXGttVqX5uLOVys1SE57a3ZFbxJhHvwl9WdM0ZCqWWQflzuZtALjPu
qOB3He6uo7XpqD26i9uZzs+vU8rKdLtvaU76fuSspxVmVhzWxyfgEkzZRqPcoCgcMhdsCXZNVnWI
LzcuNwe+3IMVCtzKQY348JJ6wFuaO8LQVBNC46JwG3wkE6SrVXECy+bcYUpmQ9QpCd+O3Aygure9
yRYDK3s9mLNqklH8zyovfa9rcP55FQbI9UIxJaN1tfv++YX3eaJZZ1RglMDHD1ugxSVSJPrNYkyo
npzd3GyYCrExFYorhkSJBJO7JCofAp7RiL24XUITxQmM5dr6uj2d2xfMgOB6YluRls34h8Maskn0
4VgERNLBVwyZyTXAi2GqYx0pvaWIQpQ/qvXcAomH7taOlhgR6rHBbsgu0FqRSqWgogFTvuunmUEr
wfmHsi7T/2/ezfq/m/Xp7VVC5P7+NP2wHRY3KjUTMy9UO6wOCIlxIwGrss/xwKAOXtBnGyTGdTBn
G5nkEyx92UjxbWsyKXtdFMFu8uKkI0trxPFCycokc8EUVeFHq4XhfN2PK3a/N/hc7u06uSgSXxcf
LtBGNUaMRbSTYaKMm8QUN8ZbWFSUms2z5XH3skGuE/pNDkPA7abWtucJEpatiSiULJjPHJkOx7LB
vID9EITNk8Fnf3uTC6PC7jmJn/VH7iIfpZA/TtpvXJDe6JbToNkbAVK0rXWDeYiBKJ6LoqY4RPYw
z5DkwNsD4rND8DqwL13I9zsd+vjVa8DOC76pUOyhn9uHQTrqy3xf3rxm9fMvy0q67HOh+20oalzL
cU8dioq9YyD20wsxZt5z/sWqNvTy6mLS3ffHJt73J/7eJE64jOmfiNIAisJOOeIvSbRrKm3CqgWW
di/FcWwtJBtnDca74lNw3aQ5diLG8yqPUGVLlLWhRIgZz1bI6TRZIQpInnSxSWO/DHshKi/MkTgR
lvAKkCMCYM16PAbrGo1cbz5umof/6MtUwqFu//OUCKlHsEArU45ofGOZVgHQzBt7e+FG8djsDe9U
dhHPv4xx06baVRRKtvJDgx6Vcc8ije5Qp9l0UxGQY7JQNYgcjKe9T0AOi/TOYLIj9g1v5QXwvdvc
ZI8OEpFqUmibZL9A3IhkfLjUj86iL6b73uM9L0EB/EbNMQ6DZEVKSX8Ly7ENpJ4Ff4JlZ+twnuXV
lFMjEg/k283mxX4L7ofq+joLZbrV4jM6pAEaYM0raA4GVmqDnDQedXucf9x9ZpV965H9uuXP1LXP
1oX/7UdKU4rdKzGASFFnk1TQPsz3qOPqwS1Det7RrVRDcwhqR93bK3crZ7JSU+YrEBSsbl+/N+nO
rTf7sliUi1iQnTgGPK6iSlx1l89Pap4L9bycFuzQQlt8AK670xbqFYcAW4X63qKjgLRurKSheY/M
VAVJzBzHMelKiDvs8ecp13lSMAmt1KG6yeu3yj2CqUbt48shZyc7FG/g/0bzThahOsl2recI53ch
miM3Cdy78bnSjAAhMYxfMTZxZwvasG3svPbvRIuTOaDEZWIogowm/mCdPJtK4z5Jg7DA60A2kKhn
oWDT+WoZxTcFcoFSuZ4hkNSX0rVw92voQZgv8sDJ0yrBumaZuJQTSHr89+z0mwFsl+cW97CBUNve
yuTjnd4fjqRAU1Gb4PJDpfd/G2LNUqqjCniZZv3PUY5J408jOouo6jOuj9kUkUys8bxJ8X53HBk7
8px+ZFcj8yX+TNuXvGVBSfOerDOPJR/qhiw6rjXuNrd3jCublTW+t6yJLILIYNREEPECVmStdbpk
+tH6rIrxBtAEzwbzneG3T1krDwo/1TwEZj6KiAJk8aYCF+XhkJS74owX4bGASDEKuzHy75DT5IyU
n+qM91l3KftGdmQkNK17WEhfGnN8SiER+6b37EVD75uz7OkWoLcCJWOnoCUjbOT4QWIlhnRryFDG
i8HMcBarN4IqMeBZoQUv/xgiOjKUIhZpuGkDHSxA29FxHNdQ59xxd0WSPq3KfUznIv5azdQAAkeh
TF6Y746ftHA8QuSD8pQduLN36WV5dP00/qb1j0CicjGoX/ovGOCaYo0lCdmB5LTs5SwTcoiN6SyK
JUPpPaMYVay3C3rRw25cfIFZSAvl+mdNVvHGzV3E+IAww8QuWDm7qa8ZGQtXugcy8fsSmmxwXxV6
YOiN8Q9aUZiq5gF9b0JSu8r59CS6/lARMdBPPSjXYS0FNJhGKi8myjI/GvrxCE9bVXMHQor4QSKb
IwCky9Zbc7Rcvj2XGFy3hCbG77y8xL6cvVmL5J5FhvEE8z3Gwps3tAjZFS6HiaOeUpL2FVVttJxe
pZfzMN4bR9Bee9QIrwh+kOSg6Cp4j58rBAn+EEFKQkc3ChllUAwfx5/UeAvc+tvDDkMJSafFflvs
zGgGVCnXlzKcCIRFIEdzhTvJhyahHgwFxd6cwqgSJiPlpIbfxk0Q+vcF4PmCmGRz9oPn0alx14vA
4OPmmgtH3TN9wAp9s01h1BStNpKxa/384Gw9rxTeDSpN1HmNRwaTQW6X36HKJuU+/SCDxTwENC7m
I7375C9EV9AIg+POCK1CWLOj1OludJ+y/3ZZpZtDAx/GiL6VryBPxBawKnmGsPxOBOu6WdGtOwog
MixcJaeAQblo0wMlAstiyrKv0xBtxotqpTBV+jDoNum29cM+kBptkBHY0nmBHcgBYGD064+scIa0
HhlIvFcfDKvn8ZttC0n0/xuHfAaZFbjtTMqfhwCKQY+rSeV/OgVMqCq2fshSXXlAjbJGLQcsXJlF
ZXYNX8+bS5bKafAXlgnC/p3uuXyPNUCIx9m2XVCXCw3wjmoAKLLZ60gwzvElJjKpBsbDwhuxeqYn
Cpk5P/sAPkgLdWMsnWHMjSzUav6g/YKD720Wws5HpMLzIFGz5QPoVVPa1JmqtIHHONIUDW3m9IXj
+j04nLSE4/9KV288ime4n5YieKlmusbJjeMShnEMSCEBvBBFdf17UvbQuzRVh2vtSCer4Hp/ReAR
ikhNl/vVOl4gHplK+EF/EN8O5UHlhbzsULQDNIbYmd/DRqViVqENyh9opAM+zEkhFYgT//ShVCZs
dEsIl+rm0o5mM0lopTX5HRv6kwumtVX+clpov8D/XNkOsQUiLhkh/9TQb1AXzCeczNLEinYC7roD
VNMwucmySjYbNsiyjsPDUiHH4ZTMjXiZ2Jn04r10IzyNfMX9BDKWD4VEP6Prz82ShEHwROX1GBPn
HTY3LgFG6M/BseUuclmN7UNSvFwpv3c/TjTnkbpj2ksdRFIexeWA10fAOd88m2ryI11UbOYAw+CZ
tdcowP6FGYChweh0qcAsS2DNR4vksVph7k+Ru2Q5t5tOUnsdRHMkgfPMPTZwnZo+uCMTMnqduSWs
FHeM8FuzlTwmKAzIq64sCASQeh4bJb4fYgpXpK5LsWuTQ/qbcWRzIS97oTHwcu/Nz1warfARDzD6
uVRGQTN2wZpaN9i8Tk/TkRJexITE8+rPCXDs7fAKeHSRChpWOUugzEtApp6ZYeMu5DJ8Am9j2DTZ
QygbtJD0PeZDU7fHUPjBENoO1Qsso7xj5b9pT+z7gwtxgcAR9ePbgj5G4Sckt8TE3/qMBMrwyoZh
1PNTxK7Xy92EYb77CNhqrlHeWmAXpPPj3dxNen5mtz8RdhUTpXIytBv1hX5S3HMDDZwLwtpQWyBp
1LbvrnH742PImC3UZ2uftOw+eHZ6UQ5fyIp2oOswacZXXyf+FKKLi2R9CQH/sOJr7gFYSXk2Xo5c
91HtsE53pi+z3HOAlYNH3qYeDN1Q2Ky3UN8cWFAdFQBwisCxd92Xw138Xe8iKb5RwxLkmeNmLqbC
V+IZyWk4wC6tKdNREJ3cHgJ3rWanr/x+daw8niL3JkHes/A1CnceilcrxdWdOKeVZer4CC4YYxDJ
vIQReSEc0skyKo9nfrLsTWLYfo+NEXwwABUfYN4GF7+UG6YvC8VhRQ6FJONhWqu5uXRV5cfe8oj5
PNm/NexF3TYQX3euZwnbdMO4VAESWa2VIKX0wTFoT2807aoAK0SwNk9VMWyVnYdFlgP5TlJEC0rS
0icIeK10ugOQ+/qQfU42tAEqGCbzaeR92yeoe8zVFhWxak9bUEp7n0SiQu+okXqQUNlojldhRZfM
KtyzjMhDAIaFYBc89a7/Iw5uK0ZO6ikCu2ApofFJLqLxmhBkyJxNV6xsb01I+4yko8yZTEk3rR3n
RTC7NH2n+9UqY58qUIjARa5oRL3mBpkX7PcrN4j+vkA9jotlK+381Yey5Rc38Q8juxlJw0iK3qox
wbiW970/OVEK22ejHiabQ1MeAv1OpGtJP3BY3h5MaFnYJbnsLKouZ+JK9EQJrPKP1CmUefb2uJeE
3AZCUuX+OzphVLsb/nuDgsqgWUGXpnOYK9QTuGVEEDD4T9RzDvXICVY8+jFii/8y0CRYKTEUQJzv
/unos27G9sqB/P+T3YxGZUht72eOZf+5xF9dDheaet9lxhCX+iJ+pnex6u7b/HW8b1umHNncqpo7
g2NGcGBXlhPowjJoWNhPFXM/1sYVYxERpfOAmPsL9JuKlyIA2iIZ9yq1pu1JSc4GHot4LjoQECdj
r6k+3RmGAhyiAFAXtC4BxfMPpGszWdljpYOdEMcPvPF6AqDHi5feJrb3Lsjiay9en2jW5DPzgWQZ
KO2lPbwMMvMoiBwkUWhSSfz5jj4Vm8R2U/SZGGOJrFYH64tZwXj2zvT4u/A53JQIfWzeRFDY27m1
1iQrDT4XiwwUNrub1ns76Ruv1zmOmQK4TqSn4DdHndmWje6uoWHCjUzTn66PlJZzFG/0MConQWAT
6hRJvkxlD+HcOcvfp+jmLgMIdyBqPxPnb5Y5ZdncjBhlPT1Q+TFH3DTDEyqSU6rqn6ozObKuopjx
g+LybGE1UQygdlJCn6whBtuTiODbRVgm4gpZYFVMZs6kqO8chJ9DZPBjT3gRSkjAEpls9zwpVGI6
FwhdQaa3VgCh80+T8GuBiLIlgT9UAe+1VFXdR9Tik5zzkvrX1beyWN0yiGrcb6bOZ9DFHmBcsNpC
wdHMqwCocj285X85R2h670Ub5Om4WFQ9rsETLfYPP/5+ZiIaV1V3bQ93yj7pdsfWUSuLtpy11ZyS
erYxc1T3XPAeVzdaUkWcmH4obSmIxvglBPbNpeRP1aVQC7vFGpduemjyMH63FRfVrYIdqetzeNia
91rCxuMS8Ic1B1i4zJrGR+5Orm6b1okH7G3KAr1QHwoWKqWRd1L3MoDX5BzQYBVK9a+a6BwvVnwj
MtqbkHtLvwHmDOyL+NECmPd2so3qSNh/59M3CabM8NS+hlFPf+hHgfqTPBM+DuEPyFa4QCaLHSMx
pf7cXgNUUp/q1aY0YoCcrmFTeYZ4im2USr6p/wysmELvJ6TzzmV4P5oLe5iBE9Tpa+9SueBipRKx
W4EGc+SiI1aYIkYXl7Oi54iftfBQAFIQFnduzMYJ28nGIr6Hknj0moAUQVFx/UYH3k0igudeKbDC
ZmJplwqH2AGh9u1gOKof7yIHSv2mrO5r/lVdc2Upha6oYWGlkirsw4QUd2gxCkNLi6hjTsn4NGeS
uOZJJUHUkHRV9h1S0grY40ZtBaR4wMFJdXOf6m1HpYGRkFHv1+WmUhwzLmcnNmv2L3nWMs6eehKh
jk+U+0wHMX+KUx1LufVFKmXMohebOiRqRS1I786TQ13vdecjgTSwNmDjsSRt3Pdek7GYdf5K02xi
SM8PMyJKbevjabvXJL4e7OyV/qie5rg77ZbMJnBTJE3iGpQkzjAI/lmLqNQbXfGpVmG7Qp3VPOnR
L0TOjxcKHgl3A/ZMq2rnb2zSOiAWMANr22ovNOlBV9QNfIz22ltcF24ySaVRFG/KyAzR9YVnFq5D
/f64/juGKgBBXFufjDiestqLp/9K+HH+gor+GLsF3PryGXQuLxxV0DEc1F+H/cLpXFjdRCME7rs9
SlkM2nPq5CWirbQyfSUTdcUkN9xcI7EwHbeCxc06nf0GKTNGnZ7tgkNzcQyTpbEGB26IqziDoCCV
gzxumQUkaC2UpFl7zaEfjiGywS7N76duFsVs82Cw/0kblDtbzZiZwwgkBlrDuc46F1eRm3CzUa++
5PcAkhU3V+tqV9ZSIzWsZztc6PW29u1QAYdCYnnW2DBiouNEFzLgBgklAD4Ldck1b5Xtx1yo4F5h
zFpXMqjLkiAjswDen7b5FU7WitrQYvbqcVFE//ffwtpE7bsXTehnvRlhoaIDrOlOPk6ROiNA4res
KGbITmeJz31ISWR75iPmgva7h4YdzaNQB2uVzIl0c7j+owkI7xbaDnoDZsBHYJDFmZx49GZ09BAf
Pn0OhtWkJpoTwZxN4dYwF34MDPdfCvC1N+hb60mEORGzEHSY9YULKBydFF96fTkgUpDmFZ0GgGLd
1nNMH0GsWZeKY6QoIOvNNa5WqPsyW+dS3dcAElv4BSdA6dbA2hKDkgj87Su2sXIWYlOTg8IRyyp5
W+RAf3pjkoony4n1TsmwTkCNyXiqqvlnhXBMT4XvbBTph296a+h1dVnV1kmRqV3Lc4fTm/Ry5DZE
yXpZhcexPqayWDdZDbcyOx5/v00Uh1fYDbmZqLhKcoybHGqNCGbiHpzafZ0EeThhXQ3mQqJlS1Zp
TU/37lkl3kZNpb0G8oH4nRJhI7QEBfLhQ20j8gj0pStE2/+584v2BRik1c3VzHg1SImp9d/EwdQI
EJfyQr0oVoCy/uJ8lL/eGv/I3iUSE3eYNNHO2pVL50ZPL1MrN90MrJ01PxX4YmbkETFyB5kJdSmt
A9sGiavHOaK5V2s1gCe/OGGWFdws2vJPBBYKSwb/R5EETce6vjO4NTlGfxsXI1LUlV0L+8CPaAOJ
koSd2hPMUeq+HUcREPPmM/8GMld8pVr8k683Uxx9+mcqY+Dk4Bzf/7ASUv6XpJesQmKoSdOPDT98
3Q/P8vOE4HheQqKCnQpD8HWEKPsmxDN4Ep4IH/RQgEJzSODjYYedh+swfpz8N3Q/M+ZtVnbsqBAd
mtDai9HT5ElNLAx/Qcuc3F0XysLvXVfUan39hyMe6KDTWGCFE8vUdReWALjB7bM6Zk2kFrk4Bs5S
nBXDw9e89kUd5+f4F6ER7nq0/yJe8kT114s86Jh5KWuO3tEDmdPS1mWNBDIRpjyNgXCHuKr+fmQU
VoOjbwE9gNNOB/AfcZzp6ZDMg97zGwRPHqbJtDG8X6i/psRvDBpVacawPHgEYG/lZShY9vpPnj0n
gROSK+YRgl1kddbIeX8N0L/0bUPQDxD+tvZn2k+GuKLK8cfn5na9I0N4/rzQ27IueFxr+95Oit4n
1vdpG8PZ2r9cXCzZy7BjcxQXCmy+KIoTU4LpHJenZeEVNc1h/Y/2IVsQjDdHpGqM852cZdg+fUSY
QWodc+hxdtFPWtGIFQJYutMxYvC9MtXABzCs1i3hE2mSoA2OFScNKn5AqEAtY3YBJRI8h+MqLAiC
deVthZn9h76Evk2XARB7rfVdSRl0F1055gbKxstDSZSTao33fPZaMvPjWitkTG3Bkm1I1Yy2h8Xx
AKG3M2tDurgI4vYPPo/Tzwn/n8pKVLDy1z18e83T/GSkEJ1+1VAxxYi4D9IhlfA4nYPy0ynK76+e
/PPj7NrXd+/izoN0FRBUFfoeiu4JgkIq941QHOeG5aOIw/Xj0ZHWfSe/UDEAuZfOD9QxrjTE0pD2
A6xy71p2CFgkHLDVW631FLb/yz39xovK6la7OXCwzx9mLdjSi+KSWF3mXJZsqAczhDe/M75Jbv7p
E4TyvuLjFhTGcHw64cAmrxen//X9sTxGM7ubWB14wDLS2y5QOrLIkHdUKN+DInQGvwVH8L4v5Z9B
q0SsxlCCuLRQ+NMF3UYw79JaFpQnZOLG0bnSQnFndgDaw9dhYWbXUvu/QxmeZuSP1gBsDVywvuTL
Od4T7wl+MGmStO/rfuEb6Gl/VUzSPjyoybhQYmQ7VyRCZjQ+ZhBJIvumok+CwMp0G9T7VDAwIbEC
9VQ846kRY1uXgl33UfTkYYt8s7tTXQK304Fhh2weKrpsDUzgDPyNuzpABfg3lQFpsEVmgw20+3R5
UBiFm9CVfzZLAmrknwlN71sStffL3q6sBPqMOevWH/Gxpx/1pja6q6yHMzyBmcAlkcfnBhbqSFox
bfF/3w8Zg65ppVThfLAj4tCZUQ+Ecabgz+Bzau2BlZAJOZQTJlAkGbsZ6GeYCPKJpF+eKSqctJcc
Ia6BwXC21W8lhuNb0H8NLzrxh6lshxeNfk5nDDidaEEK6WF8HoFV8POQne64+v5vdptA44Svr3X1
+ogPJP1FKly8lryRGNxD2CXaM5YG/PZtrmJv6rnMCNvEIbigPwF4VXlLg9nspNzNPZbYdqjTL5U0
ewa7k2mlbHwxYv7VuunISPl4FmTHQWE38NOiepdHxt8suWIOiFJmKu2Lk1c1cboh1FkMwEUV/QAt
qqXMaqcWdBAwHArazGyJGfM01Bhbf0z4dm/NVH9A/cEGT9rdc2IFNTMBpPumthh/ePtz1U3tVLUf
WV4CjWkBwF6udorfVz+7Rr2xnFXh+bFLZZk0vvQtqoos8+boPbcW3KHjpkNeN05kOZahbsjX3OGg
QU2LUMd9vb0zKpZi0iYmKbp1aTlOOigjlHtyI4us4ixFD8LE/XzBRZ4URaiPZNCTFYWTRNKGsOIL
sM2XmYHIqWE/ciN6T0rGFaf2l+C522IeFWx8J518DViY9vnW3dHYC44SPNymfnMTmTjKUg4qFPgw
PT1YuW/IITnBszh/Zr0WbYtzpkgmdShGisexntlUbGg5szy1rgIogECG3IwlSbfFMS4Ev9/HkHRW
OEFTTQKGcdVJqIP7pAgAh7wOqQBigz0nyYi6OehBbmR3xKpebbAkQoN+RRfQWjGdchZMCqdwqo5w
mZdpUVOUPDhLLYWZwee0CrVCdGsa2laXvntTLuaUXYmbsWnzjoibdioNIu8SsBq+4DVvGgl4jd2J
2rj2HxbyzPwpbDibbaxE6JtA2TC064JypcXkrR8pePIYOzJzgY7rWhFfjLHNx4YMNDVCbz4tJSfz
4R8M1LKWfbPr+8VP46f7CLgVBnNu6Ku85I9sk9lYNmbID6SF6aRPAByOq3jmUCGoAtSMn1wucRq6
u862O+fNFaDtLOwvQa9XMb8/qUAvU7o1zV6BxmmfHQD3TY+umo8cHOQOE4vGCh/hU8MlW24211k0
29sP778yUUGKxdTjLq42sShi0SyEDoY/4g2mqQdKT0fkVzCw3QJOPuOfJV3Vub+giJY0SrfKSWo2
vAXNtnNHaCK3OuotMQw3pZl6buqPieGgZckktdQ+4UFfF72uSIq0NSXeF94cFWPJ1XTSloR6Q1B/
9Jm8aQD5WQv4X5JBulUUc6wtpN1iMB9v0UvB1bHHGKlQU+CYhCBISKgmBVgovTyNHh5GhVY3h8Fs
I2Qa2CglNb8ilxbW59/PQu195fe6+7iMycdGAHrne/uP7clLoNWVLilBZDy/F+dchy8/2Jeqvj3S
ZQY59paNwgSbYejqYNbu654I4tEASPeeJhgPP0arDcSFdA/OZOLjoRi+SjS6cTaADL/C0a74RJ77
r26niPcSSDy1bumHbOqTlgyALzx5qGh5Tl5ds5+DC/SGG5MOdBDY/Ow8ddTSotkgvHeAcTm4i3iq
wE6tG189WlUOb70i7qEtW47QzJaR50hDtM8eE5d6wgmgsJPNsr1uTM4hX58vgV78/TmI74f8TYaQ
g6wzW0Iy51xwj+4x9zAZOepcg7Ptnv88eFey3uFYGnes//LTmgtknKMCIvqS4Pcc69+wRiQ1tn5H
/rzasSKMp9vrL+TQuf+kLx0+JxavKhbS7Yh13YA3L5ckxC51btAAKc/II1Ldgqkt0qhP5UESoM5u
Zlmqda8BytQLOo9+MevpsAM5sWvnChRh8qfV2O9krSkTTE+vI3wpQOWdHM+pcYDN88xP1S07IpTb
yuj2N8rOeZJ+fp0o1jH7sI20bDcOchBYy8EavFHoxM8TNaNzNnIUoWYWUKPikWc9i+yqkPZSgjIi
fKydyVvyVJ3g8pHXE8XzXkeA8qvtN7II6YJfvaFZAQMFa84h9W7/KhpyjCyoM53gZbW0/bZtsWof
bzhc25wqN6ioNiH0yVjypYv6XYz3fBqJnMEKQNS5x5zS9zYEiANZX1a16kcCs6oPKSaS/rKGZC9q
TuIQ15EKZPVk8g7BY8x0J8Ao3tt6l+gb8ol+2o6475ObpDpsh/JSM1QGuXGZjFlz4hJdgb5I12WI
bz+H+1ebN2GAvzOV0crTyHSnieRUwRqVl/YzPmdGRhYcPk6iEEJMI6CjYxckD63SwX4VfU50c0Og
lrX5BiT7FYvtPSVTI5UG++UEPg0LEEUf0Xl/z3FSAtL8msLut91jrVd9L/yV5FI/wyNGJIsIgCzY
0xYoPLWgt4s9LpKCNVbOKmF5j2Dxyp6QCxmqV+GT8O61nYIN2omIessC3V7sT9JEFjv9OKAv/MyD
gXla8eNGRz0GF9cGoIYPrsylxUa4qxlG0vj8bRZuKKjYpyEremIKEjlawPmwhLn11eXtwVc6PvUZ
2a5wJ6Wlt+p68e7LGYbXkxqG9Gf8hPuKR1OAjk+IoOrdndgP8zkDqo77Mqd3g2fiBPIWobth1Dlz
y/K4KnwXz2/wmacCic+U1g2CevoVAg+54HBux9ivXhMC3J+OGBrUBKXB1NUSBLqsrbgcv0yKE5bu
51Y3cEGRFi4wppHdM0T3fESeZ6J3xhf2DX4sO619Y/eLuq6eGrVXdUBjTuDQ0Z2g6L12r6z4jxz7
ZNMOkGNecjGYnSLAqMa7B/JdjmMYdn27gbVvYYXf5OXMxGTBRuFDUjN8jZSlT2NY1l6A7nHYj2eI
oa4oOwA2PTmaK3dkOwAoZQurcTNHdL/xdDI/2aACJGgg8l6QKlkAiAfomu1B57eZNlIEj2T+Tk//
oFvxqb/bvtfCwKixt1xGSa+2egzp5UNq4+GiMqygR8HM2MEFIB6yFpy3VZ4JK2Aw4G9009bJQnbv
HRhWShwjWUX4akou8kb+YEuymhsQzKqqUzzCMQ/cEIBPx/lXUNGfCfcWaV/gcNsoOQuN/8RFl/w+
tckWNB5DLMNhhaAJ7W+FXv/SHbzlINpemttZfTpFkDZjhpu1K8lUvUEzK5TRYgo7iH5yFo0EJuhr
190gHkyPIIKzkPwj/AbgyBwqPaRHWtkSYaGQF9UlpUUcivrRSNwuVIEDK/FsxNeDf98eqMqLa6TC
Rabnx2Li4tSsUgykPxNBe4B5/So3Kl4FIQaDFnctW3NWH72RsaYj4drKXWbomoyTWfPTbDLXGsQr
vT7SwcKQH2VeWWdiw1rg1w/Shu1dVUVSpK6uyfqmz5Ej4VmY5MsHS91b7la7PE9mMzC/I6F+CQKV
DC80gsyc0nqLBlM/3uAlSyCyCtdZ3KCFJvgXhRUk/5Q33A3jAS3vf4cy+GBtJ9D1BTYCWP0jSQ1S
UuG28sG6KgFhZtsz8OAzeGeorkuWUi66DDQ9rwAmv5T0whGyYqBSJomJZt1je4RrvlzcDYOmzGbY
K8WpmSBu0ekF8EThfx3csn4d/HagVKtZSEXdeIfX0dt9GjFCAGwDUDEcjBHADSP7Kjcw0wJx3J6m
dCDoUktp8xtUHTpTRiPKCmPIRF2KvfEq/+UfX2vyrU6bqCUDy4+SDI0fpXSTN+M3fuNPLT2q5T6Z
EWcS3Lc2xg+63ShPt8xEg6flGUwpmbZKkPh+c9y6zQL8FtMWBxuvnrB9I2cQPhWhD/zJ3xlM91Q7
qMig/1qUGEGHIUa3U/cW9HHzKjx9jVMIMTZiszNCdOYFw+geLfrKVff7GtDU6CtToQCSc7O76aMO
ssE6phkaNLJFrOu6sMcvzk3cAYMxH+iXiS6FEhEPoDdegHV0o6aFPkBKZm9PCVlKLV8ipx/NZz2k
3QV5fSLOYNkQxX4PYIeo6+CGJFBU2yxr2K5RHOcOPx6ov1C/0Zx4W4xaD3SWJF4182xhNg6H5p79
L5h1ZCKUbr004JCGW3YIJ8Gc7jxnJ7z4AS0Xlm9CUS3cmLW0e5Mz+Jw+tzZB4YK+/OMs0bOOHzFt
tkkJPS8CNn61WfNpAKfAbFx3r0+tKnzZkRDWcgITMnftWiMBOlIk39JkUFJhkeXjoqa+diZbQ3YS
9qkg3uB6vjSHcPwHEn31g79LeGcHCBzBrQCOp0pgu8PjQHZuu1AS+9SXKgwaGAsHD4D4kn78c1ko
LWXXmnOnIJxpqaH0nJHi3ve5pZRB9EmRRVJLSSj2HDZ+QJ3XzIok6uxiDv1tWNuhUfy5JSKePFYS
pF5ty4bYG/JvIW6X2kEcEEiNRPB7xWmIYfi2oTGSoEbAmc8rWH87BNfV+Fy2BEylxdY5/cn9IWZ0
60FpbcaC7VTvXfGsPMlzoiEGmPCZSF8ocZS6BbZ7br7BUz4rg3O/w1ZT9PlAj7mQ0Q9rP0ITLPQM
NH/lW4REFi//MfxmUTDZhenPkwfty9eP/8yCZ/cTquEbSK7IY/zjWD3/NtryMbelcq4nUbxhKFwj
42M5fAKAkXsrOQqQYzMybN8i2RiaVKm1CESLmKTNi+ribP//QOxHJSfsvcCE1Vw52xAyKoakH9zg
AkFsuzhGu7tCMCKaPXV2lGf16sMltplmerFpC+Ho7Q120rl+QBN7ZIJJhOM5TPNoBjwB5D36MqUS
f1s1uVxRWmsdq6VXF57kwJnU9rsD8fTCkziu0qn9LpYKohz5MfxIgD5we77FCkmw/ImUZAXjUwuS
cT6C2/aShdit+TiFjQouq7OuoHFNOml563GbxppevwB3A9JxwmcpSUGm4YtEX4OcNdQLa9FHtjjt
mwrcnDCeKH8lCieRsDUCQ8cd8VrziOyw0lnq4kR6wuH9wXliEoqaHPwQTAJZEMF9qracQijq3uIo
mBVHLgQLp1s5weZLLEYxQa+L0rdDz/rwDF1GgAc1VsNldNl64cGU9GuJR9+09eVAZ6K7DBOfo6ci
NvGIawYjBGzqx99t9pDL4QEHgkIJSKC4aawLfCqITMHYHXisNstXejRFOoPwt7fnCfwZEZDHEFmW
5rew5oZ78t1x2tgbfDtcs0EGc1Pg8Ui5qRne8qd/dSXRqAgIzYoTVYeWUqMwl1DXEH9gr9iM8PmK
krJ8dHn95qk7bRA9e77kTPHTvuNs02QShUuZ7dwt0YajiTzGLf2tVRartwGDCt1XKbvGiyl8rbss
LmQP0Vny8a5Q0UuqcfX0Ro3ZQRulZ8NdwJI+UmKhwWU9LQxxcvA9IIk+0Gai+vvUmU8LSm/2rt4r
Q/4X0X65GVatYFjKWaNK1mN7oQXCMUoVUEr0Z4k1xt+bFQogyJR9wW9irAUlhrUFVinDhdJZ6Erj
E4ocHdk2kxy7K/BDYyIl+/YpRPECuuI5lSx+YmNeL+xTS1Jsl3uG+v2UyqtXTZq3fd6iRJcP42Zb
i2San5SdfOKVsfyICyww4P1sgYYGtqp1fa+nC0SbgrI1Mu5CzzD8VUd5emrpgO1DdX+8qURMcQZs
7b/HPFVVBs5aPDkSUHfjqmIGcjxhb+Iy2xLNni07aS7RSQXyvH428kcTUPr3JS9R5nnSKJGmr0wP
jq0ry9dw3+ofNenURdcM1IDEwHfVfy7bB9m82R0d+8DkCjbE3YJgX9Wroa80gMZ+fLmYupN1dOIm
mfO40EHna8u5hLmmUlGrrGp29y0QPM+NAwxY3PSXvZ+JM7bI75ATZSrxzV3sCemzNOfOMncSNOQP
X+JuI3y+Da4QgJebri0hTyB+BgG5z19ZWUciRWrnvy8f6xxr14xQ1KQ9oM3jJJLOZHMr1easzHQo
9wvZBtZYalAOWAvxjKZ4LyVZXEl1SWPvZKM6ZdAbzXxuEoFOb4tXOP5VMtYxfDaolEttDhM/dC8V
WdpFJ2Fe+Nu/OHuOCQOG8pSHFM/gBnmc237iEYAu1jtkDKB9NAQHZIR91236KVIRnogXA2Y3ivcl
O0oxkYbSJuiAXJsfn0X+gT9rpPSiwrsJkbaPmYVG/IEcDub6ovg5Y9FBW5cw90MMRlsRSW7sjcwG
Lx4HXI+avK0I/csvJnYv/Qij8psRWUGzdr8xgLWxlw2rGEQuIKnRlheNAvP2juRxzEVNC51Y3t9d
bNiqAvtu9s8rhLt9dvrR2ydFIfc3fZx6BCeCPjbdoQjWjoY54I0J6Uo9eS7/umU6TzCA+Rmrudsu
EspE4+DQKAZp5v9OEsK1wHBfj0GoYGxW+hdIHxUKEpaJAkcQHNbmOTwFyKRMAJ1vbmPCYlvm/3wY
+Map2rZHMyUmUul1Qu3Dnk8MtFFgooN7J/AH0XOx4GKe4Dyc7NOkwBuh234TvQtqqEbo7vUSYKl8
R1ADAeJHtexmeBHJ3iST955PJpH9Xz1quQaAIH3gGQP9Ofsyyr/Zo08EpU0ojyMhWbJrPE5eNzlI
nPQXXaN+WWnbr637BIhdm7zHp1L7JJffpXQi7WrE2h0JqVbGmrkX5vn4OOL2poV6q7bkmIZ6ZYsp
twmM5/w6tEyAOeBUZSYSVjcfQJfQZzAkV8WiPBNnJYNJ12tsLTRpuw3z6zyagh2N0pliqwFyt6DA
zpV8BSOUT8rJ9Ido9FNaqz0ujt6ISxJ3IcIeYZCktTHXCOV/eeXL5wAMXk+Jmv5/aiknEOjP5SUx
3n6eX1tExI02+05wlgY33wghb6zFvjcGO5P+xplLFGwqmPcrjrwXKRAf7kVIVYcapc27jFJ2tO+v
I/42zNm/oj+KAo4eOn3DWhlMljCvA9XnCRCVir93tbL7AC76G29ftgSo74JrDXsGshC6I09UAY5W
0MW4M/0RbF/mRe/iqk5dUyn+YgewHMCIzuINJo+IhUVPCYDfRlyh0jOD6UctDyg8BeR+m4D+GzeM
q64+sfxUTQaXjR9Nrdpg3gzAZJ4vZWhYV5zvpJDc8ALLZomrm/nQy+Ve4coIve7vC/YSyolfQrsk
xLyQ1s0h8kTwp3XAazI3Yw5LuwSCWM18oLAyrXfeTtzIQiLZHw2ebFtrtxaQNxVRjda9yRdlc4na
ZgP9qVpSsw7NEI2/x+nCM8/x0YdrcuUgIcXffmuM1EhwlJnpSkUuCrh1Rknm5mZBLKiKts2HpLDZ
XlALq30+8Xfc6lNqenra1BbWL/Oxivw65m/1IA8ASdAY9P/WeRAIldR821BnRAdPbvRJnk257ogr
WhmmnTivIeftVF0jvh+UN6y4RCsaePZFBkTrifT3X74+xk9txliVWHcXyowtuIhSzPoGlU863AnV
0DIkgmP3IjN/8BcC+MIfgyDMoyw3P/AHM0JZU0Njo5XyPB6Kk1kknzF/PG8N/SpzDZARxQdXZ1jk
M4xdHDJXebkmGoKKPpTyt7S+rJRAuvBQWUcNd55/HDhhqOn/yqxZr/hKjBQMFBFDbs59rLONhm5x
W3O/bPec50jFJZHCsbqzpZMLFH5POHyIbCaUMYeUfM9AOyVDkf3WmggRosTLhIXWKwAyXNskmZiW
JPhPUpYXrvIoJsq8TMUXdEapeInkmdF3pqCRDt7Q+JmBpY8MPXNRnCor2e7EZviW7+Nr+oB+Dc+C
F51reNUJ5eDFjnqEvwwgxqW8tB82h5CbDN1jXdihx8cqdwuHgmARoapNskRbLmzlnyxXnxmyhlU4
gD2cRqhb7jB+eIQ/O4Oqufr4c9im1gnlqmsUk26mY24N7w35586672eHysX6r/B3Jd+ErvH624i2
zEmrOInw+n6rwRF+IMWeAhJuMPNbW4uC62xku04Bpm3M2A73NnCzBoH5BH1R46/cNdgTc2SJoO/2
zZv36U/pqaVVP9fwQOlP8/BSKF0gwDJ+5ulZF0J25GOr0vMDfs3Lf2ic6oR57U44jEsnKgdmipxE
n5m0Te6/vrLIpfHNTeOjj2WDy+oaykZKaiKRveswH71+knZQ8YHEeSPhkm+DebNQk7Ot+hibywcY
VKGL0D/+B2JjIVcQTQ9n+qJTK32cKu6gA8DtT3f/RzbJ0lF5Xp0sC7uOVZRELEA1K+K47elUA+sb
ho6/6fGRgVNGbKzyZIUGa2xbE1py91hI5cjRsHPdvx5Jp/JvVXBIdAYtVAmBaK1WKx9i+y/A58xn
Dq2ZjuKHqBng1aWRvRTsEI8vlE/cuBLG1foBZFETf29VYrh7p3iDpbNsltSVSSNWvK27unHEOiiG
s1efHuSNQ8fpbRq6zUo04tqX7IaTiR0A2c01WC/ZOQ/f15mMOjUsP3dMUASZ/gLtyA9BEGRnW+MO
pHY9k+ptgjvoWzQn3K5DhjHXcWALxU0Ap2HNBPbZfPafXRo0RsYFm68MY+7CN2sW8kLwE9wLIk3H
h1qs+D310MYYVjI+n241CNrwU+KYTeL4o3w4hRr6fpZrp9Jg4X/WAWyp2AcF6Zgkv/Y+7aIgFwjd
BGQfcQ7WgajI4sx5UFO0o/KMuN5RA8U+aotmFd47icgaOBvJRaoMQC2raBTTMrwzKKXrMe0Qfrxy
T8ZW70xYD7IQ4bWy3/N5jw1hC4GhDbBMZbI11or6QzBni38yB3/vtmwOK4KBeUWeCJxOXsP/8nO+
eMkUF6P42ovAKQG8JlLD1NnaxCHnZvty/lSqqNMTeqOXXQ+Ek9nHL+nAiQKVyAfsPygwfenrO8Pr
Vc2bzP/02UYkkrhDWAbN6VTLyQ3yCgfD/jib2dJIm5b9LQMGVy85XocFsBcXacYjObItP7hMn+fO
9rytV2WrTW0vkq3s813h6sVKwWuFz5D0b0nG2ypuV6P2n7OX+1xAaDZc9vn6zB7dnZ3i2gqrrund
QemuU86+9XO15/i1cjVVMGAzZhrJHZZ4VAWzDMniETCnHitjt9i0245p6uNjFWVDnITHPP/qaQ47
blu4IuLf6wvj57/wentUBmaeWlUx+nGRJ3E3HmEoubEOkJgRb9SRjorBbVtophMfrBDxlqDUTCsx
52Rk1a5N6uBZbU10xVD6c98kqjVjiAN9N61p6VsOBLuiW3uEgbBJ1W3syZE9OIifhxyOUEt6UItR
hIsj5S5qKhbUncTzCmN3YpQ8gon/Z38TaNWe9TorlfY6M/cu+NklwH3M26BYbLmSpzb4m6sP8ryG
g/81MADnD22wuQiARaaeUIyjoIUaeY20Uu/30doP2l7SsJR3/amlSesxc57TwGzH3rKMCpjjNDRH
OVjLCL3t0VwDP4ewhT29rVfT6mIMy+Sz8UCkZpWWBehZdk7YGRjfuwtD/SLY2ONjir2X4ZaBxmDt
F0YnmnK7RQKDY+Ht0JxBCa8bQP7vkVwFbe13Gj8jshB1l9hhUD5hOGKseBiZVAH9Ibgs0DOSa8OD
O5kRB+TX1rFTuJ1Ia5WkQKLha88hv8dFtRSUXZgu7+UfUcmQ39H09FKyVAAKX3iKVj3IzDLu4bHy
Z3TSHq7vY8FhBcOU/vM27S2Ob2UcM3R4qCXMXAI7JEZ6ueBK+uetd0Is/WNBCVVSw6r/CG0pFgYj
rtHwMRstc84ciczHnDeAGsrJSPH7vO4wfexwJS6Emu0jMgRTyvkGhfmIqaF/sDiodO7/fAtJF+mc
bXpNCQKklSqtVqCqpXQ99AZAndcErT+lNgrvyjSp8AP+5l5E44rdYDAS36bbBI4z5cfYceZVPX2U
YL2/mnAQPBVzwHzJ1mrzCSPDCIF/0kmhJtHJNIsXY/tyWZyGVKv7zM8DdVkRU/dWrzl0230HAzqQ
sfCmlCfkU1gNoz029RdF1eojLwtj6PtPvjniHaN1X0eqdpN2ntWh5Iuqn+rnf963AaVG1jSZwtgH
jNoaxJOMjQkXsP2zRM1/w0fOSPJTmKR3XWsqoUwpTaU4CUAuC3FaRGvtjHG/l7lqUqZ0p1a1D9uT
ubM32pQveaCksluswT4LJz8ye9Oa3aRqDNbK+2U5s401YobFDx9Tl1KW+H5OCXfEipfCp+R2W4+E
EV4ADKDsdWcrFLiLygIP/PLh3qDfvpkuioJzgEjUbp5b3TY572unQFkaw50v6BeRzZzLH5NKULmi
QJxZaaoXeTjJbnS+8SV4elxlO5so87mCGG+0hDm6fdo6PGevAoAaeeVH/si4NHLMHiTpas9sfIjO
1GHF1ehMcHdgHOAR9KsObZZcmrXTEH1MD3HKpSI1z5P0OvlxZJiJaO3Jxk7rCb+TqH9Y/aoOaMz+
Vn8jZa6va3cwznQMsj9oD0J5pAkIHlKJpMilyvKxEfyZ7Z3kaXLh/xT9xu5nvBhzoCpZlr8lvGDx
rYN30a2txMu70is7VXPehg2KEBMyNnNzG605n7d7B+0k0MInjwJNt4ZduT+TDAQo7Rn59OMKEebe
BAtNOAPlKCI4fD3mdRwgmseNaInMq/Ux+AK26rZ5nn/N+vWB8N78layGisWx89oO/52fFzBbORYQ
lj5q2ifLpEUSmf36pA3463L+tWbrw3hJ4qaELrMN4ENKrS6215YQ78qefQz5aoHpHE2moUgQsZtO
MTalVF4+W+TNg1ZZe8ufC/3wbuiuC60vBuGOKkfYmtb7L5cxWvWzsndYNxq6STgBtB/4v3ujCO6Y
+0e7/4XWyHgUwmwkxNes9rwiYsbHWFXR2xCXZp6W+JIG68G93AGiu5/C3OU5WDliuY5/wIW00fue
sjUnljvobpvTVzUHROhkTQoOiEJPih6HXeNFfdQpSPZEWDgvCn5pr7kSIO9Db+DkgYSNs0fJ9Fc9
c/bxpCsGkCUuFmL5NUnzaLRwmuSU5J0Rf5fhmdxi5Cei+pHgJB1qkuouUuA0CHq4ADyFNXilWy9e
u5HpOAyc9+ESUoMl8xnDgwtFQHtRpJP92UiChGPxgAee0lLncmQrRt7AzVBW5Ls9NKINSA45mae1
eVrGvOVb9eUU5GvlxVRGGVPGZETb1/Rb1WaP1sItehKEbRJYLoIphMrYpaM5AV7T4eOB5Dx/J8MV
zKAE2CmyagBbSCdyicHTlXGWy3n+q0mbwhGFYl8Yos9fFZL+a+qf/ZdpivFx9+k1+pex4J72TV9k
WKcUMtvWOrJjH77VMSuVAgFU2JRFCBm7YDfVQ6NOMtjA9rZxvlO+m3twjC4AlrNHp9jrmKXbNrnR
NR/64/SBE7RP1biVdl2Gj7U/XxCiBT4qmOGd5HCbBxlzS+ZJH54yy046NCtkmDwOyiAEN2r3HLC7
//l1hNwl6FmIx7db2U5L0fh8v/MnS/qHFSZ6GEg+pj0y3ljnp/WeRqeFu/OH5p3xNXxWssqDgk2D
qu2jE3Nmrvz0uTQ4laQGVpTsfM+SPuikCWSje9Ewwk/0kpUg/yQD8qxZYF+YqLdIFS3SNylnhbH7
NSXc9uQdZ/QEVDJg8aRc+m5yKo2UHCkny+HfYIaBCuh7Pog8EUiPNteCUhH9kZpp8ORGAfw8vbui
pdPTQ/1ojqrY4jJZ2y4hOGyP4TSnmvV4OGLxoglnVbRvDfltbhp6PO7xrNAOcLvHmy3ZShzVeVn1
TQpA6L2SVqEdgAgyUxc2x+FqyIah2wLdhAwnt7m2CUscIpO3xAlgE/tbK9fLTaHhiYRKUPjW/bdp
5VmZ5NnaxQABG/og4RaqYEu4yXW8SeBpPXR4vDLGigeII01aJrv9TiVULZWcognsZKB+CJvSheVn
Ygcd4mxKq0AauqQoSnuor5lIZu9hbOpnF8kkinqCUi0uKKKM4PZvl7OqaTg8g65/YLwbzBLzFN2q
LnjllNofl5w8QEyCR6g2P5F9fu9ivGfRzlmvjD6tYMJvbGYyQLQSY8/oGv2uB9JV27PwKgfPaLOL
CAZKtNvqimxRhJiE/0phhmkPX6UbZZ6u8xMcWTackLNo+JSQMIxdxDa6gY/7z5WYxYNGZ3HBYxku
gSqJYm02/oa+dcRJ1+nENTsmj3i1LCwGS+u2bec2CKep787zBO/1GfKBtOuoe9/g2zHG1mSJiAtT
DO+pdQYraaXserdKA+m9ATu/pxh4TfCPgVFPZOIOOKZ2bql6DL6uCcruS6DYJOHU5ql5nAtZ3Nxk
azfu3pYfVOHjJ4DLwSQRtvwEoIYI6IHyBqIUtLMHmhTWcuYV8JrLIt3exeIDtL/G5JOIA2Hn2wVJ
YcY3lerP7iW4DePSf7+lSBl5uHPTk3mH5EqlpY4i6PW9UvAtx9NIB0ugmXKmpKmGa1nmvamq+6Ah
8F2gkgLyfIFC6swAmMVJy9gAxKDsrkoR/fhQJV9vPz+4WpberB/o9wGas75DVIK5lIMnQ5Q2tWNn
AajiZR7VmM2Ic0q3uG7x5JF7lBpJ9ChY7lC6OlBo8a5g8A0wPxGGJHsrI51fdJziv8Gdxo+rbVZn
6i4GxawmU+dHT8RC2PhivqWiEP9cECGU6+m5boSS8LZbcS2Vrs8RSzLI/N8VBVpFxx6Dl17Xb73Z
mPZ8PH0uW2A1eEkQdNtEFYvf62ihRDKUIBT8Bg07P1xn4zcoYLFDRGhLV0cGGV1uRnbpq2iLhmS7
3zPmBz/z5GLT/Ciu9pcSVHILPUfRTPINc5qMOAR6v/zITN+V3C7Ikc9GdvM3f7ipaYf8Gitl7O+K
Ik1uck0glQAA3lgPiUvWDtWh/zIVgLke/rHdIE8dBvaLekh3NTKmxSnghykgqmz+V1A/sVIvIFDg
Ai7E1q7gs79Ylez4TRvyJogECTalrrT1uOdlHgyv7BsHlcy3YHXfP0azGddR8XcOtMGiB3eDshuk
Arm54dH4Il3WScpgsWl86TMbOlJjlHKSIEi+h1cLGrTrjdtV2edf1m1eMxNdl+k0PiCD2ajoC87b
djlcClqyQJKEItaN6/qUn8JduJF2JTpv/y4Z4rpQ+sS4PE/g1wO/kyrlov4wddZukuH77sRIl9qy
X+l9vPDVxxd0+0qXuBM2QMOSSelTKSG92O17m7oMF+zhX1xhUhc+Cps7Li2l9qNbppAzzMpjTAdj
nwvr6qnJMLvynZG552/cUbuAroheO4yyUt54W/B4YSygGSAuAqJFbnkhxwYuurRd7Tgntg5yQZxo
e5k9bT5PzSUrlXDlQYFfKvFBMNEpE3aVpZyTlMaLQuNfS2eiFvJVO8gVXUEjl9j1T8tuQWmIKhn/
8LRSqXuMrrQ2vKx3mSKcarfqt8BdyOWnoKFgejEMyU59ypNoAkCwfw9Rdtd+Nk4pt6WeUssFjpEi
Z0OBnEIQkcTT5nCDsEuDX81dSECAEMkuxtWqmcf1GFypBdb+IpEw5U1i4f02LQY6o7a20b5V6CQF
9nYOhJ41cip8/y3X0OV2844q0IiFk1ibzcpPS6bS1BX00cIlcqGj9BFDrkDqL7GZyp+ab99T03jE
WZI/I5/p3CY+ZpUAU8jEf8LTMibXlAmOxWH3np+BYovG9Gse4IoiEO7y0f9BK64QaA3o/94niZRb
VhPext6hNSrfjBPRisunaWYmNiJrHE3GXTtFL9q//ONppDecok++aZS7pagaiBhNEurvKFA9xkVS
Acq3vNsuQgxeXX6+CCYikz7h4ugO5KkCDpF5Wrgkc9J7gbNvCVHd+OmnIw72TCbSWj0GsP4A+C+f
HHabYBAEBQ6cIxJ+1TC4RnAwHf+E2rd0z5PaAGiE2y5XSuZMBYICeDrC7ew2EOLz7UDwtO0r4CAK
xT5JGBVFmGUVnHUY2pEc5hPv47fxGFfDh7kpOr5Tk05XP42Jy15lmPwtvaM3ktQD/+GsoWQXH+EK
5f1ImAaX7gikMgfGvxIziZcIWLrQdNQC7fKnHfUqXWY+AeTIaZ7K6n4SEygEgSA4t8TW/hv2JrHn
hg/I0vOskfjVDEFTL6hvgoFMtSZWHKZia6gTW/1yZvHvFUBMk1MESM4IVXSMCYdRFNKX+lP9J1IC
Epy0d46r9ZJjXC8JA5dC9TdClFy6GRfNss086y2Eee49OXUIgu2kxUtro+JltrP6YeIvxqoH3Gim
K+tj9z/zpBStSRTsOrz34YImeot6sk8uFB0U5yY5oPxchdadpTCTLuChmKVdTwX2F0bfgMc6zZuY
azcPqmlwQ8yM/Yipd3yDdLrOen7Vypp0d+QgrJCg6y++z+qFCaUQJm4Lq1uDUj9FTG0+XZIbd/CQ
HexyjnAuxnzfJ7woRfKAYL2slErkUjDiP51geWOCFR+PEl9vhqLwv2GYOGYzrSaLt4sffAEX8jNS
N5EaVj7ZN2EuYa6svFtp2K60sC4ED0+EtIfi+lMKm5FRqgdlLE7JwtbIjvR3LuMJBOiODC8wTuuP
9IGyFbRNd9h1iPWj3fV34CvUGyme3MAuT6d63DuZfFa32ZxzRs6ul7Xoody9NkefMGCuaXHihhF5
K9UGxkwXJ0GzQcqIwv8HPR27F2MAA/m6yaXkGsQubfXIyjJeMlS5E+OlOgLyJQ7ZVSWLMqQx7AF/
tkprYFlrUS97+6tTyQgK2sQEUCwWuYRuIw8pEz6bbutF02GfgO+uaAjMnjtyOrHhHPS7cU/owtBo
DeDbq14Lsq5tMgFCDTDCnwekUuTWzx6ihf2LjgKBOdlqMb4Ojtydl6Dp0Cv142gYs+9+lZdHDrW1
oRqKu0kPyx6wzO3njQYbiffSUiA6erBg8gUfe8QKa86ZJ7XNc8klZ1f09Y4+wYWYsN2qIyrHkdFa
kIJiv5WGJa5KnRxvpTbqJFUNNUZMyIW4shzHXrX7TmYAvTriHnKWntmM3k6D968P+8VHm2zqyFId
chPuUv6ZflKooM5WS2+PmtiK5hNKHQzPxo3ewVFBSYBXv5rvwba4iZRkmdRYUl4cAqgAGKTeN0/N
ujFDhmLVnvJIE3lu5+PXs3RVfn8f0kQxW2roLAZsa6ZywAjHUqPk56E6hchfjoIZpyYjrHnb7Aei
VdBNc7wLbRvvSlTKDmQ3XXOprNu+oh2Wli2k/op8FVZNRd1fJ9hDudVfSDaPzXe9mshyEkL7ClS6
WWYZ/1m0fu+ivYS6MNGErh9AQorjTGl2rd6ZaaR+GH09SBD77ayRsDqKwhjxViTnFPGBHczBOd4p
R86pmEDUipsVYb8M/zpG9HuvKBu+uLl0bfhFdMvzft2ECYzpHVyVJxXcaTl7QDGF0Ec4q7mDnuC2
Ke24WtNAlPEFGemG8CvGJMWvakFtvux+9e9y94mSk7uBPMU24wdoRKCrzE9KcIsE5MoW2yNYQZxi
syz99WwrlGlvD9Pls+AKrUBvpYJc1dgBoTH1/hpfvFV7R93m8fWz1u8ZuwzZjR/703ZDlqsq1GKA
A4S2MtT+YdC/rlBsaqIdOY3B/rc2XCWuQ9q5X8gsZ9+H373o6QQydlioOpQGS5ow6QJH7YRPjAaM
KvKghmz4MBEYXFsfW5Vay1DzcBiHCIiaQSMkmNbdSOPYyeu4EaiM615RQKQpvOlmqW21np6HAH8G
njsLqsvJ0if06C37hs8fYUsfyGss6XVaDpcuesHHEbe9zVmJXLQOPE6rnlPWk7FPcT/f7LfaOVfS
xH7vLy1RkX2vE+RntUBgm4XyyEPx5EYKBBac3AmobPuOWMLLhL2eJfDutiBn9qcfWCLNQ9gzTkuN
+zi9zGRnTzbNwjff4ljzX9JuzXHJ2fJ1Y33XBvjdrR6OmBDS1K+kaZePrLheE1AXwYDXjQPkEXLc
JRaazW4n0Xy6jfE3PkCNUmlxcTOYc61lRdUAE8WeCmPLaV/yVXJvPZ6w6JIbYIyjkIE4lRtOoa5X
ySYRmJ5szU1Hkbmt+vdUQV62k5PHuEuT9TSpQTLotCncAtNGahTZCxQ9s87wI7VtgDq6icS4aCSN
Nd89su55UuuppAmtYumR1CbdvrIHR1YlwAGme38/K4Q7d69S9GXycQUozJBaJbTeKbNW6C/YPDPY
5RWks8KIaZxxivUY+NYetGF8F4gRS4fmC3DfnBDdZFzgrvs4zOwxb/kmLyLjwNe0GGilcFBut2M1
09nEI20J5mNWeMsM4z+H004inbx5UdGMGiV8S+5yixAugqMg3d5S8iTwFxIea561GlWS0B4BG2WL
S+WeOSNJIbdEiuf8R3BAVIJldnsrWmDhGIR6sy4jZvTaoCtPzG6rUW/dktDrWyYJRI3Zq1CD2Eyu
l4y9s6YeE3U5wo2jJc/4L5uw8If5+iioQU0HirVzk+hrI4cLv/Aj+V0vczTHwHCI8PKUUL5GNorr
osdNLyAxqKEznddFsJhJz96wYceO420bn9SSDR9cHCMH6Koj/2hCRR2XaK2jpoL56J3VVhwMXwbU
wfvDfHZjjz5DGU6yCpqvaxkGZXFUPaRE5IKHaVEHwEuuha1Yru7ceszPEoyqWIBV7p/B15JBh4qa
Q5N2QHqb0OOrgp8BfAeyz8s0EfCAbxF+26jgmOSzAM9vWO7sV3qQEXU5VudGR74oyMZIN3ZmZ8hN
JZ9dUYsVFrguZ8b+7x/Uhyu4+Z31ks7egOpKjBnAfQmnmF7ODKFVnBrZ43feDgIVHlrv+0J8jU6j
MD6ctW3gcwRUuuCKit50TFx8pONSoyZeO1xqnZ8QPNGBXunJydyC+zthpvI3ZHpPatp43Qm7TKrM
TlwjxDgEjBXjqcekjaEWrZy2qEQVZPbAxr75i2g50398wLcdFVggT33fYjh1YWnqmSSN0nszj439
4Ni6Gd/Qyxpn/P7UVoToN4PHOyFrDrqvNC1zJs3Tbs6fA+FQimplYTYonsDGZZkbsvkJwNsMiAA+
lApcW3fDqGkRX6TdPjhPdtzp84fAI6EW3Ywt1a+ePyS0kuOk7GIUiySkG6pEMAEYuAM+NDrcp4rS
36UVeOSpTelB83EO/+jTFS5FlCHafTg2xAyr13fiEj9tvfsSXoAkAgAyi4vjKOEO2c0RSpihH3dL
CyH2LQd7jC7jQUihuC6h3Pn4WlbFJpfiPd0JEPtO9O7PrtMcEuUXfm/x5gWKMWcj+v11X41F6+ZI
EcVtT99wch7TWx7TFmv+J5WrZpd44uV7OOgporNou1szcSNqpYAtIF3HImCHlbEvst2VgO76rftJ
+EV6TGm8gFhdtbCECrHA1Ey4jLmcS6p3JvJsaTwEou5RwK5vlnAZ6EI/x9w54kkXbmbsO7rT+G5l
RtSz2IUqAl+teJc1he4IXlUGOLZ6bvoUfN7REQWooX68PO1GQxs8RwzHpe7Dz+BKna5bFpqKFoVE
IudF6sS5EzThKU5wIASTLcBYeIeN88/zhbOmBXWjep4TAadqFIhEgvDLHGmwfD0ATc6shL65gtcs
cQVDJr4EEL/9hGvCAqJQOLMVKFXDlRoAbAyPZImoIlAQ5qAiI4eFgTITS4V6ki+lCFOvRhIJOSzV
TYzw732LaBSfu+zT5Aa5olk34NZ0PLLozFiv0Vf1hIjhEMB3pMATjZANqDBFc2oLDlSlfjhT1+xV
5lstKFDFgc6a3bbgtdp81iM15TeEKtToYuy3ZkjjJ0mvHezBitE5pOR/W2osgK71n7wvMur2CX0r
0vnLXLJqzqwfPXVg2VBjy62GqOXKH7NO2OFz3Us1OO3g8DJk/b2+iOCMigwM2NezFY+1nSNMXtUM
GnE39r4SRPDJTr6n8Y/Fm9k2wzSpGths80w04bHsKSdiyzkJnnnryM+q3n+0bIusaylGH7/jIgvz
FtZ/PBv9QsZ9pT3mD+dIyLeMYTZYGj5D/dZhJRmM3G/dGLQY97KXjMR0aNjMk6hm3tASWIs8a4/Z
zvBpjmpcNg68F7Bk0POgep4ycrhxw1nNNKzpNNnljHh0+lQ630NiWW4fJNCb3++cJdlUPGvuWp/L
dHf2yZC0x+fAfClFdT5HBdH0YHIhLEzKkvB+aifwaWcO1/Is2fuIWOzVkQ4kbByn53ptcSArOXFP
2FDnWIINl4kvEKNDV4LWzTllwPbfo6qJRr8Nb+R5jFqMFHvUI/fSe7Utf1XXRI269mFuVR4NP585
xNU5DdUJ/hI3WNqK3nL79Von5UUsGNPYW3drf0UT6+SZVv48rTrp6XKNb1n/rafmfVgmeOXCg79/
Vbip38OHzFHUmw/utF+fKPEycgd0Zl1hEsXou46EviJuOSxkPRssWnzYveWKSBD9TkjQNCkdWBX6
jPa3p9On72xZK8sb3WEQacjLfH5yGjCciMuW4dMkpMqzO5lZDFrH8Oj+irmAyYJa1JQFwoOHRaVE
iYbgRmMcUPidqEZkWV8+wbWdPumWqfVEwmgCrVoDB+U2HpWAkVc8hSW2niDc3wiwOBk1VF0HFPRO
kcrdSlZm9bDy6tosfQptEUwgGA+sUxII2HflK932gO/Om69s/9vwK2uf+PiC77ekFclOVhdhBFj1
nXAY23RcD1UIUYNw3N10MV4+64UOUeofcge+qjahAI4HFQe1XnQAfLaelM4bjRU96TI21kyQriep
cXPVtHaxg0Wk4bxlVthdiMSRCR6N9iFZvdQwTw7aMlcuPS/6tBZKRA1Gu7ESszwQL98zXDC5delb
H8izBYfmRmMZYn3TWGiw6gGtcF8H43fSeOZ+bsIrLQEFyegtNJtRbd5drVrHmvmdLHRZdHi6evHq
9Rx12zjeXSpnyAZzTIb6d5QWpVnqfG3YmvmdBdNEgxSJ/4tWwRaBQPS1o3GFCRE9d//d7GI6kuRy
TX38HN8pPsn3xkLzlSHvVCLmcR2O5dvv18Z5ei8CpqrrXO2Sw5mFw5Tl/9sJOkeJB+o6RvhicR78
PyDTmtZPYDWnkQ/iY2buhQEQgGBIsicOf/3SmrXRkzSshWKmAjZFicrLpzzamR2yHFt8LFumLHB6
SZaV96KBPM/zOwHWMGL5cevVeVHPoxcRF6odJJ17chIFgmiGdUmirEDFg2KD8iFUI5kVtYQCX8JA
EeQJng6frMGNI9+qbxaJU5f7p3wCDg1msbgBCfVr7xUuFUh0fwjTK78yCf/5zDo5Mnq5/Qxw5iWw
A+o0IjF/jCcSa2zktfZ2R4r8a/VABtfQGQy8pODDFUdQkNGcrd1AxfseIa/CfaPjNaKbzyA6F5QL
pzStsPpi25zex+yBXhQrJ1UCX62eWkL48MB/78GuSzWvKBh9R4Welns/Oywc1zhj3vlY1Ct4WPrh
msPezuSopezcjH56b+JwtTLUDlJ84anmtG210vT8v9QYWhkVA2z4579sNlkZ5Yyb2oMUcpSmJ0Hw
sh1t/Y5POPrCf2dlfGkfB/DySlKig+v0NjdX+cSX/r2kNHZ/pmyBIfLZDBkwgX/6GoMtJx8Fqro0
P4zMxAN31gIzIwJ1/woQBs1KgwnacyhA398kAkuM0T5aaf9r5Z8NO0RVeXqguAoIhUezp6yZ5DYV
DHU0MpszsEVZ5L9gPQV7UUoPyM4lXWx/wHhqqHzqnbcIHz/wpw4ssBD4yvwLX6n0ZzaVlUntqNzg
7ngEXqzYJgnfIFc3Nn83FhH+HyJplZumtZem9gvcTnZqy+LYml+9osUvwucUqXbTZxyTVBdRJ0vS
XXnmjzQVMR1/jS6BNUidJurxNGMdu+Xzy4TQuCcYVlthjWcvw2EASrokCyReSg/O0AtDXjEaBmD8
FV5lYCyDkM66WWMjUQhpptd9oZZ6//geiMrQ8XsTPBOn4/hXkxANN+N2CULEkdsRKv5jY5eINfWJ
XFCqxfVHGixVOkdQMJ14dg9Z7T40/RvzTEwfgrcCLEJ+a+RU97FMAIO5uNaNB815s9JEPhkwSsL7
05+uu4H05YT0lWG5DvhvqoB9LCiHeVjzdUKcewIOgfiGb7T5r2sTTwEq3tOV6lxoNvhuX6Txcon7
/JIBmpYeZ461jDGitJnAP0moANFlZuZnLSW0aB4IWuPaJdKX0vJ5rDfVdyrgIJphALjZfur6IMQ0
VmXdmFwj8utvDMZaNfFbmG6uv4we/YfY3qNIrCn+xp0672ro4++iTxCCbvUtyLlbxYDLrZ0KEHUW
+RTMg7oMeCxikZpDLPbNt5COg/xy9AzjkfnKhrbAxn4fOQo2oPTGbszVFdrfIJH/m+3ujfR4Om71
3eMhOocTLGfrZ5HyGTyY3aG+6rPCnZfbQIqRFM1yfx79uitima2QB6T5Cjcw19byGttHKzuNWdBz
yu+Ygw2zTCL8QaLimdFWRUbl6RCcsyBJNBwHwozT9XTWQ3S9NgdBzJtrzxKaxrCZbeCl1F34sIM9
N1OegT5McKWWii4icCjFtZaa5kgeWNC9cM/lxU7shS/gx7oG4WZokK8O5+7+zl0hmU8fsj4xYu3p
0llhKNQnnDJ5ly36v/D1fULFYYRIfXN+SvS43eq7bU9BuoTePzNnUFYcl6ajfw+jzn/HhOV+Vtbe
SL/JnsDMBk2ack2ZFdk/lAM2kKBBFmx9j4FHSCAS6POVtmFx18CTU/IruupEYRox41Z28xXg9PYb
2Uxsqe4zhfSGpYoV7QwS3qg3fxaRAP1RKY4/r05P81xlRnfb+ygfAfcCUAOPhiym9onqDxaZ2a6J
ZreSfofl+OgkLcuZWGMdsG9/BicAM12Nl4OZ9a+ZHJHVBqxiDNQAkbGVL0vK9B8WPVpoV6SzJ6YK
v7hCMJDZeYaau01S1kOTaKD0kFA1ggnfs7xAxXdtGA7c8JlZEqxRUIPqJxmgV6jrDTaLmGQmvdBQ
CtrZo/BRqJTDIJLvMMrcm4w4tJ2VWYfthwTg/um/bidyQI31SODbvFdLcRR0Z1qfvCc9tKQlF5TS
6v7proXABFD0WCXDhdNjVBz25pvN9T+HYFkqa3s3QRnXjDsO2OlWqEIvGJlkIrao4g/XRmF+cbnT
dugFuCl2WCU5MU9VhD43dDf9jrykmnnnSWyUsRo5dBcavighlCDTT5+fO8zKSk/jcxinI+npNcua
Lfi2GDG0i59ROIdIFNUdVWAFTlPGCLkr1+RWM7InWb+gWdM3ERHegHMHZOCaYY2G61YpbcAA/ZmX
AZ0f+2F0DgeT62pEZxz69rKXJgKKBgPJzGRKEfYh/WADUnVVcFfw6k5kPKwf3Z0gGv/c7CkY3MCW
gmFLcxglscCQwKr+5a3t1n2yT0MGzTPiCaMSrJEMMpGQN6Lj/Bd5YD3P8S+Mz/bDgp9rpsiy4Odt
nGecNv2LZYJi0QvTQMHsbZYcCNgKdz60tl7x+VnbxDJI4EHzbF0o7c9UqWkt8BdZdRMPF12PGZ69
SCc93JeB5MGbAXw9bW27nAxTd9jbG4shqRRKpJocrFghYlDE3E45+iQtXvqhAiRSUKO9lwaCHH+Z
dAxTmVI9VlhhlfgrAYECCuhzH9q6vkQQijuBUVCTjOF/EuPylW0G6ReKc02WIjd8v3Wlvaoeh1XJ
T8aLzQHCJQOKyUD+P4RWXRt8ai49Joj4BkbPZJpRRuX6fE40Y318/ACQSQTLoFauqvCnLkn9U+cz
Hm/k6O+u6VoFwHdpZECQcQQbrW/z0feUOT8ajE6o4KJw1H1F7QxBC55Kvcd6eE1feip74Irvs/u7
xrPo5ykan66mQ1iKpWlz+QNH3WHD6fEfdlcm1lZG2bkLkLyhwZmBN0SPgHYhx/7Q+PBeWCtVYRDD
jIwSXwAZz9aJi7nBO07puPveUiLF/mXy6sjRLKAq6SfB+wC4WOo5Humy50XvEcgjHAtOxrdYzXaL
7Yr4f27mS6rGQpRYKs9L0waMPJHhZfiBgaPX1omNScOA1M+rQz6XaSwK4gtkwwqsCixdj3Q1Gw+N
nUx/shPVvaq0UKqcRanVEIXQwVTLVo4aluPTnWeXSfQk1cahr6MOb1/MOFGM/jvQ5dt0vkk6eWvn
78tnCl76ZbJuKbvUt0GiXGd0k5OJg/SH66Rps20fPGOrim8Xd5iipQoZhPbrjAqxUgKmhzxgz0fN
F208ysLpDu/B7m6ceX8wwxOFsuNci1hLsfsWVZRG5B1yQ0LWL7CEWrm5yZClRL6ZkVrf5YSCOGW4
AUeNbKZaoMbLO9GkL8YqyuLWD29NpyUI/n6/Zx46aKI9ILLMIdnkDOVU0La29rpwK1Q2bFSQL53M
eAf55uC5CVgS2a4ZsyYyfxGdzx28hJqADyeDHbP+Y5sGatr3YK3QGwN1lC5ZbpeXBfjzk6y9Xpc/
7V/1+YATtxO394CqKuS0yaVPbXT0M+ezw9sMyh8hNer5ARJ/53x/mCylFf/AjGjIcKW2KvpWNJ9v
PH86jIQ7mzfamfk18rKf+S5YWfqdNp8x/YoG5KCmOrLTsjhsFX2eiJqSU8W1vX3Tk0vRMsgx2Za3
wo06QvdFleYUkYqJrin5AAvTioCj+PSVwGK4d4wplSzPpBRWrFPIOZTeuvzvhsqXKRZ35oTaIzzy
S5Eu/54PtOwRN8H2bVuYdflcSSZrmCsAFzc8kiGxRPzlAjeND/iTNlCMCB0Zs5VBR3twh0yioLJI
G71OcZkK7LSd3oCYkvVY9OrWpmIEkhSfDMDIAh3nnIV6cyy+JxKuXYIMjkL95YPzrYCVUIRqDgTe
VjvefUVCpudx4TFwFxo+Ks+ZRdoC7oJ7DV0zBTgqFV8fSmYvsOXXD7ot/oQL9J3OD9JX0fno5mAe
KbEm2U723Gnj96iogwM2SZrksD1+h4pk8iDdPsaSGqr+46cPg0Z6skIlJrN3uD8kImx8338WGual
2yURnyE6NoDRO/bkmmKuy0zu1JbhJAx71f0xPtGZf+0+LoSgzFzH9lZOn2Ey/WiU5lxT5Egxe8QK
Eh6SJFjlZkOHhqsZwlv7qaOALW37bhbiBxUseirzn+hTdkQTtJUEmHcaaoYwXZnPMX5YtQNJhnbQ
0mS+IthtnxW0f4bA6w6DQ5aWRQYnvCYdXm9i4BTtduMbXumDhRjL/92mW2AsAQ3RnJwBkctxmWQY
83dFCozsx+QR8H2JgUPHDDF8L8O977EU4yvXziifCNxKTxMi00Z6tGcAfTmKb/PPbA/Dj3p15vLp
z+GmBU5y5n5ieK4RQBou+whvmlDU50EDhLhgtvQVdrePZKkIoFDQk8r41w80RwvPiLQgF3w25uUu
gTTR8r5FFUsYKhr9h0ygi9N3vzdlfuHLq/fk4lo5TjLDnvJeFcWrEtyNoaDYxb3CqyGw2j9qklVa
IsxCmu6Ankn2qtgOTOygGAM0VNS2ak//F9MhWzBmCiVQNrWcjXT+tLnra/8WCz9VRxMjStnFNMgx
WE5yczmNQ9Wb1E6LqP2178S/vDy+A+UMYERzUEQ0LV/5IWiyyKJcvK3A3oEzUPajGCP4086k4EmM
7VboyozKxta0W4oDwP+H8dsfgjXgppaDvbc4hBbqDwyPddCmBPpXy2Cxd41CtH7Fet31R8Ez+7Gx
6AgIEqcfFY1hkzQQZOCWPAD2rrou6suVQCyeGq4re6AThUJ7KF/iN3o1XpFiq9lvy1FwvZV1XMuo
EhtViq2jtXmWOZYDiodwzzQAMEieSzbhQUXaIXUIAkT6JJBAANH7XF/g+VRx7g476/fhOI+RgXKj
dCPf9p8aVmq76yWmAldWEzJ+XMwFpwHrBNkTzRnuYzcC34NEXkC/sRvL3HGnik+gOjLbacVGnLLZ
kjvw3hHiPqSwLClncTS9skaKn5ZUzX4FMJxKevQ3pJ02CYwAZAt4W1Upxkhc3d8KK76hD3dLMscd
7bzInBICDoMulDP08kLCjFnm8He4wc2YUq+dEeUiMsU+zACRQfB0P16r73iax1LAI46sT2KrX/s5
Ok5N1pvlPUVo+xdyz4bpVQ3sLFJGOUVdONVhZWDcPOP8tKfiNWIDtbA6OvMU7pygqZVbHLJ+Xizk
Z12Ia5qdfD0PPSD3HqYbqckRSYgcr259IHJbroefubpgElFFfNGGsf5jy4Hdwy7XFKybgNZgTxtQ
bGfRNq4/ondbRYDbfEGJ+FKvaqh06VHvee2Pu98d6v46OI9EC2RiCASQpARnP91UF32DNWtH8y/L
ctUn+j002LjK26WhiiIESrHV6GAIAcIcGOJxod9OPBDNqnMZ1GQ97Nnydm5BH48vH8dxfzOBYViT
O+Vrw7ljy0Hcs9oXTvzLOLHfEjg8tucOkoORAJH0xkjCynTDCqtTyEKVX+3N0b7pt5zQ03kGJylG
TVMAXKgctGG3+P7mX0/FAtfjFjbwZ0mJgKSIYnyslU/Puw77VI6H/9UAzlTFROBChuOJwrYBAD47
Q5ThRl9sSrZ17AyHciJyQgKrdHu7VZgpk/mB4XKuEKAqxaWz737T7I3W6goClT9kIkuEsirQv/IA
jHia+2q3DHGGxAbKQuxK9w5J8KesnMVJRRFrxiaH8hJdaWqw6Hr8pVBzB1pilHd1E0tlGgyzSolX
3dzGxbRF6+ZEHbxqr57/6dw40JIwuihExUhuJXQ0h7sFKq0UzfB2fI+39MceS2oD/XNxntZKmCo1
fRJY5S8dM+7MxuFzMAg8bOaSK8LrjsXUPby8s/8WbhJYvm3vpeVUuH5CrUErsT6SUJNTgtCxNC3k
Fd87ZCoTbO4k+Rj0sFyWSAzeXQ1IF3EiLIboGNPvPQGdA66BU2jLp8G7zHPOaK4L2bRfZV5LAhk2
CGdzFOjjd2qI/1+hq8VkcDQyuCgWvLOCZk5NSj+eKGEUkC7Q4KypiGtuPuwrIPLr5xOcYj62RxTc
Gxx61OZVbAJMSwQ5qZNeXqQigRRABxZsEnro6zS42Hr/epAFL1OfjdPB1cNWS33mNvre8gjDo9Hm
1h2kvUe/Q6hQniQfDVilTcVLfLmBTWgbWYKKKywfJhIJM0r7b7ooQ0KeHIM2DUb6JcV4n+3JBlTa
C8MIvAU1wf6/frMArJBHvWGc+lT4i83gURQ8RUZFGGpuC6uzZjBWan//7YqnW3ZKoUvucxMoldje
Cz1xGqTJMF2HWXpqsM0S7YcRJlq1zOELTLn6a9cjkjRrkkHBKKWRMRLiFHGPZy+6eIEXP1IGy7ya
LCZq6wpSE/lYmVWVco1UkQnFS96tvIspIF145MdIHYw1mjdNYBuHqbjYnLNiyaVmNuuKguGlV9BT
m/yyKt3/WAMlRtlI6Ow/lp1B9JSToQMW+jvm3cdP87SNyPXv3J/ceguxScRG6ehwDhCRgZ/TK9ar
BM6ylD5Ibi/Y4ofU4+wPuvvEMJdBMGk1O11no7B1ct2Mii2AMwehy03TkscWOodVuV9jP4jKYRjT
9d6sBca6VR3ygxcYWH9epS3QWLA7BGg7JO4Rqj7QDW4yEY9jQYi+yjUU7AqPthlt1Q7TXpDZ/FpQ
zx1OK7HzOvSvWQ93O9aP/JB4g60N57d/0GYbK4F3G5JAGY0pPlIBEu4VhGnfb/qLUxA0e6zVazvc
pm+IK9SESTeGJhwfCuyuGnSUwA1CuLqa0kshbjkUuz2jS0T4HfCCowv2ae6ICHZTgpMwxgkxuBX3
x6KouMkdQXOjBpmNreY14SMV2jmW8IABhLbjY0sBXZLWiFQ678EZLNYzExVZuhTAwTHoM9znGXZT
+OeoR67w8mPaldTzm4jiGHmqMoz3K5JrQ96mgXF2/xc1wZLGvI/Lf1lPaMQjqYTCd7mMeYRhlhAY
PLXfESf00ylw4DVZwpSE49dQEk7aMtJMLIx5/Zg0nrCggN1kigT05jZaFQReK+XzQDoXj4RChn29
EOFoGmvjYn4qUiou0mHoDWFfh1MZXvUOt+jdRP0LKrMLBgdeCrFDszPUdm4JKJcFW9DsYkiADA4Y
DTfyCIxS7fMm1k/fqDFUlHl58tcsF18CBUnS8J5o9xwF7H+PEG+E+MIzBc0mT0A9Mh80tpk/TNcl
72B5ApD7mkWxMU1ofcfMvqoZ8fEIvjHPAlwszp0TxDNP7wqhSlUWbX1BtyF/I/GuhYWUUcnmcve3
bLdZXU64/AJ2RaIAUjAiCpg3B5gFESvS40mUm59+UXVT6jHxG9C3baDQ7QRHqXCmIFHqVN65GU3f
jXPs1H///oK3JdDisGEyT3R9kc9i6+XkPoqh0laZwGUw0vl4wvCbvst4oJJ2hukYU2wCMievKpFc
Mav0WwsKpeNMdcmq7Q7ozjuZl8+SUi7BkMWZvLFMbnt5DAt2ER5z/CSLBeEE3isR+uluDcwa2wbU
X35s7SZT4GQ34AZgchhZ+a3vTt/xOB0mO3ZifESMLF78CppaeYPgx6OiNgcTrbFCJJGwYowp/QVa
feqjUBKQ5PlQ1QbxTutGcP929GXXB5ZdZTnVic+avsVQWUuvmIo3DFusD+iA8Qy+ZJh5y66eu2Ao
vP/9nuimP636YyKE4A6xEK5JPH/McfZzuqEZwx5Y/oY12NLxBfwTLctn+azLSaTXFMJZmhOKykDA
7bFFMaS8vH2MMN3L8n2eneHbhOMVd8WqiwZ+x7Op1ZEmVuHseQ+z3tfEzq8uapYH+OeQE7BIOzOm
TtteWpEhV0pyuzSL7CWWOiekSiJFWtD6UAucdpccLCJffgAQU6q5iwL8zH3Wukcz8zK2dpWQn7bn
0NM6T6wNymJZs0VNtdVqn0qGxJZv3QIAM8wEK8jVQBheLNDbUlyQ4ZtqRbji6E31Fp6fFZLEqv4T
JtX7zbLLNcNTnzaf2ZEgpVZthCbDVpnv2FV1JNZ/xnJpU2Q0jhuNBTwLHOl4IAgEMfkeC589YauQ
0g2Zkj0W1l59VRO7CEUzDfPOlsd3I7UDSOWwMJ7bp4BlHvyGedzvhnQyuZBFxi1awdEDO7NjzuYQ
2BwQkyneZL1NGDJ8stZfVX7bJ7E5PnH3uB2FmrQleLQlBp39H++Q9Cuur3+6RzJh6Tdntqk1+4Ar
dUufjyyNy/IabNvHEciPHBgFHDEsF2RhV+hqYIfGgbZP7tbsUVXDbj/i8wNrbMZmFCRxeUdkkvsx
U5fQlCX1mOPLRsn61SeZ7Uf7x/B43F3ZDbkGilt3ir7w+dcqnFSzoehjcd5mHgdpHmMXnmwnNm3F
iW6YldVqeSGPxrQMezIBoPI2uWBlGG/NXEebHws3M7cl8mFVJ/ARRlqWxdGUyCnGVmEmrvdT2QFA
UD7LQ8BLMbJT2NrrtAmSCNczG79dizZfnnsLACRlfJe7RxNeucE0+xWYUhOaMnQ7nM8K0LkRSsi2
oK8lcZ1VZytVYwOohcpFooLZTDcWYFGJ0n/f4CkRIY+zYCaGHhpi/DuzcCtJ04fbIai2jC3/PP0O
IWELpgDMWi//oy1nVeTWC2whv3Zl4zZgzfq/NmvM6dkJGjHXyD6QRSB703EmkqJrdcEZqmhXUl9T
yU0LH/6qT0+EanirAMdOgGiGwhpBdpQzopykTum5QS44+nZBX/6zHG8W8s+nZnujiK+K8XSpNaji
lJihTGSw/1C2qVnfwkdF3ymR7Atj/B5KUqVeIBLDSYmfizLp57g+xHg076C50N0JxlIopjPAHcq6
XmSpuCGSc8uSrkQOH4bqI3/IOu8hazHz8xMWccGLjYr/rUmo7sZSSjIbclP3sH1Fzt+A8It33kkM
WlZyTLIsQV0hOdQG5UtN/aWk3Wj7JXDlmydLLg8tp3kP2qfWYuy48UKrCbt+PnGcVXcBJ9lXjD+n
If/mYoFv6B7Tb4TWCUe30v1UxZsrY/PR8lTNhErx99tZNOVmuZyd5MiBmudi+Uxe3R3yJ6/rawIh
YBRAa3dblHPzMGDVFcSd2Ma7SbB49lpGN2reGsVgzN5H9X4qcP5p98IagLtTYiUGHtOQLAMqbMv5
KkWEActLwBlPWNEVx1x782gtChpNu8d8TNMkxkvQNY9PzYKcEAHBk/m99K7FTV3G4J16HrX20uvT
EFp5XWGOpO3ey4bnTkVTvddrc6vgaOtO2hxy9wPWPBblsjrRjKkeOlBjuNgKrKJp7hsrL0rTG7Ys
Odb9y2YAjrZx2P3TAqP1d5QkjWTeye9E4d9YtVRLeQJHNTNW8fBRbFl3AShhTYZFHnbfbl3d0N1u
jmK2Txmyy9wX55L0d8FUG+3s2Q6EwQj6GrTila4WXXzOhpBYmrrxZLBMKWBbqS6nmnqDkAIANRuY
sKu6ZqhDZ8qVkbMfrKwJrd69MvG9BElD9ne88sEqaunpTh6y4PGBe98wCN7FCqcVWH0zyU0LSFwo
FiJwJq+RnutA+L7bqoRL42eM7WY5VUQHDayt3t83TK4jQhg+k+qtcby7NSQJk90IINzHvWsba3pr
HRMEL5LDr7JQ31G8PkzVnIeTDQWWbbFcfMQeGld3beJ4PyDsNwmwAT3mkTwB9+h/kG+Am/2tTtXM
xlTIrdJlhUQOeCEM2MOCtTqlB51UILo97pf0Z6R495a5rP79+fuhNveHrYQBncO5yOQ0Bf5EuDpE
+/W00UQY0wMRCBCPq1GJc4FfmkTzs4Cg3EOrU66FAAV/6Ga5RG+Sn4tG4TSJUCN/jd7ibvI6IAGK
X0GiB4taNOLEkerZjkkXmFiypuM7apVNlT/quxfpTLonYAT9sZbcR5N9btxzkXgkarTm+0ksTVsz
132QEwIyc7cBv3oxOHVcbfMpEEA2cPnxAgKLWvJNssAeZvFQ1vey9JsFnyBizTFA6WFOjZrjUVMU
SFyhWexfqJU3aQq6wlsfDK2nFKvmKvbixnuZFtmh7cmVPGpNX7QFclOrAcJQfLYDFQYtj5Dt3T3V
U4DerWdT06eS7G2z2vmdt0qUllgFi2Z59zEu4dRyrl3WcORN7HjBsWoWOFyO3R4kpeZaXNhUqxWT
++G9nJcyumoIq5/1x7zq/NvBT2AZfOHuK8kBewg+7xI/nVjPe05/caENhTOC2dwYWLhlq0QhxRgC
QQ++akv2WzX6UEUgSRuv6WC7qCM3HG29KHbRF3qzzWaLG25hMCqTqzT/kiKgWnj18CGWaSSAljay
oaKTWwNQtwk422l1f4LJNpawWTFolU0FMAvxHgr+nfuI+vNrXUMhvsauji1p9nEYgoxDDknmwnIK
QYMemrGxL0r4ZzMMsIikXudXQ1OytIX0mNO6Z/QRyJTqkJl5li5Hmr+sv9a9UVA0VMBFrEtQirKz
8P9h452RzQ+ifU6rim/3kvPjNiziPApBoyE/5MJ/4F6xJbz3L+Lv98e5a/2gTzcSqA5g6C9hnXmP
X7GVq8kjpWPpx6pJR09V40jJMAkSZFP4R/skcO/ZENZyf8EfyAtZjsE9Cvz0oKHFU1N5hlX7U1EE
hCIX7h8mUTvEpfI8la7vcWOh4PnY8iK86AJhJ42jGHqYMe3ygrPCxe8TfymA6GgBmpVjq4dBmNpe
B8F5U13xIf8rlKNGEUxxAVgmtO+qutiLBI2RSYD8CP4mEZcfBK5rDrQJX0bfk2uRmyiHWiplitVz
5a1xvuvbzUyOdhqbVCSrsEH9OORE/rrH2ywpHpJ6hdnUKCKf/xqJbC5PC8VL9i8eXZWQcvyH6o/q
yzM/lP5CuchY0PCJu4CX5siigMQsZ4ffd5xTDxP3fy6ykXIE3f5261130SGWcjzPypU4MS3CwxzV
PsSHXAA6opuYlMwC+ucNsXyBJLFbnU8Mm1+OvxCz5TzPtPsMyrld7Cuh6ly/q080oP0sn5gNHnjm
8KGT9DyzcoFHj3B46+f4YToZrOk3nF82zLaTngnr53t0eDGay3GVfpro9WLh9LJUGlTcSvzxc+Iu
cpEjCZ0x1gJidBbpDrDUfyYoCj4JiIY+KwOJYbg/NfDFNCZSOu6s++trBRSBh2Uj3H7AYYymo47n
HnXQvxIF2ZlCw13pZ9iTcAOaSvPn8F284siRpjRkDRyTeHMZIOH1/8Ai4uJBFxCwiLaf7tRf9G9W
NuuoT9Mc+C8Mw/4Cj7GYa+LWENZCqNqWLQiMVYkb1XCUZag8afz9VzhoicomvfbA5zx0YkOr560y
IZ+Tu+Mpis7OF0TEwa6QnpKLtalRmx1qlAlQViSu4A+77//qCt8D0wxZbaOtsTWbQyKa/vfgqJqz
A3YWJXvCwf37s4Lu8ezs0t+lOEbbABoog7kKv2yNNMdJk4ghrk1cprzau/FzRZiCEjxIhFpVbr+h
4S+LbvlX4EZ66CcPW67b6GwI7zZLKRpDiKxRLhVA3DuifM5NY5abjkusoLtb57zuWIoi+R4TemVU
Wv5B9SQjenR1ukTIBncpwszqaoyLaeDSrm7CTDLQN0oAm0mQFGg2pyVN6bJMbHwTmCo2caeiGk51
AMxxKf3PDeAQsrxjT+8D6gPCupFyf8do6oXNUNCvhe6m0lcLhi7axG4V2mGd5JFFsMY6C5qyoLM4
rVNwGpGYZG1voZ4mRCyRvPbpIHDFM9fO+1cb7JlJBQybDqbDPgy58Bb2rejMT+Q6Zmp+c71tvGPS
UP0jdtaF+cnLV2N+l3ncIGiqA4++b3XCPA7h8kpBPmuRjrhy21fcpw6M6+kIIh2IpYjKkHNHwaZi
i/FL1INyH3tJib+2VNhhLvzoxLpM3Hkrkmaj3vZK2iQFD4tJ+Y28DyVUOZh6+Ctp/ypQFgkmuGSf
WrWeSpj2cZINVwILmos9sbCXESqG7B4M3b42I5bBfasZfw3G2BTHGXsKbN47qwYxl3S7Ko86QV+B
lJ5EpoqPW2OzowuekQHdyHdi2T3atsK7Ar7Gx9xLB2IdKV97fQV/0uiGQ1AEzpDhkYhRu+IYdmEP
ELB1ApvaN6r6084LcaXxVCOhdCG3A50iTszqfm7HETSPjIUvwxF6qbQF+21sKVcZ1Cvddj2PE1o9
qzVDqDv/dNvDMRnIR23C9qXOtbssEt837ThgFuLFCAumJaonBQXClfm+h96taDznBkE3JqD8EQWT
9OKBMwRY4ao8V4x5s77zQA1r3Zo2ApXLl1Kq21bQhyk5G9gjZJtD8Ao5NeNpzxQu7PeyDKnhTBpz
QD5ul/ltg4k14iKyYCi6gZ0n0XtCzKhDVh0RTDlbVpaYjQ+NaaKDkPk/X0sk2pcAw/WecndlnHzv
7hT+Sc3gB75B0OT0GbMGf208CzT14H8J3VSaiJLXQ5QsabL4EPl0MizQVg8aYoNk01NlfAz2d0ee
3c/tW4EY45X1fz/VP5TH8Wk+2+arDX40DNzxdp8muGi8Pny7KryKo48N825ueTijzegdYboywpDa
Q+b8VG8BbdUB6ohA/sJFaZ+hntPV7Rm+mi4Tm+piu/th2fnL742LKyFviG8AY+A/+FYiNNvYIIff
6E3t9+w6hWzXRgAQHSivrS+SV32+PNOL6dcLtynWcuQ06WylTq4nWAK/uT+/uPq6UNKSQsOEKmdQ
G5iyWObjHH/732qIHpqOB+EEm28gqy5txSphP4VTOwIxczqVAnyDbVfJQKNdkkSPuLu4xhjAhRhi
maRSTs78/Ysh4W9yYrlgL/zto7HS3SKptSVwry8IR7xUuZNuyVfl8oSz8SK1w/hUzX67utSOKaQP
MQfGRpqJ3e40syVeZ14+dXrx4/B7hJ6KGJEpB3HK4pShIv5vwXycX914IQQCzrqCfkI45X/7A9sC
lntxdSAodYjx267Kq2QhF5/tMZxCFrbs1ksoYsMeazEDYwynpqEqTV4pMwQUlnL1tTIN2aRc4rbQ
ZALIt706fUiEiM0NCAGMtwyv5lyPPRTiHXHkol3Vs1e8nxSWwiFxqEoknMozo4jG7RRfR64BBKiU
6yRTLhXuvvs6KeW1xL096I9C6qI46vRXQAY3f4TrJfUNuBE7dXUD1Fv5R/Pvqd5DAoiXOJE1lRh1
G8gdymlpqnD+bXwdhh8FLIh5i3GUYzMt6FOQgMQ38nuqCqp6vT77Drf24hlpgBVwYFvxsAR/J4HG
f5wdITyBe3dnwc0YlfGJUafs3BDJPizBoRLLZGJEWd+jrwQj7hIwfCkM0ahizUqYf/sZlmXj5Bw/
P2e6qGi02TLn1EjCA+RjRSUkY6mRSVZrpqDy5gFe1yxyjcYNw/voYlCTc7YPP3VeeTp4DLG1h5GH
CVtlV2fb6/UwMmTJaeogURyiJSY5vVYjoF4AAj+6ZHJ7VV8pMzZkPrPZSQGBMlfs/N0K6Vq6Pc+o
BvZjITFlk69I3RofmuOi1MhUlpEPp17zJWRDH4ZKTiey1s4KHJUJMvnZG9DNGdyCpUl8d0y9UH14
FJbu3ryBalYoV/QjcBgKuld5rjeERlt3aGKb+jzH4ZdD/2CmnCsdPY6iABpSadZNYbsKVo0kMvoL
T3vSTsF0WVbWxx4WS6kUlCD47DAyJUe8pMGC1KyjDJsD1pnMwZIRwxy2M9WglsEtdTBtCEdeft8i
hS2CSEBjxIASjWI4GDG6lL4GJCvcKK6UnTTEbZE4g8qTSO4H136gm1EVtiqICTza3w/415Jzpbzn
29yMDTE0xdAlwL5+1+7YR7akE4a6V66b/MWoZLxov3E+GPxes1/R51SOOif1iQmSNetN7B84+1Qn
gIVthup9dxuU4oQMIE06FcqYjgw3/wpq+2emS6X3TxISQdgsQM4WBGTBPk0YY92aslRxxqqiLZNC
aIH5rRwit1g50Hy34aJu+NRXFaNzVQT2y3RoZj2xIl03/FPQ3uDWcUKDXVXqRcAeQiz6VliBkXYo
S3MdOeDDDpwqrIMQ7Mlo3EYQz7KiNrxUIiPyqtsB7iQBZ9uLfTkk8wXzTZ4Q6q4M6jkKdbxWWDpj
J282Yw/NHwFs5ZAvJ1NIko6s4hIoyn9Quy20PaKDmV0ZHOObdJngGJqJ4NTlic9r0H2XkGSIzpXe
K6JXKTfS7GcmQvIVAXwYXLtpm/hDb12EzIYpu8aBnnMxqPOJABt3r0O50w7gHbmrip1ruExfXBsE
2nXs6tE95OOJcdRSRGQ3znJICaWv/ere/aSTznaz62LZhZ8fE2uGZ+ASh1aW/4NAzPbXWGegrmg1
imPVqghBYi+P6/uto1Pre/nSUAxjkkikfzy7NyWWw8bCM0jIkAXSmxSVRLsqQO2TTSxOxV01MPAh
xvKSVcI3KHi+l/zUWOwszopjD6xF+KNKae2iYydeEa6+ZjC3uf+YxQZYWnjG11GEzBxbemRAbrlW
bgArQxhmfFc5ulfYDmzmJDNrR1WvA3TYHd/jd3PkT2yQP5J12ns3JCvgbF13D9gtgyJO/6lynW9m
ZbSdDqzhdByhXpLp7H80T2ansCPhfSJEQm3hbqFQ8EHxSdGYMzHQTVCTiB6ah4Igj4twNhowgnLj
RXNdHO9t67BjIZL9GnlAYfNhBQC+oxq9bPNj3xRc+NSFJWcV5qPECFXIyS5+cwRbjN4Gr9LEkWQX
NeBOanoQf64qeIaZyE6rlnH3H4HbcrboJKj0uxB710CeWGpQ1BRvRYhIlLCU04SEpB03Mz6epuJ4
HebjqbrmHsh9fbbOrl+RvfP5r3HmsneEQzrgkQ2YTfM9PMf5JJLgBeP8TltzhFY9Gu1lRXOCSQ6t
XagLgScAJQxwoplQ7eIANXyCYb5PFFh8ZJI9yfai+CV2X8JkqYS06Jdmt3xa7qtV/RmS9bHaqOv8
C9tyxz716kSS+sK5/VOLUKjSExngmdt3KgacQybmFPp+6WRR7NlQPbbrR6UkmVzRvdd9FwA/VIxb
EjMc2kYs5jRDTsKxbcoy+XV+HNdfDJRe9Pdk6pr7k13c7Io9QSoPCqMmURSrqMk8aVW+A4QgWNST
0uh1tyEGk10xnCSLli2z2oBPV4Ck8WEOGpoRVKSYi07WyakNq0JKqP8CZuTkspP9md182OLV8HSZ
o5t7f4OzmbpMUDVan26Mf45UhXgy/oBXt4bbquRbnfufa++0wU0Stbv+hM+Xg+xgAyUEiD419sFG
xp4OP0I4uo12PvyQpcu0Q5jjQTf1xiB/wUTREG5J9+Fm5uEk6oXHL8QUSloA4wQc5RRh0CyEgFJX
9iDiiYzRz3yeecWNYAF9Mpgrf45SvSUXuOmrbFEy8SHk58QuiwjqxjIQDwU9Ne92GR9CgRBEKEC+
iBRkkhbS9ATHQp0aVb7/3QEF3IK/bJduOJHzwkNqofSqYPfwpbwB6H1Pau+vuxy+0aVcxpR/cph6
YXR0woKWNSewgbDUNdBGZn41g4yBqObqB6183OWutoU6NXEbcAkaYX3GPVowT9+mJbgvLblX132Q
3POiEV8Hcg4EMhmis9F7wDQB4UehA2JtcSbTI/BBQMkvgOe3TBFvkt4hD5bstLddHl+sjcCC2uCR
WL+wKdhrmTgUKhUmhc4hivrnFLVRi1WKI0jHu3xk7qWQEO4ijSlfA2lZSW45MvJtyXPGqFZJd/ij
22MUa8rvsJlClVhyS0ah+6df03sODtQ0/o9VMQzO7dPSlMA8Sj4yS5Q07aiXeKTPCiwnl5XSNdj/
fqj6N/5lIY+N+0BOwPBAOF7N/iVnrJjDDwo4ByslL1at4YDz9eLEaYe3mPysV3j/bZj/OLEVFKeh
bZEOBNLtJd8SP+3B9CiNwYCC15r4wqg2PBowV7dZqYkdGWUUAO4Ck7SJrFsjOrlo+CEZ/M/DULMl
QQiO4jEN4Qa9agQw5Frc8HZkCp/ZeFkz+oxubgiD5HXVfacKuNtsIm89LMQl+DG4ZTO1JTlSxGRQ
2aEYnKWMDSzQxrCBIo3mH2ZgVim0HRkO2MKc8PyfyRuXL71Rraovmv0JbdUKyat7Xnq5ITBFbJnb
nu1oF9gIysbX+azTGzOHwJ57vlXzsYYNsOAJOEWY/d/ZaHAhNX7GuHa7kXQM9dCoHqjMILEzGYvF
LOEl5Csio85VS99n6iF+aLg7t/c0RKFN2QouwtsnoMRv4KA0uSAHlk2eyuUJLyNMDzC08TKeGn6c
xiB8CvXfK1h3xlup8GENE0J53i8DXQ5B6uqgD9XF1Xjvj2ZZFXib7PmSalMh7xI1uVeNXMWzlEAb
whTteyIiWix90fPYmVFXMcJt16OQFbIMfif+guT0yHVnGG5OXzEgUs5hEEzV+HfmnnHWW4UzmCMn
L/Uzt2WsOktCuqjJfo1Yk7wTY2j6eWPlsUMGbheb1dW2vO6OtPnKdk/5+/EoNcRVB1KRZev0mGDl
MBSFRvZcBUsATbMvaw8CqagUCb1H9HApjzFuPbJbY2nO3SMfzXrttdfRzxgRUG9wLMFIxUhFXKok
HsBFQ26YFkQJqYqjX2weJvG4fo0GT5YEvOcML0P5ynSgypknhHOd3VytO+W3/uqCk/8PWB49+80x
Aq1myrQRO56BS7oF2vr3TdKl40Ay/zwrspQE/E31YhuJ3V67frrIHJRNbFhYi4qT3V2UU9Iw7Ouq
s998ckhyMvY1/3aFQwe7qqttRM/SSSQsVEEbRx8tzVnRHfwnC3g9i3YxsWwRiJM3+v4VC0DkYQB/
VIpROgw40Kq4sFtEl5JmNOr3y2HF60qK9TZkTAbOjcFQ1dbu6EKwbEIPB0C7pKpygsr717TDFhVi
UWLq/i2EiE2KTIcXaFyrm8QWmkKg0KZQ8bcGC3i8/Y5TEdXGaK/0jy090yaHv5GO4bSCcHEyEvAJ
6K/rWt1p4A8c0C2XxazzPBHRUu38osatkDNOwy96KAH2Ug3O8dVllvtCvmHMtjBxIzDsb3piTFe5
UuKj2g8GS1rWgB2MqdQskpvAmOeKS8cz+DFqU/DoP/Twk/HKeoseruNU3uvwZ1qEFfBLywwq2ycH
xSOPv6pd57VBFIUjQcE8P6d6evlEsnnO9Of3qroJvvZDOYyFlderKD8YR5vkCosq6xaeJ0r/jg2s
0htrTLn7082iOQqo4fVQzcqx6VktkmXhYnOLa7wEqdDWKVvvZtpyNzfjtfYTpWUCZtbSVh6huKU9
U1jQ9my7zg9rpdUrEOIZF2eAB0GJb6m9AtjoNVEzG1cIXlyxZNMR8ASkfx5W20EcIVyOLfISk09s
4wtwwgUoV7MdMlLbbx0DZvhVbY+2Cx2GYgW/cbpOYVEp6UFqJtA47YJTfwFUs6VoLJyzK8xBBgiA
4ELbtbJVNwzn8asXcEB42mSgwnJ4J2rUlKsIc/QMYndBH8nZBu0ZpWICJhIylJb2sBhIbjnoAFXu
A7KFqtIjVUaoI5xb+VByvbNfNys4F0xxbzB18EVlfiEdyyQfbnMUXHA1f/Yb9Pg2KyOyDwQAf09Y
rPl2lhTpNlMI6YPrSgl8DuJC9IhDW9dz9U9RE5S2u6limVh76EJDE1fvqP9xZ+sys7wXExDkL5fW
bGW4M493e/JeiwbUxp2oYcQt+gs+5DY4i72uJ/7eq19H55hy6Q/I5fC99rFsgCu6duACxfKuWfs3
e9CmLNNqIWK3c/cLWaph4LDGnHUSl72+4vzoQ0zsqU98jlf7mSENX2axHuJqhfVLeUOhyEanq/n0
KjyG/IGVDcD9W0iZbXNy8GqDHOCUegZvuIRjDh1KQm/ZMNn4EZk6XVqhPsPt4b63hNUa/zKru5t7
EyU5qE1APwoEJDN/Xy0ngMAs9hvGXhWl8urcIpqewGAuQSM4DyEwSSramvaPVHG9WPWivVSIpbJ6
55XpRZ760r7BxhrN/J1QAGlSCA+s0I1nyUYRgVOfJooorLRxPBY2n1IkM40KWzQd5FpTnGmhquPh
AI3RexXMkDRaQxeZjkYPZwpuvzH2gcUxXy9GW03fg6TiQ/yH1l/PdSEH5GL5ICVykFy8UO5zdwBJ
eF4+ESIc+8WDt5qy6rT0uEvhZuGl94r3pnUgtbvTES2a4JL7Zxqn57IVNDDOHxAjmvJ9hY3KScQN
VVxlGwg62jH+0iLCya1qT94tsshbMyZb69DTLlt7vh/5hwUDwGCWrjmU4YHHkWbsVZdqa+JaD661
vGkuYMTCRd/Hs0Y6bSiq8tvrybgJ3D/TfN9qWO3UQBwtIwaOPuk3txTDvFzjV9+ht8MHJq/YHs25
IX1H1Dph9bFLx0NTH6ZjKhJO3YC0UVD+SzVFQEisRLn7ZAkDh7OH57t16XUOnjp4LS85CLI7adCZ
spBy7IbxAPcBBaJQTu3dmGGifgb1gMqMb+oKYSBJu8dzT+mrjoyOffxZzilKjGe+pYFMLSMXxGnB
NIGt7YwVvqDo1co2fTM0cgSMM5SWSYjyGJ6PjV2rXczpel1Un1KHwzie4DnY/VNTb3eF+0YUc54e
/JmGCBCBGvAm1L/vu9T6krIMIhzSn0Kp2V5wSOiO2lx2tGxBtPJ0kHjQheIs6lno0nmi+srXaaMV
zqYQ3SbqSyMcQNCHmcgtrDHuYwzBMd1GRlJHmX9gdCmMfwZkOL8qke8npXfuCtWP/NE+Q4zWBJnb
42TBgfV0ET0Nw4+iDqB8ohpnGDV8s9+V6aFZPrfJY8HIEssi19qqJKG0/Pd2Kcf9eCnk2BVg/iut
TXVZN5X/nmNfFqagRB/rzU4urpvFTT0WJnf4DDmw3d73Tq/EmGDcxmqz3K9JxerDf5XORTYXMQ8C
87d1r9d1jGIAmthyTpEIu8YQrijfjr+tov1KInvnNkIFIjx4yVmUMKOjiVSMcoKWq2eyt6tKJiJd
Xs8w7VCcKSp5YvTAb6lumxIEU7Bj6NUHukDI5q9rQvCSOyVdSTLda2aQLF+I3vEMy+YWWfR1Qp+Z
sb433zT+CBvDP6iz5iaJgYqPhnXvk90hGx1Nr11l35/NPwbLCCNSjqjU8k5MCdDkJIO4XMzdxm9m
zQJnY03RYTTIayZ+2ZtxKtthWoPOs0sZphVrzdBM2XTGvmxnm63ojQc729Fc9cf7rLBbxMr7mqiw
nchDnLYkPm58SGNLqEItwUpzhQy7Mls2IsdrXKTkULGT7d856XRgRQTeQGAq95JKRl6+E+5zQ///
Rhen0OO7dmnt036lsnIfn9XOt1rOqRfhrQCXiBupQaDn1RwUp8c8h4fouw4ocI7X3l++/3+h5JgS
ngHWt2cvlJu0h9PQeELZVv4ydf3925rTjZwTPxL2QdFHJEXrjznDgoI5k6fq0zbhiiOgLY51wOyg
F1r+U4LMByjS3j/rMZiJPiGUv9d2lRSakS7kHKSOE5QEPqA5uN50gIKv6KFsYLZCrT6x53W9A5OD
1W4Mp9tmSwZQDPX0e+Hty1OBrYxynRZnrc7rwxnZsHKoUpkRGyYmVBpus5IRav8cEhj396LA9pGH
B4NItv6iVvLeXSt+uab3DiEZGWLr5Yi+prORvQ8WyKXZGigiQZvoaNuOmS6cp42uA+aUxdXns2bT
xTCBe4xmOG2rwdQrYJGnN0b4ZfesKECPKnZyXksak5hlNS+2KwzTMWLzdE3/msy8O+no44f2nI13
wltjm7SQ4ET+qtjB6L7g1Nx0g9e5E+wXECz6WrXrVaXp31JAmRG7gl30ojqFPaj66sdah8aCPmAu
bRI/Za3WAlf2SFrmtIpF+LdspEsNzTOaTAjotmPQjfwhX4sJ6e1aU2xu7K/2MNN/O7jJUjS/1dvK
09GrmU1zSpJNJDxYJgi/99VbC2bTzS7QbxCguCkzzhrBAv2OYm+bF7ugG1amH7gMvfrOelk89JOO
Aeap/J/+MGqYGh6NA7cRMB3gPZVMv8TBq7dXn7dR4MmMVzPsufDGSp5hJbKNCjohPs4Y961xBbG7
gCbaLmQ3oG/7H++V+ppv+mNzI2EgF4wn7gJeA379rhBGLj6FnnUUw6ao9XJ6TT5jvLVnEqQ/vY8u
CgxTUO0DXem9wn5jKF/HSjlisGRwwB7xUvWefryiUsvEoLupAFebB1rePs5I9L+h4+k2kCD6WZ75
vrRl/joMzPi/DzXAHU/joIlfVYxVBFYsCNyakMiG16ojhLrSMVtd0uLLz2FLmr2lk9R/wxKw3AgG
sSJjh6xDF1fbOqYXSF/u0bhhMccx+gsBjcqAmGuN4YjlnoWc6kSVZ9h580c7D13JC2VL/iu9tahw
mk/0plRm5XV51vAQ1cwhT5ufn6GYBoZucVBhomXvrkNRkc/nKb7d1GSYHNyk3XYbXbtsjhDf/zzW
xB1k5zBgNpmh/rpxhV2PXW6m4Ve5SSBnOQTvPCX+BPA0FkHbUBRvHh/8cHE5xSzuX5fWdXcVhMAf
DQFeK37cuItBz39x5v/xrr9NVLk+1+HBQUpuk3x7pVfdbxt7fc/OMUFCjALRfeFV2LZOWHajraXT
GslZRkcv7Qvkytwl+E7VVTxMZ7vuueyxcozHJh9yshptxqse3HbVZK1oUyRqIkW9ZOuyCWxewSRR
vGU/M1ENxQSAiShRRWWa36ElUzKBkP4i16/fTKXXGLvv3lbecQy6ZXGD7HQFfquy2DQ/GuvV/IY1
w8+UG6nhFt2f8IP1KCnZMeXXKcU8XBVDg3aKusHaMtk6NC0M6GNPw17xU0/9VN8KvOqQiYeey4zg
DDQUq9vRIGdPpSOL2iwwkcZWHlbVlgQmBotSEYf4uxGssSnA0kbXqC3JJLmikT7Q3h5KnUDPdrD9
xpWEcNx7NjZSgZn7nuSdcEbr1QM7KpTWzemz8NYPo65Pq6AjBppqYbfsFpWYie9YOC/aBQL7BCqu
ZyVQ3NZVpU7E/w1aZomXCTk9MJ+SUhaSAyHFV4W8dBrnivfRVk3mekBMI+94JuXwGXGvtoQmH8ZN
32Lv0V5iRa+wIISM+QAoCZq4G+1xO6qDMX4dxi5TdtKmBTbM/FMd3hh6Vy9JktLSVQAVqq3xJsOf
COEmqdgNaqMaXxes6rdo2a79Dtjh9lqmdBwnsXbHeNrnDg/QgFqdCU/qh1o3Ok539llvODS/Rs+/
wYke/YDMvNohO5+osRCaBmlerPUq5wJ2DsZKoJtrnG6dxQBpVZh7o9uEYBMTJgPQk9tq+InbGnXO
PYELq6zEXdWUHekGsDTpHnw0AZYuRITXHJwnhUgTsrTNX6G86fvnb1YGs0PLEm46hg7POkcTXDoG
meFqe2Us84/L+x6mMii7bD8IyAOUH5RA85KmYdBqBw/a9hUSeGL75XQeQx6d06nzGX6Wmqqey2+e
u1wY4UZW0ZRjx68HPwT59SfeH8wmA+t4QiQeZQBPFi1v+lYQM7zxR8hatQzkEI34FAq8+wugihwI
ynNgHQsaa7Un9HZJ5NdTFV2P4Ue+lXOOdfPdmXA/FhcbJrv7lxLXxZlzrMzVsaCuIGVOSIQtSjQz
ZviZV4djH8YaE1iSz9awaAQuHN9jLZ00rXN+MwKaMVqt/e6EHqnqiGaPk+FkesD+HFPTlpMAMfqO
vYWWxFobvDOER32yyQgS256k2qUIo7hpNMGF98jYi9CkK86ksNrpC2gg0Hk793DETGmNudttxN8l
bxnc1cSSxFRrXwDLcqzIhQ1me6aGneAjurBs9QZoNiuc8PfzBJVMcqOqKkW9/CI2+Z2YQ+HxA7k+
zpd7qQOdcL6KWssvK+nTcg48uBVY4CPmPsloybJWaBjhgi/Yv8XMrhhBZ6br3DzbtjR79fMDpdgE
ZVqvnB96u5ihzixQK0MPBbT/TXFhmguWPHBvv/mhFxkxfp5sy2B+a2EnVSR/HhZ5HRTELK+tLHSs
9ISPV3jRiRuDi+NlsqrcDNbyqSP+5+y2n7vHUFrlFOCeYbE61TraN3u0YDNW0pvc3JC3kwN8DAFa
Dnw0wkbVrBOIcIwqzAzoX5M7hCV/6/OkWr4PAz53uNxlZJJo9G6V/to3860PrtlNo0qe99z4eOyy
Jvog3A3078J/8ZYNXStZMBoeCDCVVIKt4c88PXQG96MHovCfFBGlhs3bAn1jtOFy6sKERzezkAoC
eivswFX+OQj03TGx8BSWMjlYDoOm39pgLYKRMn9MSySeIoA8B4HEtJvV2aUw9UdWQ55WnFf5bYEu
b5+ZxKSWUvPQ8MTPSCrcmr2p7HFP3egbnaGM9RdY5ObGUVpldfj8xrFtohQEssjgZT2HD5EZYlM+
HIMETB8QFhOwnaKs5B/ELB0TiB9NWpfxCOPv9tmda2ySiABosNHtF3b++TNNT7mnbUZFnyItBK7Q
NSTKfb5XRW0BSfiwUsn2i+6d7OHHAQ2TVU5NUtRZ/5yAlrh48vcgpg+sR1Zz/TpcJDbNE+JvTsif
J28fo0VAatSHeJRXEUReRKB51nyD1x5oGfMl179OF+hXh2HtEaL5d3QzTigc4XdDXwoM6oQ5VJB4
P07zf0JqCFj8VE/EM7uXpNIQ+nZEHbZ8gnMXfPaAwJq652GxshXqyunFgYe2DarF5mnq53bByyNu
vxJ0v5BFj+ckXWO7IYeovSlf27eC8R7Xbe5AZVRiFUIq8HRpC2VZzjN9qvic/pcWBkAXEz8N3M0y
0/dr0rrN1U9wtzLMe+ynI0U0q+0rKOTIYyUGkWSIEHZDp2thWxKJXUPwgKQiNt78z1y2SUutvkGP
3lsZKbBx2mFzKDtJnotJENfEBfgOw5oHOuFR9hmNNayVCJdUAFAsogTQ66ElYFktiLNbfF5NE4Yk
GW9L7FH/bfgT9wShH5EdzdKVseuo6Tbpl9CbK3BkDClLBZrEiOuyLZArlsm1OEnW0UhQDhULhP3l
QWHHH+ZeoaPAVfQhVtxOtNewKD9jYTPcHwix7/ApRhvm7iM1ujhPYIsFNAVKnqz1nkvlcm0LVaMG
6sdsQHYD6ZNtD/U6bcVeU84iPSIE82V991VxOi20MlMcNFro6DADbQ0kq48REkIX6loxjw+TF2XF
zNWOQ2osCFmccYcgnQOhuzTWvLCjCX+pvbGNIoobglVQYxYMBgAaDqHO7q5QkbusnaV+AVW4hwxQ
jl0wgPA2elElPumbfZVo+ak/BMbn6WFGaFgNTrzhST5clhUzoYSddo2O0ukZ6NmwbjztQRxd8XTI
nyxm85HclHJ3Tmv9z11PnEze5FNyzjuX6qPFGSTIJEQXMCdHElb+eCUE5paGcimEs1yrsXn5DzWe
Jg8uStmaOzBlxunJ/zMi3naIXgJGnvW51P+fZOq1gfDYu90zJq3fnlBPpaT+btzIU42jqsFoCANz
AqwFen33mST+GfzMoP1iIahT7qkYEBz1Tv4QzqYScrAvQqJV9zvfWsURu8sUe1ZbNxTk6HqZXnJX
EoGxq+a08qT7u8yc93xonXwp+lPDSshkczrw3nONsQNihC3HuYKWZEeIbjm3NkUXkg/VTc15BFVK
zqfHInXM0cBk1TwLKtFiHJxmlhA2JsD3YJcp2v4uRF6jed1vZ4fM6bnpUROjHvCay8ZM6lBfl0No
Er1GCU+Q4a85qTNmfbMeaWg9PYmiNSmJ1ZeyldZht/EvEgu4qcl8kjTNWBgBzn2BwCHzVq8M/eCV
RtaG9e5D3xhJTWjdcZdCm8LidRfXeuBLe/gHLVaQMDdxQn4lrLhK3jzh/BqUlwzz8sdmo/SOdu2I
aUlXCUWLMpD0NgpFyK77uZ+OEQ27Sekf0wv81+KtccSZOmgf6cLDmXJ9HAJN+zm25xnS62dNPZQe
kUi88SByLQcjvUlbK14Asce7BJjaFk+dP2IsvfB5INe6ruTBLEBtJ9DHmHfegI1X4y05x1ohNpV7
xoAXaU3KK5zkwHbOxXklTucWMGPrlEqdm3A7uZu7w4hyygkj9X8nJtLBCywHOhn85PnSxBpI/Plw
W9dAjrX3RI+aNqDIZOCPvSRBdG6WMLZUmoustinOtPEkDGTWFdyKr96jvi+uDquZw/wTdUX91zEd
eAd71vrBSjzQcB9j9aN+9MGldMYCkGdf44biDgxxBynECllMIV2OObzRvBbrWUPYoxX2uMsJmKM8
EcbS55t6l9yKecTuhTQvL6PPxSpBNoCrNOrIsCRqZq3sxWrvSW8pH7iWM63WlQxbFmB8Hq7hwUec
bxacKOCKWj4P6Hs+3mtMX9SQK9AQ8ffWOpMTwEipPlADvfnqsBt/kEWH7vgIS8CRLfewE50XcqBx
PDxdV8zZVKhoSBVYtW8naODGo0gAF0Ex7cbhiH85V7lmGCsGt8PnxH/i8C8rJRBL2iFqU8BE5pNr
r9X3HkN6VuZMKG5ll5XFdmoMI02rakuPHfEbVSg8OWgFPit59rAXmhzeO2ktovT4joZ+CTZvXSME
GuyRaOXIMleapM5Bl+jV1kcwZCjjFWi7A/qbOrN7rzYdlWSH5d8zpuywXqHl+rQjQqNIats3ykj8
/T/TpHVlbPZoSfh4vauZ5pkmbX7HovX5Pkn4lRLWUkK0fG9hxHWj48dY6jYJ8qz3TMKG0oc/dyeS
CFcT729oYB4Zd8ohbcUadenlYBlzbF5IrACLt1zV6YD+ylcBt0XRBGW2041EyFauFoohPppUzwqe
bn09xAKCGux1QyYZQ+EYmj1z5FBZcRmglyNT60v4zFCwG9rTJE2C3TayzscHSzG3lrOzfQtahC8h
eQVlJaD2OkPg05LZkbkomQG5BviXWQskJqE0I1dlArcoGeT0OThdz9oC/U2k2tUcvhNFKUHMgIVA
7jeXz4bM5/1py4I0i8iVYUc8G9eAoXVPaBwmzf8p/iaEFTIMSF3CDh2mWcmMTpnFiNK4tkgB5d2N
9X9GAQZXCnCFt6oeg5uQOh6KHlISQ7Utpb+EMo2/mZYi6jy4ScnLqWy2KkQ4mYCXzu/mtnmNA6te
GFZGwA7ffuo5nVvCX3zNlmmn8WtsR4bJAXbUkl2YnWQw5M+3BiAT0SpsSFUWRCZJ+KCXpZBREYZx
bJ6HZ+KyIy/YZHLuLhQ+LL9XE9R5eFgvn0wEQ8fWX2UZmiSbzed3G7SsBbTooNgdWetXiUvqlvs/
+pwIY2Gq7uFJmZCasXMfu2cKnrLNNYsZUJSdLeuYXIg5HWB5bIr/3gkpgf3R/bDDZ2X8FQ/Y3CZN
k2GBKlq6BJSOk1qqQCorbeFiAAjkNO+K8l/h0Kvu+cMHRk61SNhN+GXkr5rSAufg5c10avm3y8Pm
EvjE3sGWLcvakY1GM3mw08v6+qTKDMMlfSPXNZ/V2hKUgqsCKiywYAPRtrbq+APSmiT9WkBfs+IK
Eegvj1Bx7hR86ebZ4GdxBCb7GUiEgXeihDtuVvy1ISt9/fNEW/SuAhORTXaVsL1/WSvu2FcAsSGO
/Ggr2L42SInJePKX7QNhuXsn9KrL/LFj6yhIu0rJnWHqRb8KdClZ8f/4Go8oSxTpsLckGQlaz5AD
8hv2f0aK0V+ScvtCktsZFLd/+8GbOCeF95GIXYmiGkoUxSmTZXMJAytaWu1wokFhFyC4o669b/1b
/v8wHnlVSNDkDbjupHh2AsaqjwZViLpC1WNGGO4XmVXh7YwZkhzqcX8BfqDx+Q+bBTYcwzfLMsoG
fmkSf6KHEsWbdr9qhrZoun/b0e6L705K1FbhYbVu7S94ScyYcDh0YZmOV498Sc3jdNrLS6aI1aJA
gMgKtZsJBUo4QX+IOvzmcudhdJtMN5ou3pXnVvEBif61lFTxdCrZiVgaHd0NF9oyc3Qqutj9cXm2
aoUHskNjjhCxei6NwABcrJamSi5v6vBOiIQcrrw48pxFGOpO0t1un/faSwKvHGMgyDcM541+9mJu
yAuerb13Z27BDt8zKy99O+M9HS8/6scA5rZyDGf1RxuUCu5QcGs9ih2SYgHPCUAQg+AHxMar01AU
NncPaeXrwVF+nGxnJllYQCxuPm2zHzY4ZXslXQZCGKqBiKRLql1QTSk3GZYBBQTB+70SJhFukwWb
RH+c0m0nHvKGDhLMkkc4snEzhdAT18XwLr0jdY4j9Q1T1cEwi8UfmoXysKJW5GQjdkvb5wh2leVN
sua4UMhlQ36+hUF3JJlEZL60S+r2MRLQfm2VslURG6ItuIn3W80h0I9ksyd4XvSWboRFa5qlFTwU
P2GR0ATFV9lU97uanAPbOaN2jPwOxxk6oWYx0CDxP8TFBmFsInDUh5fG4odPqixTWwxWjcYQHnxZ
DuCHsQpX5syFb451Zj2ZwR+2D+HDPRNOlkeczgJGoGQY85CSU4m0DEhiixf2AQFznL4KNwX8SJHA
w02dk0iifIEPZ3zq7tTCEvLYM2CRFkn5Qh7hpE0libVJkdCg5HYRJ6eNae4PSegC+4PXW1TQtfRe
wngbP/BNYCQn7cl8KQaRsZqrQoVjPupVdprp8RYje9X7ipjkWQXVS3vs1kflqquNdewTZYybCFtu
gzN/wMqjtGquaqMWsfMIu0Gwtu+t7eNNFfnbcHE0F5g5XmAz5SJ9lNYbOsT7DwId9sIv2AQpPGwV
1OP/Jfswc7wBR7lUsdsCgYSTtbpcNjMsATNBV5U6Evp4esDjDk8zcb1x8K69/9oi5Jtw9DH4RLYG
mGGLwYJFX/QVfU1kpHLWNsSVbWNV3BiNF22HOY1vyTBI2HCzdAKCGvzvJvst5Th2DBwoPxONqlk2
KgQSwn3+pmvouvCRsFwHcGItdEkni3m+3r+JxFnWOw8LtQEuE6YC/aTx6HEIoOqPpKQxq/3X4ayT
2WFW6Pt82XgGKTw7IHvnaL+++uS8nE66jXxiQiWs5oUIcbx/eLloh9SNoQE7uxw6fBhw9JrOCcKB
I6NfJ+gmqB2eb+DMAlEmtCAqRH1HrfYIT00of6z0MCD3zlgryMAv8Tj1ymlLPe+ZsBCbZJFMPUdT
UzySKWdkbUKEjTQiyAsjUZdZ0pKUah/qJYdpn2MV+4Olvgd0ltyAj+kJCd8QPJYKbH/NnMiCcnNy
YkgeWcmz9X6lIc++Jha/UGcvBwlX6P9PCdZuFZr6do3Wfc88VpjJ+dHLAFcAyNRQpL8nf6j1G0G2
E8rTbWRZYlFUaVQgsC3rjDu5UeVkSssRiUyrUFs1K428MIWjCctO0mzAHUpaeM/Wn3ZmNEqT5pAs
Kg5df4hd40VbgUdgbjKeLAoHogdXyiCMGNIWbIzKyW5R1ZcnICAyezyGxiqr7Zijy/ZUPhsbRwDX
grC91LoRwEo/hlz/YlRGfryA1EtMYEsxVizFfQFY7oc/8s3hFbO2x+LbsaN0qZ4bZ1NlvjVmAb9q
vmPy5ihZH8HYYvz2GsCzwVK/cx37ANzNWnAbRmF1+WR6ldrYyMjsdG5LUtSstweR7BRs8mw2EVDC
fL6srIepMqytsV8EhcnerXh8lp8BrgSekfYX6KhdbmFSp7ZMZIM3LnInsxpgYS9Gj2Btg1l8eYER
GNK/qyPf4S+xpvY5r+nmtihgKz1N7nBmACDrvGbgpiOmEl1Mc0kkGprh7wCfmrnszennbQvElaXO
ZYRqCbfpcKhavGhJz6uDnnDEvrd1SnErKoS2Wk/EZ73/RFgbIn9BG8Y2I8E7j8d184XJga4FMVdb
oYGLCL1Att/6EsdrCRMH0H0yhWU0MJhYTbkrilsMdZYH9D76onP1ZQkmhkQRO8zh78ngGDGujg65
1R3Q7B80T3qO0Tx4UBvaNHvDZdwNdX7pFcSJG0wYHs326abPZ0KR5635my360PjP4hXygbxjedY6
YFnYsSZQFq+brfLHOy1+rWw/AL3U1mtUpOlkhWIFHk53SS5AUhEQ8YX0HpOB7pUgGlRz+X2NClqL
q5hAzp7sBgGgfve7dbCdnrSzqWKXV/rBRFApHydY4vQ3+Tyq4gJH+bQiIdYPmp14p3adEkx9d1J1
PHKOP391tzAqTytTLTIZpCog3orxsOZZ6w4qkEqsrbwivM9ESaQfm/zkfEsMer7wKJvhRF4PLpfG
SMdVuG+1lwyWYggh6ODZWlgZC8ZWvcVjW06c+f/3q57nNZWXiq6Hc1rFT+t1ASb2R89ZD8lRBUX5
uCoQEuiOv6YH9A1PbUfSMM0ec00Ie4Dw+fVMD0N8eTG1l5bU1EbAYiHVv5LS2i51BI9IN+l/EXrB
/SbrjdCnK6HpO6w8cu3OyNHdEOsPsuhTfBhDqos4A1jvjpuDltAbyOspiDv6RLhK3x0zpdlufP4u
ENOt7UeFHNUwL9SZQTYl1m/d8xQFVA2Bmi1pXGrYOvTSbEQPvWYgp8nC4NCVR4+tmbp3FMrtUowS
s8C+tW2WNeOXrQsvdMM2sofT6Y6WRooOzRBODxYJ7ddFkkoqiAE9gU5bwNmHCIFMbIliGBEfJ/sL
ZJIvenjOS3ZOTSEBT2SXql3GwkFt/3JXLahraqX68AenI62e5lZsjGSlXYRa6vI1HlGSxZq4QYIh
KQ3v9CZJhE6nAFNuxoGkmTrfCOQ9U+tArCWdXXdWVwmwULWG+XSXlAvUwGYqL8pT4/lltI0CObL9
+lPhXO1ZQ80kQGE36j2e4UfkV7dSAzLEDu+oRg5uqDn8M4m9+GrZEqssbxEHEuFE/qQjCiX45PYl
FJ+z8iRVJfa8FhraBUuzRYILkgvms/vbRudqE0g1renVDGgU48jVHXeiZsfsEBzbTym4zLbVgRQx
JAi+5eTHFU9y2S/Qx3dbPvoenvj/2oZb/gt9BfP9dPJw3tJaTvNOALczu2FLyBbPNcowxzJoz+si
oFoCPINDFdiOX9PPdkBB+EvxJCLeuof405lhDZlb5ntHQGh9r1AcwlfpzCiXUGq7Kj48rr9jXxUY
LTml/MVODx/cF9LALOR0LNR6Jt9zRwLLhc1WO/q44H4U1wk1kUw96dCuP6u3VcXDHwOzSTJDVoJP
Sw57GTG0T7MlpfKsAVGAsPgbevQZyAUh/t4yXLBzn5OmFnidqUhyzcbrDIAHta9NG4YK1EoAM/B8
T8lHjtcvZkd6vrTgNYO8hkS3fms1gcGQMJG161+Uig8xoP1bIVArBcs3sNAaZZZOBCvwQ0EnKZJz
e3irY+khLP6/X2AS6+tniJeFt05/JiXJEVQzlSwoRMe6aYolt4asd045XFZGZHExnWQ2SNo0Fnzh
rCgS1HOx3Tq4TiDaiZpB/VGsc5snpMbinff/xdADD7Q6h8yDMK0wzDTsRI4T0o9/+PnApi0VvFcc
1SlBMMXBi8fBToVGOHuJGhPUcKS8BiWV+SqUNLatVNvEHt3Dwjgfjg72KV/pm5A2tszkd61pI3Kk
xONAgO6TdC6hNBwP6peVcw42wWgXVvJ/iMtejil3TSW3ywTHW20djBjEM81yFQsN6BizUPdATHWe
keBCAFbBsRXhH1aQlNAxas6ZDoJX+XeN5g8U3WIH00HLgaUekfrV+7V9nD43FUJPpftCXUX3rkb0
yF6+KQuQ6+wQR9nIVMuSNaENSP2g8vmWJ6U5MscXhBqXtdO+RS0JXCxty/yXbyUGSmPUyvhEkvTi
ZGGgytAuyjxFLhODgGPg94wRZgHCunCt5HB4XGeCzRbxMdRAhqwR9e1BMg1DpUJSqQbSFUrfj/4h
SBdyeobTQIIUxqNybv6uh1zYf02p/6i5DKkCwz6Ki2iV+CgtvQiJehRevAvWgHK3/1EKXQacPgHX
WzzkxbpSOLFBcnNC6Dbis86BorkIaYdo/QtOXIX4xoCBc4Nbm6r6zNT7sjCUmckcXEoh82ZleGSZ
2d+JZn6cqoRlvFJXpGZp4lnHYqTY8GJoWx3iWIu2HBiki9lT3CNPk/MNj8IFS+9ETXpkN9gSV14Y
oM2eDl45QPAEtD3zeeXxjVfAjxW6FplK5+YEMPv4Zivv9Kkr/Tx9TtWUShs5IWogBC5eUqcwK6dP
28SYcfwQOxSvVWmUVwROqtWsvoZqh9V6GJUsV0lJUrkRcViRobaRjdEk3pEGTe1xCbhciOpyZYSr
+Rvafga9ycY4pfEOUQuA73rPghcdJu8BXBk6SLK6HA3PTW2qIkpBiQw1StKfVdMWtdQwm7n105hc
08NZoYcgLLMWhBg1jQT6F1YuqiosbLZEfHyHSEEp2mAo4kAufB4UpNdVzOdEVLZagzZGmnRouDpS
lNa0PeIvIuiFL4994Y1aesJuKsN+ggvoPVQzBvaZFvt8JC2Td+m43UwfmZjYSMADs9VYKyAwpgMO
5CTFUnJheQ37kQVIpqP+GnQwh0IJc77lBmuxDhNu6PNPSen+u91gcTqXIzd7spimfvNlXq1Mud9w
XrWHD6MwRIdL/4tqhCMp+EXDNunBb9hKTC0VNC8wEKO6T7yijFFaV9wqVIJaGMWH7rExT6DuyzSB
XG3tvU5sI2lrEaOa70eVU1YBFXUY+uPkTClg4AQ8RAttpD3NjyTvCdu0E9aJXv7HVn9D0Y52Of1O
lAogQunGubj4PfgxhtyFEBSz9sROvE7v5FCDMe05FLf5c3RgSuUOfHjq9GhNxRW1EnwePgIuFNo/
OYQWvsrDC3VX+sqbTNWAkZQG2NrSAdiy10MSkmMAjSewhpk3dLe2LOnIXB18de6TJnL95vxGoinL
MZVtsyMyvwqWzCh+MaAINWRlN12l3CZKB0LBEX8VTx+9TXIzrUusdwOUvKHYGvS01rLL/MvtkQij
LVFUCv+THhShqwQxGtTFSMK3lQCgjDNouy0YpimjMABzo0/yj3MNbryt9jXERYjIaUVMSItj6I6B
ZnmBvdbh2sn9efUd3+2ltVqjSO4fKK+skipj/4w14RX3qRIPZ1794fc+XwtJfi7VG+QF5v7h02Wn
h1TFnO7t4RUYoGK6GkDZycAujVp9AiANDRT5pRLRuWmBRUEaft2KgpQENNynQKu0jbpipuhvG8iW
YWCb/u0z97DAOuGrdl4BXp4z10eQOH3tK+nP0BYOvQIF41/17SLHhYqW0gWwmOKV5oBosn9zIGZS
peJiAz/vsqLTipncdJtQMrqo5LyqJnu8XgMLQcu0RXsXUs/VdepuziFuxuAn7IWagUmuf1tt6TUa
QJyiuhcu4K4T+7R4g1EdSfqCJDhStkrGqbCUKIiGEfdATBzRbMspKXfU6vg/1MHB9pULfAj8x8HF
XlBJcSEfH5sQcP4uT8F+3Ou6Ib7e7FcipT03oZivqmg3XBqLOkwmhBAe9hkPK6Yu4GSKyJnYBOS/
/VJZZfqcPGOXjL8ITvGcPRHwVXapN2w01q5gouwH9up7Tf0QDAPRW3hp3bz+2DDAHxvuNGIYzs2T
T7VJ42LpUcolaJoJ93bhr4u+gMwz/+OcSHkDSjINFKfCQNj3Kw32G7JlJiAHdPRXqqVu+oprP7xs
aTA5HklS0WcuOOwz5ECxyGbLi3jlsWPQlvlNMkxbscpr7tTBxheUgjDNYqgE2lwY/2Ns/IDdyX4B
NgaEPRaS6NAIsih8MaIDUu4/Zd1Uuj4mmxLY+YM0nSRtV8CBMv44WoIFW+EKYBK/GNyDGQZ7+JgU
QCm6qpYg6YShEAyOL8oKBh31NUlcjp0QvnCqGLZI3FBY+8Ii0mnNj3WD6l1N1pZbL7q55TIf0qsy
Agl1Ilrk6Bb914UF6ftpaDC0ntqyZ+UhmgoGoc+KDpt8JikagdDiENydrPrGMRMPGTKZDOMXt9gp
WAye7ckZWR2jm6uDNiwrNHO1a972LLRXhtdKBaIJCC5qDp6BqHAmyCXDCyA0XRq8E8jCh2roHI52
GbSysUy5YVE9S9g7bRMyHjjK0Yml2W7Od7ozPsbsEiq02e8FSrD3wZ324+VEH7ug3i1zyT5pBmbM
Z6ef5nnL9XU89uaH2DGbOl5t1VN0VXHl1hEs5RGuDYOzHRF2HuzUOTEUcEJ1VKg1YphZ0tuJ4RAi
f1HkCg8qzjhywhK9jlXJ1dVy13iNa2CwaKD9mB0sBE6CIK+Uz5ow4XOE7bNehlVS5sP5UHz/M/g/
T6rIYRky/seRFQAiJUM/EBW6SfcAAry/KBUN3tGoScDc0bTmtB4ATx6xmDdDxkWIJ3FPMklvp1Y0
6EF6zcqCyArLDvuf29Dm0zrrVfOiWnGKCtgddw8rM12VLFgSg7Ytu+rsQ6IU+D0fBtYcSurqTlDS
E63zk9dejxIvlykx+giIyo7gGppBtNdWq8tG0BRZ32HGtheuZ5bMK13m1AJZJOBUzBzs/ZAzom59
KwP0rXdwc5ilXvdtEjGNOV2ZOY0unATXry0LwO0/zsCc92xR4YqfTJcj2exVCy50s1QsaHZQgvpo
77Gyn4v0pnIznm88iB30S0EcFbeSr4k1aF8g8RmH2xuKS7InsbnFJULlsPU50m9bEA3N2ClccL/1
xFx+BAzKkugdtEwRXICnOfSBD2yy7LUYUg6pSsmY4T50z5SBJsri4a/ApxkON9EqxpzxkMfJaoaH
62y80dMk6r9Pv11tk/OKbeXAOkIEcFBzli+Yyy+j2pSgGkCeW0O1kOWRJ/SBoXd9Hj/Qa70XmACu
cWIToOEZZtB98tiAbbnwl9gY454Lu/3DE2wqiFembrY8T8KzQhsMGNjL2bMPSWzf7RrmTgqStLoq
MwfUxyUokoapHHucukQSEOPhMTXsGEuQPoBRUdIx4FMuL0vbXYWl+gPMq1BGpM4z8XauZKoNeV3V
C8dm3Bp7EQKzDlmeXQsKlSdKO5hlV+d0vqf1LMan5XZoQ2szkZW3GzUX07Oachs27+bnkNHguHOn
/qLctMGfF1YGX+ugHQjC/7uUxY2tw7KuyONHueTZkoOT+SgbZrugSAPHWY9iSoUGBX5SZfGZ7JPr
EfgrgYp8nXGJ7CxvX+Pv6U3OgaGw+RZy5xPw73FV0eqZgM2tj/zNCUcoQC98iZxgdgZBXnESrXa8
VcTyHvzZ8MAiunPkIe2qUCY9OYbHQKRcVEtK8o48q/yRpnO5nT9ov5X7eaYjIxF3f1uoZhyumpX5
pfO+bWSof2azztoUNzqQ5ZhR6eqzVnXvXZy6Xi1gKLcUdsYIZfvYLvdOYBAYbm7uBRICFd6coFEf
qzBvGpsrj+tWIFDVKbcGL2eV0k6tg6TtJTNryLJCAZWzsxvcIzQxHHw+hhBUf6D/llsXFsfY+wl7
zVhA/1GhVNASaoSpykGfS4dJ7lI9T6aWEGSbb2oqd0LpFfjAzGREOefj0KBb7yKzVVK63oyChJna
niZ2gq/7HePMdRFYhOi0fxPYDYziC359+2s4odwj1xGwzGCFWxCAshdstiX93r7ZL8KDAVHMj7qb
HsMgPek3Rqmrz4U+KsenAvgcuoipFlHuKPnL5HZrR9QcPN8QqwmTxj+8M09jyjnKVTgwAHCftmaK
8JAN8O/MyTIARexFw2DuEwmE15dTSg+eC6/tSo3LCq0LzkyrhTg0ErdXB5KSVzA9qDtodisls4tA
bZx9V2u5byJ9Aa+ZwhTJk/jGWZ2JqKiuD6hEuKFtzry0GPx9AxzYqOQ4wcvX0PFEhBs+isKR0K8l
Zi9ynCHPbVWBm5nnt/whyY6CbLTavbWnPtygJXWtoV2L0lZnZ6Gn8OVsQBU1zkMJbPZUEkRAo0n+
SVJ1pkvZCh5MAvXvvydXV0WskjLPNVmOdADlXP8d3cg1z5WRQSIJ7ooRngzYPNNWD7ZvIxfCyAjJ
i/y8kUrbn5JfIc0J+nWcTFl48HPZfpqRUeaKR5NrFy8NC0n4UOdglO7Rq7am4VN54yug5/023PVW
bfdd/B8wkPElZc8jZqJba6voHyC5/kIIPq8tw3qxruNkJS9P+n5kZJot7aQP5YRFnlaoPmW0xKCJ
WdogmH3Way0fPxdi3xmCj1mXcW/izp6jzETATVp2y08+c2peTz4fiosn+xFDARixYUXtgMxbZgJM
XI7d3IuGF6qEAsMPEvXpUrWj8RPnajq8N+D3D2r/HcebtzOU1C2QRumdilmKv/X8iLrrjlJhtp/5
0H6y8Vz+qKL0KDcYjpl1cE2r0fB5gx6yiXgV3iltaYsi87a27x7tc4BER9i9nH/Z9JuBsMjW5l2U
DbnIbVHv4HI36EPI4guvqyM8cOUj/wwCUB1qRE2PEFyMGgNd43CCijpuG0qfqcQlI9iuY0KHFyVE
3EKPxVEyFew8rcVh5gCe2WtQPYHHbtsTdcRIWbc1srM6sWaQ/E7s5wTR2XURkFWSjnFECjcGfCjv
XdqMM41qO7Gd/e/eXyhuNk1ESMObGUaubxsBnUEXxV0ASj444aaROCCIhLKiHnWeZL/jbkbj7Dfn
V7V1aEEzY0pKHR358ZgyxnQMQM8ZgcNLCurGnHoOSDbR8z1uOICI48vR97y797glRDKGv6CCvdHV
vAwYQpZ19wTA3rueoju7+h8vB0Th7BqB38Jr6PuDVREkRvYS1fQYRWppgfxbRxnE9IjV+x0++rXQ
fqal3ctEJgbK3Sgdjzeyv8TKjHttkuvmKQMwWcLNu0SOC7H2hvuxGAM7ru75fxG7l6i4zlj1a3yv
1TWnYJwR0Y9r7z9GLclgtfWOKQ83q7gaJpsdNzeSMHhIm8HxIxFBTDOessqWZ0ojuPOKCZgKBBbg
ZU0QtvIHdPtjlKGzC52dkO4Oj8JVQQDCCaue34MCmCIfdBA0lZ2D8teuGLcJOY0gBi+RXZXdyBpt
IO2Xt7ra1IAO4qixUvw5kbsT0LnRPQwABKWaKaYziiVJ2ywz1VwPFzqEkHHR3DxEoFillyJ/9y35
/4hH8evTW2MrIExEWYYnAHTwLxpol1o6yM84P2vKEQzvhaLu2KBok0zFsckBXvyPsKM8uIBhRRj+
twqCoD0koGcuG1LRMsO25RFUJtaYCdq/JvbhgGlvQOY+AEpbsBkMQho+mtqtIIFA1/9GQnq8Dupp
FBQVrADFX2CWTXVUdTUubAy0JL7I3iXE/rnNG1bYTuYEC9XOwsiFzeS/LW3nW+Y11OdE4FcJH7Zm
7M9n/qkxDgJ94FHECELMCKcXq1SE3rxFHM2ovO1Kzr6/r9V+3a2P6GbPJdhmTgIhSUSExysf0VY9
nfgbeMR3i1noQL1TPBp2YuicDS42JwAnxqzEL8qLjEZ4lFJ8Hjtf85ADGkBO6Eajk2AKEvzvrC35
koBMyQzJtjdVf1l2M0rjGCil2zP22UJt8fVIxnM7+4s+lJ47l7k0jqe8Dbb9Mnx1mS9iGNzIBRnx
u/1mbGfKXVKWssk3kXQagDdqbHoO+SBA6X3wGE+NA/9XBILDPWNrGJwcDFaT0VfJoM/Hy5cJ5bPw
U57E2bsEu6Modj5phVW0WU5QKouthRKoIUVmoelQwqsxksSD62S9IHI28MAghsNSSMzSnbym4Zkx
YeDwk/xNvU9xZVWo45P3WbFnMsso0FgtqMxFy+ibWz4U+jQmMjPVsAXu/8PNwAqypstGe8tRGn9+
xxDrNfAjoIhoUs2Jtn6y4weCpFSBK6e/hYnV+xhpi6e0zk9xj+cJw5orNACYSVHs2S5gBN6fVYV4
M/oF7CIjB+F6TxpPDcffiZ2YA6cx+grUkqckkvQ7aK4Y8obmmyf6xsAF4MlwFigyw9GjvkmGCGsQ
0PdfPgzO0lmVlRdxMHch1SgWolpe8h1IA9ZOgD7XUHQo0+aQDIdvU+ZZoHW86VT3u7uLAbVMH4JT
H6KwFVQOyKjV/EKgF3QPe8+BNFa/Pp1syNYXDL1HupfHrptVom+eIrw5frBCNHXJoFMLIneQLRSy
9Bu+sgh7MEv5IYnvOC+DOh29dXNm62J/ykLgSZ7ATR0pMftin0EgBCmrZ0jLgR2OsacNWfiuokHV
9ZA8EgipmDImvBdRIVH2RaOW8oJNm5nBUZGFLdF9/hrImP185/obaJMkm7DFD3fUo5XOeBWB710Y
venR+8goUd+0PKa/JzyMPMfjYV+oWPAKtbP/3ONh1IRuhyAw8gWWfsgO1s9XlF51+PxvKVYUQXLF
QIAcc9Jy3vQwRAl79kv1ez2mBojgmZ3iIM8c+zBB+Ww3+RzwjjDJEvDASP7JEq0ZRs/qz6nJ5Fw1
tnKzl7y+pIGobeYS4TeRUnLrW8oJjGgF1qykXe7/186iLTXBsINu2wpSsRzOQV2QThAEFQdiJ5tF
EKHiTFPUS+PbwBiNce5PUvQ1rojlQ1UOVifcQtim9fSa/PAEMHQIb5IPDsXkybQsF29CegFhqKHt
vryQgNG4+1zbem9RZZzX9x+io7fF8gnFhMU6ZekpTEuRKUBVWzmORAJeQh4OjJirjYZ/CLGy1KZy
vOTLw1habBwXAaUAAQc2rcV2wBcIakYiO3eIaQBy7BmntkHMhPknlRDHl0oUH8rIGj6ecTdStDx6
sgyXqVb5rLCuzYv22bNA84RY4RHR2pB79gGblSOsbX17wRcbi1kuVmyYITWNd7hcMx3mF4cPf3yU
nGtMz0rbH8JqIowdoh8uLV7x8mF04rsqTX5BOY04PRW66aL4Ce86Xdb+Of+xbVCy9ke4s9ni5nZx
rBZAoCgtz3WaHwc32g5FJBzjDktu3AJYIXDgDpXjq+6/28Uuh6Qgsh6pwS/bgz9RJohqZQLQL1ux
YSAdJBHmLrzIkbe1YG2zft3rcZ8jJWQXBt68KHAFjCg1ooyP5gJmGtTJnZLhwZ59tMYK/GO91Zdv
X1EwcKSMQ13HRQvE+rVYod7hGayTEj92oHoWx60hQAC7mpsmGrE+Xv4y+4kZZy6Ow5fhodR82j62
3sS+pY1RZ6qBhKAm0Jg7/zwclSppnX/SlhB5vb99m/9hdNR84iybePA/glf+J2cPKPbM77Yna2Gi
2+aMzp4NfdqlyXM56iLPG2SCpGjACes9Gv574n1KmdRPdH9TD0FZNS5ReQ7waHlPJ/brJGtIVtPP
n+QzdCeIais28vBnURWUCIjq+IMEkY5+vwSod1TPG46sR60Rk8+eyZ35slfdYukjkuVcZvQuidmd
Dnn6kzZ+9w09a6hVieUxM5exJx4UX0BPqXufvw5rT5aHkW9iKLeL+Oac5/HHF8Rj7WvgfEJwjKg5
iP4dYB46rZqhOtKQcmC+BDLqGcL7M87NuWQTwpN0HuLdB4OeTZ4yrglRwawWlrxM1frAgsaDzVLt
ySzW2PQI7BbpvOV8QUci6l4lpPXy7R7X0lDCXgBbgn4uA3r46a9i1d2EsEhYp5VE+ZkyLlfSqtZj
MI5sB/m7wnuGhJMGImhH2nkONoPjDN16d5QdpigB8TJRV55/lINo/0w9rhTrVAsFa1uophSuIzg2
bB4e5kLoNbC8S8GHJwFEPXoeabEQ2CB70/CyHSxVZHnWSq+wkubFeWyIm074Wlmg/+oEnlb/BGz7
QA6u17SNzZ5+m81frSjEHCUMNZGh2gOwrRFp/ZSmatAS5ZTIvMqA62zGV6yTF2vzl42GTJJqljzI
Idu2OzwvmW0u83S04XSp1ikbHTh9G3C+3uCHvndj2ZUNNgbqabHacnHQcP2feKHS6R0CSEpJhnGF
MUkEWckOV5JfYuL6AX2PeRZ9KDM/rnQxgw8T9wXbtQkpyWSa/6XaD25t2+iVoIQZyRy8CrcsslPQ
r1IXrrC/iR6JUGbOn/ZW/xHJB+Sca+Iss3U5iaEcDJ5xFcDv98fXadcIg6SPmW+7rToxD1ib2hgv
bdV4LgjPekMxAbS7PtViMMLrbZRxJ91j3o2pEIuh7sojzRibs/Sf4rLCIDA1YAnezR2grG5wJVKK
OeI7ab6C8tMKS15OwiKC6nB3FKL7BphohZnTENN9n1zjakRD+evVxnEa5wdSAHM7QTL2WraOAJMF
+UGOT0+k4sUOupRjoH8jWsYZZS5t4fASptLEksHoX1Ql7E6lCx94V3Mw/I8+O+z5liyHKkSBurmh
PEJeXTA+7eGWwNReVYzvoiF2YgKwmo3pm3F3+/I4m1ztic8RdpXV65TaOaQkt4YOFbOgV/41k0zc
xhP7OPjFFge6o9vvPifM4+2Qf9PkyNHLH2Rc1lYISt6QqAO3E5y9ABA4dmi2DbWNhkPvC1nGQYpq
p+Q0EmEFz6QQ1XezqnVgs5LpHkNAWPFQGwAdBle7RFsdWJMTFXrzMn7doCk58FKmh511AguwFC6s
Fu/Z6dxER7jdKOoh9Fb1GT8fwmu31+gMRHbruvbyyG7aZssEIvK9yGkYqWKAMWPP65EpJ9RkJvoN
GrClWQllY+s6BLAUrWeePJAn+FWxgpZJ53j3OKgaE+qJT8GLdMVRL730wrYZ5YZgti/YZwRPDSLq
HlMMJNibzHYRvKXN3YnjveqNxOpHhuk8OSBq73iT0crh5T2SBYzH1NDy1ZcI57rYZlOuOX0ZZQxF
Toq34yuFmoV4BgQ4f8GrUIfUZQ5VVEu7D08GihcCi8x7nAxCaUfl93OdPGvL4DiCKF0dwBEEYGZF
RauvUI1suCcKEYUgYrRYukC96ScB6w0lTlbwM+rAaNyjI/l4ilPLBySrWDUM/iMvyuWD3kr1bSNz
kltLeLc+grC+8OKjpTSgFhYvU4pCr5mbRiER0jZT/gxT1/paz4t4WEPHm6pw63sOS4MKnt3gfYTt
UQA9YSmpVY+BGgkgQ3WiCppTc9yjXel/t7XB8GRup3Szphi7bi4UBN63q3ut6lVXeTkGTglbKyif
hsUDxak4TYdREM3HWoDzY68gKAdS2cUi8WYeBlOlvAKcs5Wk1M5bvAXxDBR4RSjxwyrmBaMWeYct
tIoMSrUwYXqvU7bBgPmuXDM+wyBxGdk6K1yGoNNyYZT4TwnvOx+01L8VsNKnO0C2Jeo/KjRfI4sW
TWaZC7a2XgieEed8Jw8HRv/f3s16UETV6xWq50/qSZf61JkCZY406ayKJ8L84VPA5Y8NY7gfoH2O
YMnoLIJTQLrXE/Cer5FjaEqVf4YiesSyFSciobd7lfair7+2qpMFBa2WdF4pFBrLrh+e0r7MCiGu
hT8r3452LNfTmGSSFH1RChrYxhqf4VybjB1RZ5o31TdiSe5Y1ftWEc3KnO6Lq3fH3q7bJT8sto3I
U3lirPQn7oYsDn/DsNUCUEampvd5KQy6+4nu+P8ivJg/G0bI99Ebk0vgX+aAoj61QpoJa8Onm6qK
/kOEP3A7Pktqc7pVvkrCOYqYHrihl35pZXvYUCrM5B96WodqvjQzk/0jpeZYqiYkuu3GObvcMFdU
umNyaHD8V+AfnUt5OUdYOvqwMhoWjzXLIOdG/oI0T/dkefZKozP53sS9Lood7bD6ZxMDSrtbkMmg
QlABQ1wsoXGDh62XmbqdfNXLKSwCo/gUWGXO5mFVW2akoF3srLrqnfbAmdiOJIKQU67nWSH2UKXs
e3FJG7eqOtSvqMJW3JXfv5INYjWZQ8NGELehxjQBkBIE22srOUNT3qf/Nbw8qiz7EMjEieaL6Dvy
aXe5So2tkkGuwJ+MU/pxuBMtN4gtQ1Fn97i0KC013RwbO7cZCpZK5EVpeNP050I4YlfofiSYHoS0
gA89ySwbMCtTq6YWegepZ/YgsKej3qkqshTY8GGfOW9h7LZB05J/lOIxbf4O81fWWeQc2JNs553T
sbbDC7m7HnVGlHG9l2NA8O5GSS/2VtV08Dw5jid58xw4+R5Dy0LFD7YyLLekcs2H9CmX6nPPUhu3
gazy+br78qptKBVL2S6w+OvDLAHtA+OH92JyagKNkQOhpUl8IfkMeSwP2JiFXgkleV07wJeDE72D
9V5yJmoAbzhKVlQcvwUHPMr6XbwkaCI9tBbjXU39I+/qnhts832BBqXZWj2JA86jmJKShEC3aE9N
6glzaSLsFbxpeklIeklIJWk8RZR9yeId9TlT4VPOgPLakWmxHtzr8wJB97iG513m7YEUyecGZyP9
YXwmNyQIvDKBuNbCFIEWuVvUSveWgcGBNVlca1chAigHWo8K+nGUiA4zcHXWa6SUQOpoX0FmSmFJ
hcJuuQpDT1YUCEBFOL8izo4XHGiCQkBxVrWzEbPtq5ezPrPVj/lY55Ym56aQYj5aFQ4xaRVCov3f
Sw6C0XYAkql6rnx75FRPDQu3JNQ2RK0FptqpcDtP//4eZ0ZDTmqiBCjz5NOVlJfDBmniIEB09LxK
rnLceb1BVJPug9pjUTaFII66q+k13SW/SqLVQ4cUG+EA5t0NlJisxSyAnertOn6SDmKsO84m6XfJ
X62TcQV985JaPyuChUdGXE7vgTTZXxacFntp6Iqo+kwaypVxz4mbprH30NFVBXqyP7xsxZbyBWye
o0eMJ6Es4z/WoJkUida+QxlSYw9yGbBZqO4XMeLK3AztMYeN+xMe4GFDwfnv0iEA4IpFqcSqyaqY
JFpablfxCIUPlXGM7USdaMfZtkquWSBie0ZBGVMOhqviRABZCLzBelU1MZMxlbHPVHHRPN1HnXts
oZIEw6XBvA35bHkxVZUN8Ix47YbI7kY7jASsdGMOYB7P8y1an5wPtYdZr4T2KvRMSfJ8v574UI5T
MRgfOfJ4fqUqQoVgrtz6YdRZuxoBHU1NbKY1WW1ahVU3gK0pe55kt+gaxVBF/GE0lEIZdQWpqYcF
HIQDYK1fT5YxdrY/nlHb3x+Qbf/6FZmLlCfVJlzyQLgztJnQYZrK9OoheSXZnf+fLiyNvnSVlPGJ
ay7FTUzL+41zG19+IUbgPdIIx3FY/Ow+WRYQKTXmyCwOVo4UyIRPB+0ppZlPTci2Ja5fbvZNKAmZ
wAqiS8/shoD0JbQzk1szqo/2oOUiJ4M9s0EMjQbp/41yUE+ja5FvIHWzZ3uL/KCCyzQiToFYg0L1
8t7KlhWpWm/RvusDQpc3tVekFUd3YFtfkIkxF+MECofE2LgU3cYwn59xeyp3BtYKpczipoMJ7sL0
ePLPcGYW7jdk+mtTYKzSSPhjkUCAPidgbw5uKyV7bkKrAWlpXXq21BVgHMpd0JJspIyLgBQ+wJBh
spJCMIlnM6bjvz3h6I/OKI5hSiOzzjxQy7vRoECyINptivU5Pd4IPRZfMDgWB6b7c0sa3O3BiOeM
6OtYYl9yuf3SipNcY83eUuy4GaGa1CXCqs/+ugEDcAbvyzstl76PGOLAl6pnO0fbyKgYxxaBwkLg
paB9QU55oVfshkm1b8dq4zMgV8R+bPICb/kfxl/FNYAQgGaUXHhMG4bT7LNlQQrrKgQAOW0gMlAy
llVZEsom2MvSXUSgnZFEQxdswG6Q0GY8aPl18oVYI0BL719t1prle4Y40xBbbYHSncAELSYXLRtp
rznkTRBdQ55Epe+E+F+eGs5zB70rvnwQlyz2C9CJTuYzpwev+xLpwrHcPhTz7wgdeDfEzvMs6dTF
62EmO2NfGZzRgENx5+MXakMdmd7YkKxB6ZGfp6pD0BfGA1HrtSO7QqjU2K3KukwbVgAkGClDT59W
vhMdNZQEqAnLi5t4M84DHG0LpOtxmyY8m36No+HWPdATh0gozDWSod8HWPUeMaomoYH3XkiSbidj
ygPc7yjq4g3eqSlTHeURT9kJwX1sWXFZGHqJBssyHvUDazWKnOs0JfuR6/uGzqbpHKiO9CK3pniq
qozg+2Cz6LaGXSjyIDxauoYHLVEN85Rf1BZ6NCWN0QqZOnKCIB86XsdLhM3NyihsAlehU5JeCL22
svE5Kli/FmBiIOPs7qbsO4NjjVSPTVNuAuZkBF+hy2eGbsvAjs9DY/OXchc/NaPCXIbJfYHjZVHx
zHqoZDctwgqVJsWV3/N7vjhLO2tcIu8z6Eue5x7+ztZ/HnRAIYI2BNVIN4M35BpOjV1vDS9dqNkh
oxf6yJS2GTLTTvmSRSnUGgTbYXqiMgbj9pqXLEeXr+1N0WL2SUG8nOtzvbRbotkDwwPbHqCxZMhB
ffrBGmBkaGasCkX15II5ifw0pK9BRbNjzjkatfWUOtisKBlDy1rRQdL/AkbfBNHJXT0SoEKBS+d3
iQG861ZlyRbx9UHS3b4sFINokJ1/R7QMOsS5mR18v9wpb+j0+0a7NOLE0/G2RexkygG64IaWUvWc
Io20nvPQSVQRhKnNaSVU52as8jo5gd1t5jzG9a9Afs812CfOuK/PBtdnukTxPGI8m0166mOC4tU1
EdRODFMaxDGgTPjhIJcVdhIaVz5rIGKWsguYvpPkIgbpmvXZPykBqH5bpLQwF5bL+V2J7Mun8IE9
l/6qsoFMHYcw9z2qcyfessAA0UhUkJJm92z9pYr0azXt0qRsARIzyBwnb6nnL8wWDlTOrSGIgr37
sC6LAfrUB8SoFdo4KnYuuyXfkMwUI1Ag3k6RD0OvGe5TgUPll3X8rXo/ybY7s7o8AQZ/dmpYT7F1
VHb0At/TJ5jWjmCTPPgRFFB6JmIUs37r2KWFjiAH7HspGR76sPxDgB7yhVuMKxybdjTWfSo+jJ+X
H3kZPz7B3RXNJ9f1JSnUevyeqXnvbBjsgPZmmrXIgIztTb135V4Mza68y2OnOWzMl+uiEpVOdbAr
3QeKWIL27qbCHGae1Rw75zJV2r/Rxv4INF6J3vpYAJlSkbA/PnyztvYUi9D9KH2BLhjPS0gi+zRE
22iFDaHuTWQb6IKiqITJzRYFUeDvs9mg0Qq/nso7F+Lrq6qMbGYU77sZcFHOSimdBYOIKMC+mFmX
4AllR3FPcLTpz8r/S32C5BWhlB52ix6SlJAv1zD5xx44RIBdsdy2o78Yt6o+cvFfXH3EW0PG9n5n
Mm09c1sAmjV/dH8VTtRn2C8gcpz+l+IKQkSuTmLkCuAOwjUWmP/cp1c7EB4UABGDy5DxljJqY3ZQ
V9iOaIvR4DwQxU9qUvlU4KNVJQF4mwH78cffkSTpeMCLMb+uvmUncAOzPyZMD8Nkn2JVz7V6Pg3f
rYX31D9TWmcJO8DCeSmvIzabdVQIxNLaV7/uuhlIkT8jvYYAzLvvow/+5uoGIBftdQg42bABfWUK
WBuoDgUrL3T7lMl+4C0JqNjWR6dev2+UTwcrV64fgJ/cgUK826xfj5NSWmqQnCMkV+U7ItfbRl28
OPTuyfKehH26pnAKX7OECgJNVLDylscebBxysNPT7qcjB3jIhmiu0Qw87Uzja9Tgl9TzJGYwA2qL
bTmXpbx9bX5S4ZLmbAhRwiC6FcZJXzyw3tUvtplNyuf7Xb+9lVEPlpj8U01SRUDGSgYictlzEjZ7
VQoOTHjuGZ/i5IeReAXO9dHnlKJRJ98fstoBahdFYXeHXoaHYy0P7DNybgVPkYKnrXD6yeHdBgjF
mza3eKlX+Zr8pfE2MRkw94rpbyGp1DGnSrTtsp1CoVcbs8ovpTv3xUW00zNzlNT6ijLGz9/ZSVc2
LJCByiQ0zdqpz8cForFCU55M55GggSfoKkBdyC5SHA7Kv9dvwQEvI72c0D5174Wgq3TL+nQlrt20
dpSoi0Bj3unnQUVFmy3X+euEt0fZgi4xtXyRK5uQBxa83q9mLzxFb5IalJ6mKq2mbWENh78JqDIK
pmWeA/g4bBuxcDDZQvBDc9xXZWSSvn3bn6t8TaD0o5zbgDtRjUv3RswwAKvU1pIHWXi97h1jEuUC
7pUXhkOUzjsve1xiII72vyRBALWK7dJVW9c9u3Xf2STXDr0oWbFhrWee+hyCaq79AA45e1J5xR7g
sJL6InlMffCHTJWV0xVGf23ZjncRJJlL4vDgiLmlB/zQwHGzOwq+/hHI8kLtE07bYFN9P+C3SfA2
CYHgbb7xPXmNa8lg1aCiQ6TANvZq6W7X2IKmTGn17V/1kVsQI2ovdVunRrCeyALTfZD/ikWRwjtz
COzcWSCZ/l3cPYng7jtfjmIHKVfCn7e1O51MvC72uOCbDUHwaGO5Mj2yG4B0kIR55WNXOBSKMMlO
j+hvZK7+SJTvn4eKjBq3+7y2e4FOVoKhn+YD81ER06aOMO7To/Afd0PfFIB2F3+o3MBWj11AebA8
qMSOPvY1QI1NV96dYvb+v3HqPWTKNxcQ80pNSDbBMPI0KeDRFp8YklLQvzYPqeUATo4tcVx5Sodj
u3IDtSPwcWHpOFVH+FZ7+Kg9IqkyoptzU/BbGJvK7r5m9cWMNS098cy+LS1bM3M/gUmCXjoSXJ4+
N4sdHY3Z4CCpN93jY03qWK2DPvTeDr13eYFrfvlxyjrO9tZNDNg3K8z660Oq4cqeOYE3s2CjzFPX
KB2q00Qwnox3y8R/8TZIp3QzuhYmLLjs4QTM+j6zX5TfmiulrQMHEy2tnj69metv2wAumIM1Y3/r
0uv11BuTiB8dbA7bjk1GT6NcfmB/PuvCDDRKvEDrWQR+F9W7wUFWCAVkvvnqfLXVJqx5s+L9lr5f
SvqAH8sZceEUUfauuNGZ9NDIO7tQ2XnGJb7urCpXO94Islkv2M6pG0rlsEG36XTo4nne3w1aBbHh
v79O5M75WZvGh1wXzDxAi3G6eVizKJcCN2V6I3V0yHqCVfdkO8PraQ32phHn8Td8cG1CJXwVwwOU
ZB/OiFaUUSEVb0H7U5VajkJTApKy3A1U5l0G2Bp0gspD/9NTEc9r+5fXF8+GZfpkKrrqXaYrDNcQ
EUKaZw+W214D4USx019YtnrDHY3jkZFniQYkKHVmcbJjNRkkOtZzjNnW2HpWsjLA3dOPFpeM4JdP
DjrRJV3fhmkoTVxPrdvOiJcLWunZnFIsvk8WyvmAFPVPQWqkVmedHYP+jMs93q0L1RlJCTpGv6Ka
wpcrXtm15AWTGBzfn8r+3/wDQyliHW/ZzmgRZc5V+r1jeE5PMx/R18s7176zZQkZYd4yB2L/BJfB
4dx0BOgLPHM6OI3yIvW+d4mUk0uJkbRfowyPpTRBd2gQfTtWD1M4hvUhHrxImqkyrwX/x4lytYvS
vA1T8VJGcabiz9Z4dVJd3AVtgIkAJgifk633MYmQR9KJxpSCyOr7wzonDXa3fwblimvdHAIU6RAB
b9+wpXoUnqyXNhLyACgt2tZamlyn1dRqZB4uv+gW/TcFi6qC52nSV2+qycHBR8wRQquEMspn4qi+
eLQJU5fhFZCa1DDmuTwlMM8N7cBudMqJ9Nm0imnAXyOlOsTH/68FUcIn6KwaPles7R+aYwpC4zv1
ShdofogXCN5/kA9KuEsb3KNT0vuXtJOmHzoZgwcmWPTRIe0Pv11N+V9/bYKiTAEzeS8M6DUqq7gv
OVHuu/GKIJKdY3OPVJefW3fKACaS0GJVs3yoD7agZi2kYd/88WYFCUnQWgSB7k5ScrC+kMC7y3So
53k44cjOJYSg0Lq9DakdjiK5iTc2VVfxVLWIMCwI9nH/ZgpRvp9KSdsXVh9WcYx4W2TMtoKxTBXk
yiylLeSsCTqIPIlByAShRRilHcTCHPrj3zLOai1IzMad/bzMLf0mV7mhdenhvGthD/0mFZhbgobt
MwktkiUY/983LN5ANAGfu9uqy9sX0xmswYBrTinEgd+5pXSeEJkwyXKfK6AhlUWpEepoWqTivTZ9
Z/8jPYz93yfdcm7W39StI3qrJHjqZx1emA6Mzit+/C3UziRIP8X433G5fmZUGeuV3MrTP9khcdUd
+2T21yNiTO+Wn0FIiDWXCCt40VOkskCRTRLQYcisu81hCy0z1OqIXg0CIHgfu8c42lT6hSu2qOAc
wA5Zru1np+EXPRak2dgpC+yF0J7GinG8Uaz4v2A1pcKAQqH1ZyWKM/FrurwHiag1RqsDM9spvkRW
ZcKb0GdWSrn4RFICGboxvqKDdULBZ/upf8w+1HPN48tNVUVHD987oHmRi3syCgHCX0VaOwb3QYM6
LJsXH68UnCtLju9ibvOmbzJHBI5NGAbe0hiBX8XFVL6b+g4nMKrJxobqafiidybT6yk4cvPoLL5m
U0WoA79iEoQywAhW0AODXI0sARsu7JPka/1tvCIQsXz5W3rWQH3IKNeX2b114jyBYFls0Q1jDj7c
QUTHmm/mD/0B6nUdA7v1iWeA3mXiAdlWkzCoJH5tiYh15shq7XK/XVr/tAm4iUor+TveZw2Z491V
DpwWkK29Fl9j7DWRzcBKG69V7lfTf1f297ShJLdBuRIiG5rN3S1k1nbPJJkQEMFVoDVI+Klpu7jN
/Pr55xYtMAEvlcc0/PYwb1G0Wm/KPC16CfZniFgH9ijpLoNVfpQr0J7sv8bjSeACVbp2ovG9csDE
prMgeGTU+smKQ35SY7UL6pW6JuwD5/yTypQ6tjQkLXRwomVCkLgX9wz/GtKfji06chHgbgiKnqpL
8HCbVRzobFoV82s4yoErvg9vJcVfrkU/8oMt6yOY1Hf2RnvY3iJ0dwryz2DLakHByyJs2P++B8Zn
1T4o80X7M72W/KHUhmj3KJymmYGHsSsQV02pcWRaKgCPb2GdNB9n9LO73/MCrSuZhxCTXX2oUmg0
fk+tOwxrA9Fj4tA3BkGg2NPlyHTdnSAPV/phVqEuaPvbZxHyw6SsUg2NEFEw/npAgTAYunXLyk1s
POPWtJF1HbFFk/9zQFn38y6WP3G9zR6ihwnkZ7Jl4eLNoUP6BF3zt0dBvwmNcRg4Z6z17u/SVs+k
kCtXIRZyWIjic0pklcBT5VY3iD0gcBvyYhU3cjAKlvOr4BbCwF81MxVvO0vA4WBLaLPAcWBna9aj
2Cbid/DC/C3Kbf8doVZyLvqJThphZ+xscxGhcRXcK7XDjqo0pRfH2yHRr+6d+Oz3hbFOoX/t0+CU
2IgZIMGA0wPRrFrJZQEVZBEA/gTMISdoxrZQfodylc33+Ztyd6bCaA7ZMV7a1MN2JwZZR5N2y2LR
gtU8gCX/inVsOVERzdwo52LrtNoQNex7m1RjbWH3VgjZDc6myuTgY2PsYUipov4GSljHAVggU9Qu
8mN7vbv0RwClSvMTKNXv72wWjslXivkVJMAB2IWUPXvNGmhqXhQj4/H8ZXnkOiG6rQnHkxtAApSi
TBw3lc091TAPH61wwQARHoks9RwTnq/CdwqFceGKWGmX2PGdaBBgvkMCS4p5wEiI09Kn+X7/+x4q
Cdzx6b+9HVPdrMXiTtJFib5PvBdmoxt0i4dq9Iyj6qtV4BMuLD9yetsGS16rwSmC8xBqZ+Jh4AZe
j7WjrzeJ7voGVdbkAiMJIINvWBkVT/W9/e4D//bsRFKKrHkIIfhrgfb1hmSwqrszHmVcn9oMggOR
CpCNtmEXO5sD4kF/KrcFxBw8fqeTnEizceh/PExNMSKdDb309jBrzXLiLBOyixuasub/koByXagG
2DcxitCKwQ2usaCXzt/Cb93GXg6VQf7uwuYComnt3V4eATHmvZ8jg7keKToZ4W8NIPqhgiltEPwR
RgQg5cXIEMFmEXlEajX3sukNlz6AQgc+BKPm//GrrfiV/XAiDTz+/Wk9rgIxZGZEN78FL69cWS3I
YwJA1wvVrixqaEFpgy2yW+BDBtBXCWbJiBGHigFrNkCD0LZBYyKiteL4TOpQejHInFOn9Y5OtZ6d
YVFvNQsGdRGw1PkjRID5yHetQjq0Y+KknYi7nJW2Eok+yGUKhsfG/A3IOdRp63sB1GxTAS+NMrkA
unOj9z7HJB5FdQXW6NMG0Myx20MVTRoEMxgXG6/kr+QQCaRcoJiTX0uVijUoCTH4rq/HJ2raQJb/
RKhVacg25meQ7vAfXwTNbU9YCxiCcP1tSzZbq0SyHwZTTi7zkx3ElAXk1xKQuT9SaXheVpvUTSfD
7evQHzvRvX7O5zuh2jZVnhpkhgsFWhQB8HAGgG+z2o8vQLB+0QzXkk2V8SuKQiz10PV8y9e4wjEz
2QJP5g6M1+8Vr3jCOJEP+Mk0H9FTycyOTAald8f6HjNA/LijKiW2aCREHptOcf4r8U8MMznNpJW/
Bt0YiBlhc8Sj/3zML/s3VfkkpVwHjx1N7SmzpySHWjtTAJeKk7PVPkqfGrOpGRZxIDR2RiMmw17e
HhS6v1YDJe/20M+H0U5wDCVux3fZKLwZWhKarXItl5ktt4QuCFYzXhEpTWdZu+uoo6LeLb6EFc+W
UzJ2ZN/4AnVFAKESDAlrURyl3gXOXEn9rmSIh7lEjeehQ6BJvmu0YZjQP2bBZzp1HbR8fcrQFVCP
Oyz9qwlsXmPHDTKm7e1OG5JZN3G34jox7IsGY/f2J8p6wBbOrwGW0F4wEbLdUqG3dS8ekmx2Q3B3
aEgYSi+Emu9I13LDpUV26pcf/VQgn3TNrnCvDBqY0/uM2T/5eEdHztqA86YleFaVeJWKlzOQlibr
HRYOSrjFYGann15igA0LU4QZf6LMQQfMd95TQeDB6W84V0BLf58gT5DBQMzx/WX1ZWRX0ftQwDBr
o10UP8KcioYxgAUpnB0zBeNzYhlWQ+dDpp8N8c/04Y6dA831JOmvZqAOwAXqdaVMqShHi/xDn5B1
NyoHzUXhllgpI29dtL6LPUXOXlYNkLpnPd7ENY7imhhvpBm+j0Cxy65cktm5IlP4lm/RB/1cOFxU
/LwOQ68SkcxkI92bu1Fsb4l72HoImdCfx75+jltB6obPfyd3ZA5IcDr1wPvtsCpRudVnqnRn0dBQ
W9Bo3nKSf8Q1vJ4XLC+Du9d9lWmMaWEzFWfOvPXDggS0DFWRHQFBJfnJbYq1uNy0KEjuxBks/SwW
q68hzQ60h2QFUnNRAGDU8C/gAkswV4v1WXoM6/UuyZu4+uVhmUm2UAR8/2luA7twgHcbaC6a/CBF
H2WQaM36Emdjr5Yto93Sl9+uau7iLrzyh0rNCZ+KyWL/762fud+5UH779E+59qVswfU5kzEoJa7t
QgdnxzRVSdtDJppYraw2XU4P6+jsCnShCobPQELgROj7ZiP2nqYbFfYBoKZrKeyAAV52VHrz78ce
5SBrJkNjQOkcOE8DfaWFsjEXHjBhVuKK0xqEzdRpHXW7rRW0i3yEqwFLPpsBMHckrYt0nzKGjoYC
UGttITDxl7F0Q+aC6ytv8/b8rfbbuLkQj+MG3KYSDqvkBd4fX+vBTmoKTd3LyDWNnKi55CtFpC4X
pquP/ekdQTxEgzv2aDnXA+ZH4yiRRXpqPnO8I3pqbKghl5W5xutQpsqZTyRvSo85G3vdQZvMYVpd
ouDI/xJg8Nnb1rNmZg3wwOnpjf/hh66CPZzD751jikEjJJQlN9bNMNZgq44AWSbgqxhPtIvG7ld/
5rgq4IgFzYk5KclIxIYk+RypWaKPTWK+ZkrogZo2FMjIpgwTZtlojpLByptdzfT13vyi9p/tFa84
CA0DP6Zjye1O4bSCaNfyY1O2blaT7EZzEWtCIPIGfs5hFsPzmmw6i8QlUudSFDZYgx5GOeF9Do7V
6hs94cdeiRGawSyGO64Agm7TqA3ST5f2eovE2LDYXyA8kBm3Uec8cp1ZJz4pIPcd9BraG62zvPC1
HQ4+CeCUQhZvgsh8OfaAtRoYLss96nqN+QCMxc6IazTHnm8Osz+Thjd2tPycRfmMObLrDwUGfujR
v4nYGH+upkOXw2I+4grjlnvwneloKxftfFhR2X/sEWlYGNcpYeBazAGUAp+kM8sb3TNeQl3uMlEl
uthzssmqwfttzQGJvg8QjqKSm766Dl0e6aTHKBaq7K/FnlqLIxh6HTC2/Chi7sME3/s2aOVFTyBo
nEZOseo/ecuQFypaNG4C2SXbpcvP4sYKl3OXXDIaNVH+iYDCV4nhvY7exqNf20pcABy/5e4UVb/m
VgzGi5qjJIxfGUDCkRItF0cHRawvamsHKIl5B6n/CMJ5AIJNf0pdwBADnRM5g/FlMSj+T4C9gfu6
YSqpM4urS07mBAPGyZNgrtH3+zgFOfRSFKGEpotKjc7lwzhRjvsXa1DSJfNaKl8t4eIKLr+ULxUO
ez88K1dHv0CVX/EP/WOg94nBv8NEDxeQZwnTRBejxU/fKiDijcHTWP1SijSzd+kRz6HvQsTuynHp
fSBowDhbgK2VKA+wliOTU/Mm31ztm9EuGEpBYCFAt9oTw+G3z8to5a9JiHJpX+dKekRjQY8qVKcw
lOTTiMTY0ryxFcWDyu7NkRiwzXEPiodcxwpI1k/eJUZyA4CW9VesA/oZhlGDC9go+YdEUYesPoAI
kzmrDlP9sYfvNqsGiDdraFpCzux9A16xjcTMCoeiCdEZtvA7SfMq4DCoD458LXDfo04ZFFEmaAPj
G6+gJknOgWiMM2rm1VTufgH27dNmgDgkZAKsUkklwKTlqjIz2IT2/jVNsFQeNo/vAqndQ3A0xwr1
U4vckICex2eKjC6PJTKVQYbnsf8HMwoSv5lJ4fLX468jCXT+hYdqDvFKuP7rqEI3dRgSjBUHUIuJ
RgZDQRtmQpG0DWO6bHUawzN6SHvSiD3keFkJdDZvjchaG4FgiiciWq3hjcwd+tMi/aIGDgToukKK
EmCzHTk5zVARQzKII3foAu8BWc8PL6MOu43TE7GM9/gI96H64mVehPDrShJkdiWGfiVdvoeGMxq2
XvNlbachWXAC5W70CkBLAC+KgB4Fv1dcO+73Eu/ZiIi1gr9ojZSdxcdm9QwQg7xwk6BSpgycBVnQ
i8lFeQYJw6xdrZkg2q8E92UGpl6PHN8jj9PRtIOnuC1+FwCUcrh4hoeOq84nx7URFLPWgg759FbW
okCpNhCnYCjn+mFaCU99gNBjwNUtmsCuPkJTM84qHSjH+Tb3m6zepLLSZrLqN2JHNg5hCT5pxqUR
ljc8pTotQEwbErfCtoBS2mnDunMMfArsmvXDOpPZe8EXwvxGiPr5BWTiYlsPPzArKaQGyiw8xT3G
q/F+9cg6Dkzbjvhi6adRgFIuYST2CbK2mYoZ9YCT4R+c2D8+5QwfPxH7GWaLp3GghYA6aORgS3Dx
mjsIxa5Z40eWJ3taKcwhVNTn3S2SaunViAS0fR4RsaGuy5K/2QUSEgtmtKliI2Jwk81Wifu+LsFg
uAOZEoXCX+/dL9yeSUwiaY7aVTwayTf1JxSR6lFLITI4YwFuV2GcUNYxsd0SaI1EAGcO/yz6m44Y
vD4nfoCbvh3i7G6hczRQYUp8cuDQ+POOPMVJIVk7oyLvj09tjWsiTtCWOOzc07fJ5tgal/CqYE62
LTt6zRWUhO1LrwVbz2ZQoond1+6WhFy+bU0V2FkOPuL23bqFYKYMqxcdOrGVZ4HYHFhJUmL55Hqx
eLzITEG9Mfi1mSezVBjnUGcI9mTc8sBl9cs/buESBkb7JrL6OBgaASOAa2X2Ey3Cg/FxelPmOHX/
mlriCfnxnaZBOdXlCGGZleL2IZavaN0+9nXjLk0UmIvemWqRwANYXYhaF6Jn4qWgSHjqRm/SbXWp
8FuC7WypUdDEd4Qaw71ddUYmlPKzhx2nCh0okbSYSsy3sjhQ8795qF8XOBZ+VrYBI9YHH5wrHrSz
Qd4j1PX9RWkd0EJFxryIPHWsG5tTc2xo0ln3OZZp4GrzRzyd02ku8NNox9E30O5JsogsybQYMbql
o3ogTz8/zlVG0zqF/XWVeA9RmAhIddr23svwVExjsYL4BGhIoD0//j40SsvKhZYhN4sclMpMTc6Y
g/iWTD29bMzrF0OhchYulTIf0odGX9QF+/1ju8hCTvXS/jW04u8YIItklT0TxKgl7AV5oqOQnAY4
UAEwjqZeohQZ/bv+iRJa1yWWC73YnjpAWoEtIa9+GExZVMgurkW7MO0MFKzs3yrbAxAn0sveF/Xi
r9ASSlAYkv1IijiNfJJq0pPgWFmp5Qk5DiAoWZZRDuIG8WfpvQ/Wcg93IrgGdCrrSzVSfgfUmJ6m
N9dX9RP0ln594oa1ag3IHQvBONXxB426tNHtW7vzbSbptX/duQPswToCS1p/eeJnY6gnqprqbNi1
Hte3mUDPxCvj5Nhg5NUXNMLOjZSQ6PMctmnGk6zLXBfSSvq0Ki9RU9Fk5MYp5p/I6UtTtGpCE0Di
yKUyBM9dSNPQCA/1w5krgQt9x5De6fap8Cy8bgtQXRg/O5uSmejXuuB8yAja+3CWSdZp799t233s
AAhYQ72oAFIE7+xRlAopYMQA9chGMMqIhrvDglqAerZLWKGYhHu2vI9TbaM7KYNBSA9GtygQUk0B
2hkkpefj4UxXPf6i/tWpUgxpthWPJvQr8IZYcCG25zJ4nSf5hFJvOGI9V50OkRVFjd8FYO4IqCcv
iIW95D7W12JO1NvoqSMFhCf/6PGfERZqV22JWBRGvLbvzzIj3oY9Y1pxyg3gXLWk9A4uTupBq4yM
S+wnhbm9WYoXm8ZEePMjWgXTnpKi36+cfnEWH4yWKmem5h6Q95DPS9NHJkUKAWL/bgfYjbqJV35B
IdRNyuQFm0F5pWtG3xrxoqN9LPWH1keg4FQl/v42ENVJcgU41ejWE95yGrAc4Nu2hLZu4nRyzqO+
2Y7kq6iR38o3kvqXZVR65ecC5G/0mL9OeQBfhB6WTI+EmpYTHVxmUqxveOxO5eVwhYcoScXHWhOv
IKIh7YUDp5VQ4Rwlb6F79Q1uhNj1d+n3ixIA+wuxbzOvIUV6c9xtAmBVJzQYhGx2bS4mN9WykBHk
drhbp7jBzQ7vxa3LpK+GzugzTfJrAAwLnEmomTLtdHUMJZi+1TVNYJezujItQbYw2ALxb6S6LDl4
fbF4M/zxkr8EpwFBtJKPWlVUSlM2ohzvqf6qDAifds/SSEfTWMwmtA7FGNPxmHlvqNS6Oe67GGm1
Clcti9itzuAALY8Cwmk6Ma4/QLO7I67dT1dbNAK9vk9ObEUIRTsVi2GFPyv1iqwm1Xpg9bC9B0Eo
/GiAqEyfsJp9IVALxs3wmSC6uKLtHCh37eIAltun4fh1LqnnizWY6xgSYJbCD00Efl7jVZvqrmmd
MpNpzJ/pifhXgayMAKP1YPrE9OX/8Wz0RFmoBK+0RSp0EbNmNmVZADtKSuWY2U/MbswMQPDTtRtW
DftMJWyqd6prNTgSCqF6+qnLS6dpMQMnOha2HBW8aGTr8uA6Mr9mP5vqsHGK+lJiylqpe+heQ1BH
5mN29+OQpxR02YTPBBozvqUDO8dKEa9ojyN7JDJHysNTG1lscPp/PeYGOIuefyMO0bO7UuWm6uIR
G6ouawNJV5caRfniPR6Dgu0RhMqGdwMBxCMdbhdIBKqTT07FeYevGQ0Y00ZAVfAmqfitSdROS/fc
ifWwkSWNYhOaEycAAgKs+sdI7trnm0yvS9G1/MoP8aRMDbg9iFl9BFdi6JZ2OqUg/Hc/KpeeZxHD
tZVHsyzIOqvABY5NOnFTZEU5sExITYqqvKZXk6GcZCg631B+tcnsgaoos4U+caN2kR0MVKx2fybx
GcUOtA+fvURib98u3GmPECFQBaH65bKWYpsqSZhJ4J42HR6SHxdQRNBstyko8CSBOemxTKL9AX8e
q1nZHrKhs9unzrV5Bl0WX3jfj7wMihu7NmYeH9KMfEGqcWn80JNS1ngSXtgh6hEy/Y/fXlaSEghN
j/k6Nc/GqXi93sSnX8a93lXuxM9e9TNiAFHiBwoZ5hvhJUIIUGH4uNgfatnDETwAZOfxguXdXeVT
nq0QaH4jkHpFYv6YiBi5AemBB5wUJZLvhNJzW7/0ZwhU5nJ2enAo0zX8Ur61FTwuQ/RYCpM9BKEz
eka+DIJ5r2sKcJrHX7ei1z9dDnaMXxlN/o7gANFF86QakjiK18BAn8iTA3XUOv3RC3w0V4R3rxi5
ct3fSVnt3cug5Q0w5+I0oK95X11IH7uGYsMi81a4tYE4S3IYAZmWZ41uRUowkYX1U/+B7mh2MMdt
L42UdQofghzLUyCzb0QfI8HjdWdbCebCKaRl82j0b+SXz1nMMyLeuHeWCR889KW9b14hzQf0M5pC
JgErBMSlqelvE7rGS2refhOaprNHHwPad0fpiZtW3SrzQwViN5mRq13sV1906T+gcPpF9p4C/sgV
t+OYOTZYdjbn0kKs56WXEVInsPjq/+UJ1sdCj0GPvxh1RPXS1XwWheGsmw0tuh6yEWPnthsiPr8H
TeaUTF/0/GhoxXaoLKQEQAPd7fLDtQIRu+1upOO+zhuXUl77gld58IbdZR+BAe4xIjPo50+cFeBz
wA9ktCHM6eEHqJkwDsgGB9yzHKR4wRvpxtSq5VJOwcS0N6P4KSc+Kx6FA/z/vJCeoK4uH4N5279x
wTnQpvE3vRGlWVzEbXL0KWFbMd6ZTSRz2/yYa6FOnVvRx38E+G0jXff/kZpA/pqXMn5LikbBjq4E
i+EHGEcTpLWXHEHQQ5VeG2lHbGkYg8XjZlYR9viOgsjx0Awx9Enu1tEjKfvECBmACLT2iBIaJr79
A6Qck949ejPNTxSNws2mVTFN/jpBu4aI5hKA4p9Ti8ez3dtYGYZZ7NAmhnPtmE41sLG8eYv2F7j4
YWG9szknGStD+5KnJ1XOA1TgLa64xWqp31pe73YmVKsDYWRCMQJZa5YS30EWxXDoAIDoy7eqG+Jq
fw+lPW2pHRobR/rj87ZDhsq2be2yLI3mRT+nPdVpKTTn0TKfRVZ4WmzW59wQhTHkEIVImp2EMaa6
RGMYDrRzH0r4CyhgLqWYPYni491PbiCnd+6CIvqPIJVddYomdkbeakUfHUoGGGiBH5sOzZ9Pgwip
p79LuwGUk+/Xi4oEcFa/FYes8WfZTjDMa9Vx/bEA/8oP+FYiRsTUH4EpaN9S55nnM/Pfp3yc3E5j
MGFOGCUejflNNzHvAZ02s6Y+sHjX++64Xw2O8F/PwXmghQ7F6S16nvZuUjQ9pnsxT7B7TNDXQEYf
RBHAHa8wrS4Q0b2kRrq4TXRxqykoMrD35RTcH1HKW6UhjvJ2bknTWvs6ZpygiI/P5IU9XDLxY62n
JHZFhVMr6rqWcOG4qzK6q26pncjrbrDA5LbUaLHD8r0VymBOpKUPjGiMM8bsjEzQyVIhDiomRu67
UOMohtrtYEP6DVGmoD2XuJSBurG+z2lhg2gpNvTX6qfH/XSmyZLwJ6CzEpLv8H/l45D3LIlG1CWA
PLjoXpl5zKh0rkNGdhbccaXbWVGYcWXC+M/C3ppLD5Cq0jxfcda6Fahy1hoWIDpUGxC4kjCweEf7
0LCpKpTIR9AxDnan2+lrIu2kkDKs9N7LQYeZijQsKy4E9neGA6HrYkS2Zy3eORoljgqJWwCOGUgT
LW4+mPlh8fRCY0D8U9XIbS/BWEV6LM2oePl8CUNy5WoPyKLV/1LJidpU8Vi9jBzBTd7DeiR2neO2
JUFWwQnnuA+cOxo2QG92U4g4z9iswFL++59kFP7VnnCbQ/Am/G6Xo0Xj9frflI8gHcOV8Da9hHxn
1wJxinbuM0rIMNg7OLxhgUJI4VdJuRnuC0MTRsdLoN1/FPuxhxgMz33MvPTwXIl6iZLF2/bYrSSW
N3CTQBouVXEzs0SK2ganPbOQJx7TlNRmHMDzNpesyPnNARK2JM2BN1LYRhcdhaa3u3ZC9ThKDr0w
aetYs8l7Mx12nvvsE6ES3hI0h7dytpXtwzXumGQTxkdSUEi3BF+5+UNAeIFxllh3HHWKflY6jStr
hyC+TUdF1M8t3NMv4Lqy6ydj0ZbG/Px7IN/a+L9WfHuVsU60fnDFG+NIf/XKS0swjdzmFXgYvY8F
IrQlliE7LqVrdQeObIcETNHvCfHF05X5f9M3TS+H5RLMQOsI9AGyccbym5rL6QED6vEmRHwo0cg4
jy7ckhbfsLKRPuyE7UJbTfMI/Rp7Y3s98yv4n0w2vXDDyabW6Tdqwa2LP/stUm4uMWHLgJLSNGka
wznA1/1pCGj1r1qN8GNsN7MaG4TG0/Zirstc9zGh8mxJQznfd5GQhgKOPSIj3EDEPwmxnYMk7m1Z
p5dcMMNVH6sgdb9LSOiBx7cxi001a371heGHmaXK5Hfmk1B13aRCRFgYcMcqafShuyvf/8gSmp4U
jJSI9+AwubOPZQtN9yRnbM6n5L/m+iAk23d6BNifUHMDQe+HsVVmCbRieP5LLLwKJvCm3OVEdXGF
BpVNacs3ztgO/fpWcdBLI4XDN2JhI2agJXSkWTF2WKLaQXWfbNZSb6qe0k4H7ERASeo10oAzTWzG
WOp5lnzNP88YChSez9FAL8idpYiNxNBG5sLTjXpfGPU92J76RIeiy/eUb659r0rGSqWN3EWbVos8
XdcruaNoOgPWlU6avJ6O0hfMBqjWVH65PdArZm0/IwoZdoxwRH1gGpr+OkN+26dDZh5/1nbPSFRx
1qVndBagn+Yhixh6611tzibXYNowbyeGfjgnlFbYCpo+mn1lK+sOVJbJ6BxEYrLDdfw+5WkqoFHw
JTzbf6UXi4q/Bw87pIA4N9z4vnDKNq3BT207yAlUnQU7JF+xnlia7YB1qSei9yQ5QsPp4JcT6zRZ
qmfpiwU+eSNmL3LYYgKX+vitoS1HqwITsPGMqeieh/2DVXmBJY0PcoH+q9cKHl59vMAOwlPZh98/
jeBG9QAFsFT6cTeSxAWURrApnE+tBBGyBS+z1X3ZfCS3iCN/X9b8j7DU3EiOIKJbL7S+jZXC/XlI
/B/8x5YQ721u8+jj9P4uoqMgSFUxHqjGRVSK9zjjnODhm1vPF7yesTM4bemk7Xo7FxnWPLvtWfsg
MeW5/TlsU+CPiziDPzjgQ9kb6oTulmpoM9UiHXE9W8uY0NTRpwAZW/VboI0UoJF6ocdtOvCe0TWY
UvMvJ6m7rF0WK4MNi/sgolzmyyOapq/LfmEtAYCiOu1fXIpmbsAU5QCLtASAuW+mlQhQHlveEV+W
MtmPIMR3nCa+pSoqXDRqpgcOEcjhZ3QpSD5xDybWsMo/gF5lhNfoYq0HI7vRpyt23crur3hjjowA
9rD20qJi7jxdmhms5uPcjAgIgJTu2hJDjvkmkqKXlZS9f/1oZjgd9uFEGr4Gd+1k10ELMn6vtZO2
3jUlI0pUdhmyN93R5MZxfr9t9yz6jskuJklQHyCxA5an2X2DFr7OhMQDBMZ0GpgM4e4IaEhWKCay
frD6a4+uRzjFsQtWQAdvgW1KL56LZTj4inv0DP91RsMg9wNHXHwLB6QzD6YUa9iK1zVG1ImsfHLE
WEr8MwXuC3AA/QFjFXp535MbgFvXL8Nolbl6PASsb9SRuKfOcp1FHC36k/no+MNnq2yNLDBgEQJm
G+oxurdT82wycVFVKX7uVZ2F88lB+DAvTpjfEpJBQZED7WDtAlsrCO25cwD3toIawyO/sph6gVTB
5863P6+OMRVyFzJJ1lBZKH9m9p072NQcYoGjbKObR2z2CxZGQnt0xXw88lRhjpyfOK9Cga/XPeeb
CUJd7zyna6IVwOMKWP5Ruzm/RTVVD45fya4/BBROA2yP6ee5b6Dm383QiY7tuxmzFTMGiI4kin99
eZ7Z7UEt0W9zkdzL9voxWQw7rGh+WBYiTOE49gVczZKDeHO8OaYC6ieEKXGIT1iMkE7gnzs+Ok9s
SziJvntMk8XOTAxi9MWwoarhYGuXzoMDt7fmMHfj4EC8Jc852twNk7W+mPqlobYWrAm3egmyDWgu
NS/Odu0yVYZkuc38IxqHKXt7RSj8Ndnep6LT4ImMoWylQSl8pfOH5H1WwDSI0/mQHgRISmnVi7CT
etu/GbxiCRYL71u+Af6HHwMzrqy8dn49dec5kfpBEY9vo81rol6w99h96xXXpnqm6luocleCZ9ob
gC/5lhMev76PAWVKhB5gjhEECmH1IpCPOSUku4YyefRfCUEtq9ISYiLpwJkscR9bQrKK1PnDK+5H
BOrbnrwLFWcMSWXPkH49WtL9VJavxQDN2/c74JdPmHcJnsHCVw7OXSu1D21P8bRlOo8AkefApCvN
nL/l7FtnUsgyHfB1Wn+aOGnNJJp3SeRg3u++8lvqNXmp/csB2BysNMUEuN+pnMu84VtwiuaruYSO
quP3s9Iqe6mwmRvHYh/O25shGVJVaq7+yyQpnYSfhGzWoynYUcy3MYgcu3nWY/y8nhSihq+krz+0
VV2RLSN7+41QCiD0HA1jKPwx0p/Vwj+cZmioFRIYC7z9zIzoB9FD1foZwXlHpP843JxnNGyws5RQ
weaqMc0YY5u4UpSVLyW4TqKGkmJx/msyeCtUIvZ8fIRqzG8w+7oL40sMq0s8m/gP81P18uQPPvLh
9JBQNt75Eo2RzKPa89S4VLdZFTWA69dcY7Lkw9GpOaOaH5HM7Aze3FS7d8S013ymSOsFc/ABoow4
FY9cu3IrX0DLFWgrTIH36TgIhrkfDNT08b/zDAr1Hetts76+3HGSC1JClsi2yfnhlGFRfFzTmltO
IzWPLX5kKo3eWsXoEUWO3/5JO9Ugu+ZfQyQfB8zDVj4ajo8yxSX+jdTQAtDWpWCCvbwHV0vaVcqX
tKYXuWFdPUVwbt+7JMHuBURz0p+UaD4Q5kT7fUb7G12ko+iysl3lqBlQwCTVUcLjgOqiAlk+GA7a
/PNGTJA80OnW5R9ZysI0nzKSIE4fpQj3vltOVcasiGI9fyd0cGhKvz2SIMiF52ajKBWIF1NckywS
tNsBVsxRgODStE48rxpesqAXYDdQCeOhImMM+nY6SQ6hzZE2q4Z/+aewn47jWUuLZEzpyn7ix1uq
v5rjw3ZcaC+ubDvFxgUivenkkZLWETLiVDUuFXJeknkjt0cR83VO9IL31BLM6RdNfFRP/V6Dbwaw
iYLCtKbzHi0zGhx+f0GmVhoYn1Vq72JKzz9gWmOSp9o7fnptJMZEX1ny31bq/h+CEXhjEP+ufpjH
Azo+P/t7+q4/73aJYpCiNIGWF8TkSImQzJO6m5mxDZ4v8exJmxCXdpa37k1iqYD1qNc06FIkxACR
lM1GWY6NZa8y2ltlFN6bZ7Uzpiw99tiSdiYiToQs+mOcYY8p1j/o1CVCSpoMs5jQAvl4Z2EkPTzm
a42g23GzF8qwHDHPVNdK5sW6cY3dHZvBwWEg/E6HBbnU6GeXdSMm1bKTCVselXuMo+Qldwn3A3q3
E2UYHVRq5wW2b6LiH7M76tZw3t24jbnKceXcQA5BtsueelCrRpSJaZQFs4NhQaCp+3lptSLxYGx3
ycK5qp3PjTxSVzZspzoSjrnVhzbSkM5prwf90JdGsH9Qh7bmkW3qIpktpgNkWKEv8BWtno3653p7
Fin/wjA8KN5u4JT0fL9EiQaUJCAF29atwq1LFh3fxpvIq/7BjfrsYmTi2dZz2LcMCix005r9y7M7
XHaMT2mlkuwyBOYVXAA1pQOc+wxbethCwF3Gv1Evy/QEIAwlJSSN8rl9FqknqERVkGZf+hCMA49t
gGAW/vYNZLk68pfBDVqZQb4pH+vtNYc94JQ3OzyShij+QUA6SihkIc+bUKJasEni96HyZ+RuJx4k
jngtCjiP/ZTt9u4SylxKSC5zMFtcB9t+vPde2vRyTTuO6/HvG89kKZtfe6dOZMKZ7IXMNVgbIDhF
v8H6U+oDlbxiDTWS+UeYTflXtC3uz4LqzjaWTzfuvQNNwS9j+UvGdIy4UTJD3qnSU34ZIQwXaw3q
deHKYVyKHuPBYX4w0soq7WatNtZL5yu5wf6VNT1hBDsw+uurwKy1KDOq9WyefKYQIH33a8PvuTxc
6cSDjDP2Ynhq4GYUVPJOvOK6cjnro0cuPuK/aeETebmAr4RmTSc3yBTJLjlrHQr/lebyDagdxwYk
IjMt5OMBnh5gLmJ3OTKptB3HATSnCRl7w8f5bJc2IB0keQUQ0ib1rlYBWgC3ro3SqLuYWb8iXnSp
GatE02M9Tb4WgqcAh20im02zpwsEaLMx0whaFu8NSUT+b9Z405iYETDJGOaAbVnQH1bmMkS/phtP
V55HwBZM0oAt1T91+qXYpT/wZ63DUbFcJWaes6YVPOYOBaYPwtcMD74lVtND9fNA+/lljH/F2VRH
0CUjFdtOSgp+SYNgQTIct4vbf6codXA3HGXboWAFjkSmsgiEr9zdcuCi7i82EebzC31pdw0Ju/zU
CIm+ITF3m5h4GPKrhQEz0gg/6W+iQ6p6wbbAZhPdDMpBYhvU+NUP8bMY4DzTIQpvOrnCQfG3gAv+
Yi9xIDwtKgcJ/91VxNfp2t2KrTMwzTRJhBL7ub9mYlm2tA4be4UjCv1qzuli7qj3HbjguXIpBAxT
KXgUBxrlq/jzseQG09mmCDrlpbuKjHm/2fAc8aqPW1HNCfVFf+mow7RApl+Cd/d70CogvODiY7Dq
OsfWXy0OZkMLD+Skq/ak1cO01lQzkd7yS3op3hsxBVHmityK1UDCJOlSNWEMklFc4zpkj391yV5c
7nvkE3o6m7tjjf7ry0RLaUPol+8QgiP925uMUWDLxPxZYwJ+D6tyNqKQcesk8C6QpDIPf+9UH7Ua
vIH0iaqy/Ouy+lpAckDpNqX8q1xd9ZDw70nLMX/jTy1KHBYp+PEEg/WLZJ1de4PvP5aMWWyMEx9e
N9yU25DlmAfmc5N1JGt2Z7dDbmU3iJ7J4Edtb2FREgqSiSmKKVchBCSsXSYybLYYUqeq0QNJQpms
xjxT5iLELbtEMUxkzWqHxpP649BRXQzJw0l3pzUGPrf1B7BrNrwXlkQ0DCQjMg+uJW7aZcZz3r0L
iip3mVMeLprmVInLtbHwqFtY0QZChZWUF9bxoBzgQ9PMIlPYUTJNBN/yleScvEfjd1PXhu7K3Sw2
7/IM1ESiiwQuMQHuB6mX3Wf+Z+aKJgdXokn75tm62NfTNxRItvyPwwkHCEvwDVa+PEUOay+EfOZy
U5jM75HqJ1daTx+aTfLRCstSuq06XlKocwY4gWeZbrKvXc6oob+7wFHZJlS3itrpWt+URfRudWCJ
bvLwt8MDk6xOqAEMkELkoRp0SzX9D0qG41RTdcc61qOj4AHUlpDLQMOvgTitxuYL2gTDjb8T2zAH
bi1na/AZ9D0MBmBMJVflaZxpM5CN8bCIz4/daNRTqn3XXSvG7emuY/Jr3ep5V+mdeNdWXQP3WeNe
2IwxTwL99CNxy4d844cLDMrP6s2QwemDpHzD4YfHRn2rimeHeZ+S30AkgQliqGkfkmyv20WQFNYO
DjB5qFcMdECniBfnyvwQYnuUa7bzrARLHEnwUe7s0VnFXikTQRJrO4FBN4dTieAqiReb15pmZufT
BiLi16YMaK2ec0+hG2NEBu61Cdo0n0+s1Sws78NQmXNmv1pXXiNhyRgciq++hqwkQE6pc2NmmMKB
uDpLvVNX1Q/BCfg6Oac11Hm9Vh15z192rPTYVWAS+Q8j6KSjoRMoULQxcWqIql0uw33epLW52p5F
XCuG1RRwbheUaArw0Y4JkL3M909dh4EA0HHk77b4eFK4HNA5F5DxpEVLo66aOgQ/vhC4iU5/KaNV
SyE6KXzjlUIVA8F0cd8/gZLNvs+PNzVOgMcz5lbaRnDaaMsNT49yKZ98h6n9f6V6mSlvtYzW0Fil
WQEaJBjMjV4lYvWRbdBjlDqKFHY4fT7+maHYvobWps01L+oqCvuW9fLYCgfonjGi2ny8IJJamjps
bwdhzJV5ylXxWbjvyDVGBkt0ZHvfipkXz6fV824fSMtxuZ1BIcZBqgVrvh5XwYxDDaKVvulLr5pk
E1FbRmFKm7sLS4aTwc3rhetOWGrjemzVTfgqipRj4XyiM8ZXlPJTJBvLDbJsnBPtZwGvB7Q3jV5L
kFyW/gBhc0KzldnL/R6J5PDQrXjucI/MfSqRK3YPlfXcNVj1HCWopVqFc+Zb+47PVh64iAky+Su+
Ul0xI+4KYIlAm9T5nvU4yI/V9ZPRLXxRH/KXkiyUlha1Vdr6p/8h3f+414vurE0D8Tto+o6NSsFC
mNxkSninLCp6DhDD5bfzdKxw9cAYykYnCU1NRwshOsYwNv7/HAXsYPRHRxMrfETx3tMke0fRZuQJ
YGw9S+nJgm7/LdgXFBtk4WVH5oxgVgk3XHJk9cYMTftYjdBe3ZiLlpwTF7D3p+nC6Y038oKrj2Yk
0iyJjxQY+FlrHfqZrzUc1gfQ+pzZTtO3CjhJYeWItWm/fOrOAcHy2eO0YNw+Nhyy4XJ8LfViUKRP
fHND6qZwLkecztuJRD7jgMfqxifWvL85d6gaP80J6dQWnHc64igMQbvaThIIoNjd1JVCHJS7gTTE
Oa/JMJX2nYT+tFaBrMjUXccFVU0T22G9w6q//m+Ch7WxcB1lCBrOEK4c3+9hznJxfvRkoV7IUZk5
dlGL5zJz8t+faBZ0VegNZypBr2ezOFIDbR9Zjp2Zh0lhEEavqnR+ccnpnUdaXWRblwUT5191Pfhk
llNjoAVU0+bq1/HJqvmAB+Yh4riHvWZCB/T30uHCuC62CwSqgWjWcpVRF8xizKtn47yoK7/SDTtK
DcQsmAB1v6TRxGd72VgjRPWUgehQAiFJARf/1u3s861Ihglpsjx6pmMPGrrp5mbqDAGcLb0rnqwI
DFgCh0sT8asWYgDTizKHXyKbCmB3N//k5+t2b1XAqrYbZ43ak27aOPtAUzbkPs7y1KvBK/ezxzey
/EQSoPCOOOqodJnWdhrag52YXgLYf7IrvnAC6Fv0lLzQcWCWBfTA1CxFtiHXSmgrYtDqtVpTIdDC
x+9UeyQswGkiwdTWkoo4VVCiPFKy4L1A1azndqldGoUUIfH5cv2Z77PF9T1m2qEyHYpqKhyl8OvY
Y0RARYiVzR9t+kZZJ/Z4VDL5EoqvszAX3l1+XOvbF0iEND8ktk6kjZG99tiFHbBRLsb0xLrq55JO
j9o5w4eojjjPz570gDuOF12DZsXrFg35UUh17zchA7xJAFc72sNumD/7+3JYU7h0y2VuEVRma1ny
S6NOjbm2Vo+95EyL2Es3CIjt/uW6WX4XzSPyS4JMihi0pIvpMLQHY1teK0vxbWLxjEfNQdtYA3jG
VX/sLlL5m86/XKXuAtpqdZvujx4taNsfwryjwRT+rUpLhOSRaZ3nAYN6a+bu5xgmuCMKXsoDcpXW
rC9I0ZhXNMAcOTZZNonrekTlQN2z1zOpC3Pt/mX/h+xda5kAeWremwl39jjVTnFdVn9rou3PucYX
E6v1OzJvv+38pXODTCnSKn8FnlFxowROsOUz8W7zum0aTXEVBA/7B6pigP1iylulBovcKtzeJhmt
iYllRDBiz4tbO+RpD7cdLXTzo+N7cAEyrcArg1Op6jjBUomg4/pLSinCHEEGOsgOe8Dc4BVsNgb+
1PSJcY3G+2i8hYyh6r+cEbKzXnM2qDv1+VP/Ln3FrBhtCiB74v2qKEBUkWFcoOv9seAyQYC0mIU7
ZIDxEAdBA9GbynS8fPD592AD5HgX1N9v6OWw6Q3oU6fgm8Ke3pqqtnrAycqF5jHZO35d6rCAnEcI
SF02hjsDweuvmbk2hXqi9jtp6z7itR5n2eA+6ymODMoS5WqIbwPNzAUk9Q6Zjr4K8owK0L4VFyfu
w975G/sS7BX/CI+vO3mKMkA+b21+cWCI8gwZhPjSOE1+oT17FQKLjs+SGAzgv2Hl1uvackE+6xzD
2cAdsOFksVzUCvmjsCndjeCkrCAhpOvhDZmaddcoRZLfQakCAf4FgKDdJkozyHcI6l9boX8PfoOp
/kCyLQWRF8M+hCOTRnWcgs2KygnDoaQNeU9Ow2rXNLm+HcCaiuqxgeyjm8nzVgEUs3WTQJXjjoCo
sa5KSdCeIIta+GN9TnfcVSfJjUQjeJxCS0qVaJv1ReKoMCWuY+KPN3Zn0zzMkhm//qnH6bTuMLWw
MSV8li+tyekqrSh0SqCFZNH8A2K9ntVhD5Tq6GnQylV5Ttkcqx+Gn598cJZwSw9z8yrqJe1dVJiq
IAJ+eHdy1qkOUvteaUkOIC1788Mmhq2OKxfBUTKeCAXMpMIzqDOfmJVctXk/nRxXRkK4VxXT5F6K
YlgvF+HjlgP0g5pTYp1nLpA0XIkYae1JaDIyQL97Xynu6LOqrctJoUCl57hS1CzMKPV+RXi7rBJp
Hzy+yVT4qqlUhJYEOs8/jb96kI2xJZXELse/IWY324LW2si59M2kPYvq3Zh3VxGHxPrUAH0J4+W+
GToI7gcjcaM+usq+LTIi/2JsKPofkYQzm3AunkhyPBKoH4nm3OWOVTCDPUON+zJaKlZq2Hya2Dgo
8Rt/hrDq8i46eN4fUsEZRBAodbGgn47GfSo1rTvKlTxf0ZHz+0mlAfvukZJpxHbcdqMwoGv9pTrS
GzFlDG3v2unmzBsUaFff6Ne/9A84dQkpiizJh/1FCea9/5FqvyZiN9xN67pQ12eXg2L4Co/QZI1P
FF2Ga1s47WFrznZaJnJdxxFVeAgTPN+sW6XKnMxyTwr3P2HuqMedmU3V8YRFCSBhhjisueIPGoQP
xiML0JW3DZANgeCy+tlmzJQTZvthpDUcn8DbMpKk7izDWIQdTtcOCKglM5FX+/b19p85zOQYcrEz
gJsWlny40n/psm3XT1PGuiasfkfEKF82Cehd/S/HQV/cINL+rP1S/yyJwbd2D9e41Wwcem1017BE
9rJ1M8fpzmsasVZ/fep3+1oR9EvSyNYJPmDm4p2qs3WvX2a8CNpxItu35eDard2/IHZBwlViTky5
jnL8b+7atWhflR/ywY/TbSC2aVuyJ8wqalJkPOQVk1eb0Dt5iHagmr9svdYuQpTJMTRvAdxg1oHR
POs7XP6xtgHphMlItGLBmbWx9mm1WuZwVNMWpbQuk3/WqIcKBpyyDVfh2GxnkFpN/itKoxUQ5b82
TQbsehuHoXWoSx89A4LkxYdRjU2JAeNCJPJZ0oNSS+2vxV3NWTTl6VNFp1rnuHHiaYkke1ntmH/I
QlyqOXfBOA67CG320i3GPdHRyBJlsxQq9Op9ca2o88t7xrxTmcyxnwLMi2HCTWeFjFoKRxLVTCTC
GE6gwoWRnBOF3jB5gzgFGTDhDRV8fA0WRlmHG9loT26e5QLUkEKBFAKPEwnPuj3yDfwQ6Gesy0b8
fptmjtewhfYG8W0X3e2IaI+jWL9c3QJ1P1YyJP1OUx6i/d239EzeRomQpU2Xkel+apAplihskhXP
IPC/KKztHcou2pfZsPzk3WPHkGwRn+kt1SderC43y8EpxhoIihBiEDR6lq1+FzoP31cBF0J9BxRg
vV4G8QR0Y81AeCnT3/DqVXX7lJuAl8E9JWusfwu0lo4+VZzp9sJv3UgAr2L9/9zhczVLEyV0AMNl
PsWWVYHILwJdtS/GJYIIqEvg0LB1h8n42ZBJZVAr4dU3ETDRsL4NCvrCSJAnzUcISRHJkl51f43h
5823+llPgzEURD+9xfxnpM4/GYpb1oHTjA1ntOdasDowm2Kd0B2fHY+1P3ec2APnKezDk+tO79II
fvUetaX0e8AMDvclFYMQByG6okAF4Ju9uLyIiJv1kdbqceYQbaBAfpsHIKmMKd9CD2m/Jx36CXcU
OtgiOzIjIXa9Xo3IKxlrotZug3czKdHcL94PszLs0yEYub11ksBAzIhFGSCge9SYGOYgrpChNI9v
0Oay+9kzCpyyYsxO4Ax9YWuqkDsksTAfZxpY3EMXaSBpIiVDghj+gx2zVsi+Dx/jzVo4kKwU5BZB
u3EgN2KhsfFj30YRof5EnpkpaDM6smFeRPXMFPXyee69viefOa+CcBTLl7eOAPnpvR7A4m7Ax/oU
kxWlD6FFuaeD0dJExipQV+tXSQm1d7S/6zhmpLKLWpV4BjxGYtPFbgUJW40OJ3PEwNAI6iQswtGE
2du5H3lx03D1xj/QlUJGgWBBEhBztYTE1R62b6PokUZyMqHU+PFq+9M96narZdKouKN4nOe6yrwi
WFFrrqNlduoQfLhN0+AupQ8uoK30UUi9rp+i0Vz8ptaK13jrulphjKQOhaZQvzKWom+JJktwLT0h
IonbalvaCmfYkGVTFS3q0o81NJpaA7HVFC/cXIOZFN4zLETjanYie9getk7FgB3o2BKRqZveuOpc
aHkBngdI6iGsnK7R4C4AZOkZftpzzh9tfkZSp6/EfexcxoeFf+EGhBbICqWW64amhDspnqEBqu5u
iCVftNBWONQVR+b3TKFUiK8PF/5V5Fk1Db2kA3wiCmZEzvocjVNPrks3LKEQOJKYcZ+JqWcM7/Wj
s7MFx/VIfrSVNLDa1L9+XrjQnKzmWOg7cehBip22t56QQ8YigwFvUXh/4Y4guVmPOxHKEe8JoHOR
WW6P89gEb71ncr9s07Ag7XydH3/T1cQPWPtQwMR8LG6PUU+X3GtxrCw/jg0lacpRgm+yE1p6Wdz3
gW42mm8UO5A90ZBzyEoDgIPIQSSFe7BhhwMRvAXxP278b0gI3k0PKPPFWtvvRg1+AC8V/jXj5A71
AZgOHH/c6BqtrQdZdCDHYxwZ9ZnFrowyOZtRTg+59py+fYCChlFcLmqoNNrTiPTfoKGioVo0wNED
Klj8E/Nt6YvMLTEtNo16QOJBM2Ymtr99eHQGq0sITw3xkoFlJvUMZkPiZWLkOKOBHeGlT7j+y+nm
uav4DDeM13yXUDrc3BVKjVBauHkObI3p4ex63poY2SZ1WMzW3nCkfSlP/uYSRhlINcKeNMtexJqv
eZKSuI3k193Cexei5v94KXSZU1houcPjxF3nPC2wy0EZEZeYb2zHola5vUkouBKUoacV1ZCyFMdd
ZjKjo3bA/AZCLLPJnRSRfPqkgyFVksi/ksb5ni4bSaFhx8AHb9kAKLekYw0V9dvUoycX9Euzj8Gd
ZQpZ0qiRPBxy8fsXrfWV24TexJWx/xrU9vGoJCgjk1GE+BQwG3ZJohAWV3qOoC7uoT80vafoCY9K
iyGJWXYw/GqJYlhy9lK/P9Lw8Zu67fZLhwZMEjj0dizaXhuTaqe6VeFnUTsuRkBelvCU4gZVzvI6
/cSY1KTaPDM08k0+jwmVZ4OUiPgJcgiYJVWqdK/fGuHYsPIxNWYHgJ6cGoV32S600rFM5KgVgjNd
U5Z3gWw3on1msrh+MOcDWR/XBHZWB+cNaymU/o90K17pI/z4UJ0CD+vfO64xb3zp445i/8VbGbEg
uWgyL3qD6fkK1/5NviWqqzWyFThbChL0vTuIodJwiCyWOoDFLB9Lfgzd2zyapqKy4Heejs4fUViJ
1YjxY0TK9Mspj/zuPcnVudyZNENLGGb6hPeALm5v5Ei2Axk6LYLwVQmkX6JKXu6tEUMBzU9KaVyH
ZYBMMCqPQRdlpFgmy1U54nXv2hu8a5zrPzcBdeKsgni2o3/wEu8QGOiur+ga2h2DNsvugT4yczQT
xjMD0RAOUPbYM21cB8KRwPunGPpD4Y+FdFEwMun5gxGLIqqig6IqA1AbQLk4HlSzvc1m7R0vdujC
zaqx+ktC19lYfg2UfUOLVaRFLwowX07emhik3AD0COMgILsQcHv7oL2z/01YnuHgCHYfXw4T0NZ0
f7kMXEvHgE+PUri7Q5ko/QFt0EHMJK5Pewrna/cJHJBoqRnb+MRnjvtkkhSI4gWGcrt3bupEPcy3
wS1D3L5C8jCaMmrH2ASl5MPyae3y3j+ARYjWS66v8vV/DGebXrqK29a7sgiE2sPrlWNil7CYkVnw
E21jZkaowDL2Ibni8IMULKvr0B8JCsKRvh61MN7keDFzR6QCQActiL1hzkVwwuPBZgJC+XZFEEKC
NgwoSD/nIc6MXyvmEbIgZg/wEMKjdp/GXmkd+v84MP7aWqSkz3bVWayxqVVFhXWTAgef2fuV/7DM
jFB6BGtykdN1JSsIhzVTKhKJ/Ek+sb4ffTJa/DXjVtT8UobM176tlLZvfIc66sWKpVnUX7RN+tmD
hCy08l3uZwOqS3fufniXkv8QtXcH5ZwlnbjXC7aggqSneQSvdwuiWHdVKIV+1PLARnG1BI+bboG4
S0A931AYhUyFzNlmGEdjv086LbU/B6RD32i0w33RWbWi/IHCmLgvygehkwMpVJv4hBnzykKeVcTt
+MN+nkTa2ddcPqBzqOjPkQOKg6clThSsiOLJG9drPx5Hxwf/SczqeGwKU3JlPvMsRdEAyPzvFLfW
96uSCYNvmiPh5+JD33ZDyOPADKaGkFplw90zkPBVnLEdWhIuM+aB9R3T8IQJgrf4zp7+5e8aavh5
ytpw7TS6XADhOYl10Xx20xEOjHmW/7GD7negw0KBzRlnn85dwl08gQgcBIAz/ByNdbWmjTHJiC1W
5CA2KXj5Uo/HOS0RDMZhAysjiLbcArP6uZuiSJMWQcicsXbDtBEtseZif060Ts2ZINrsKEptmhcI
3r4ls1Vy7ekZamiUd60CFte4YJ/uqwXXdKdey40qcCzSAxVxoxJDGVDfKk1XEccPOx/Vi/b1UDK5
TxnX32ACuerX9xCXuZ9n1n5X5jZuz8kFmKtSFGO5M6+1ES7BPvjZ9Wkhy86cxROGErMYTrOOTynU
vGpCRxAa2Ib/+A9L06FJaVtyGEgBQc0kT+qSqn+4yvsnn9TC5U4hZWpQtwD2k1xCoqs9xoQ/MADd
YjDdgPvAXihO2xhAeYu8wWBfmNAPu3o+zvDEEToYE6j1w/XSm5oQQ+gvYxn5WbboWnFPeuXqSNKw
zhgA6fNjvmB45M4gESDaVh7pBlaNAsmhhtUc6pvbeaT3PGJxZj7XrRgDL6z8oPt7X+T5YfnbWQoJ
8wzBqs1dLqWN2lV9a8VAbXZp+NxSMocOLY4DVaF+xdzuwwLycP/6xw+J317/iT/GU66dvvQl0WwK
asl2GMq62x0K4E2dLC6iYMPdJ0BRvgQA7WUvJDq816zZ/tebgBXxFTdbeqyvsjjkYiFaHnzvjqS3
DANzaPIvqkqc9VM8MQj/V8I3IGbb9JbEdWkEAxCp+7B5yb5Ak7YdSUDIMftudL7aioJfDHY4Q0aP
dGx+ZBe53LP+RJjHSJJ91Rm03ljlEsWkGNovl/SAHwcB2frlJ/OywFULWAD7qIyBm96xerQxSYd7
5YJ6t2//EJrbwjnHwQVfujM9P/JkH7ab85dWewKZRzQAqU1k+/rZsAu5EInlH7WaG+jTUFbgcEUM
vr/Gk0BMT4kw6EhG2Ze1v6B9HvBlFBqCGFtZG0e1liOTYvNdBLpzxMRjajlxKskGjSctaci48HYL
mA9wVruSi0mdZ02TUb/ZiUayZ+KeJMpTdNBiMbrvjsfTkBWtHTeY3Be1y8oVBJEyG5kXqZLYvHmA
qZX0puqdzvW6WX0mCnh/so2wG8lPMk+2/uxqyxSTmO4SnOalAbrzmBwkx2WsLfBvbOJJaUQYYCCF
1l9W3Hg3v4bGFDahjfnLHbLWIOkMoxEPk7wFnK4v6WeuZGDGVeUr0hWdkPbjjGYhvXe+5f8vIXxN
6ojBtaLpCdtU5Pj979sJ5qW0GbqzJYRUs6viVhCvd3Sz3Eb/2eJQdJiYwn0zXcjIGvTNrcEYnlK1
v2CtIW24rynrQI+1Zb1gpr0SKk9dyb5Ahos7xMUPh+igybJ8ALOAhW8TAwkHaUDH94vJuHxE22Vs
HdUXhn/6ZMV2sIdzDJvii+nlKetys1Rik9ydfobQ4j2t0UxTNR8Yy0KpbBwYqhMpxzlRBa4YSKU9
W+j2IoYZhPit7bIF/LqZsa67+OG36ecojocMJooo4zHX6Xaod5brQPysXse4rzqzJ/wvggZqbyFD
L19G+gsxXIQlNyZxwnjSwJUbQgpx+wKAb/U2zbsSdujvaZsXoXvB0OIEUzhQBsnV5SswRYr6PzUH
pSLsJQ8XonKMel2y+T6/byOa4H64e5R085sik0Z+OG5DBkxO1RsFRwWKdtZ8HjWu2obapJ3MYmde
PXqEif4ZI6RrXfn6vHun2Y2Z2MrjCQ677JqAGsWfRPrfNnALfwCkZv8wywrN3s0gp1Ttu47tpv1E
iZDJW9C7pSoRsBCpu7Mk7nld4n7hMtFy+SQTy00bZ7QntNBbT4lAaHZz0Tl6r3ZzWXyJTXN5Fjr7
nyudf6OV8dJr6r2aBjosm65IncgUSDlAHVmkp7nqzMHN6SGg8SOmgMmKp4X4LxWTXTtPYhJOpiLB
pp5BVNLTwXITk8MbwE+UXViy5JDD0zTGvljwxsDisuth1pvWi5saGyiyu84z64m9di5VUb09stmk
uWKthhZ3Ylzb6sEU+63KxIkE6jT0HWFFrhqttpcCOt1RehIKAn179rrnzVLpvknJPmH0PSXDwtTY
Z6TdSOY1KJHFYhQJybLcI2W4pxQtMzyDd0+rIergTz1bQt7NMqWwVBop9t8WLoEcWqnRW0eXDmNF
QSFDzb1Y0IxGN6eamiOWaoAf/J5tgLnZoOXsTX0R+++DDw5Vl7RirIq8NtDfIBJyit7KUFwuw8Uc
KVKVN6wVsC7YKJbS7rhsdThOxyYgt1YGziPFpwelF0629IjsLsL0Kn485sFn6N1FDDfcCkesYTeX
vu02PwPtLOOv5zdFCmU/uUxkMoYFKoDzIQ84dlqiE60+7TS7ELNGOxxIYeRyPmHfdohoFPcL9UE8
cLWpYg1VYyKES2SdCXbKXpr5uDA9h8DRObRV6K/mS7NcqrboBS5AAGxvxrlvlvTE0fHyRx7uuIBN
cSjVZsUa3h7vpioHCxj2qAXxl2HF6kC+GH4g1RPhPmxaeruNBETkhU1Lvmn29EIhk1f5EO5t+0M0
zXJGBmFkfA/BuaQhpZl/T6vU/bEZkro0keIHBepigpzkG2uKKXCwHyS+oop/6IEEt6SC8DtMUJzt
so4a8eUfUaQK1JJzS139+9pUsH61Uly4PKd3hMXVY5SFyXyGgepyjwyFzdgy1zzg+vAOb8uSvINm
RpAbDVt6CC43XPne+K8aP3cm13c7IlR407kAtIOmUBv4b+hWcCEtpND4KXdiCkbTTClq4tdLS76J
gkisKNNa6QN7b1CBmd+6V86DBM3raK4auzamA5PmuFwjIOIwLHwsjvjbOVJ+0czgP9dSevWJ7QQh
MB1KH9fVUpwAnA976y2tCtRRpKGBz94v2t9w2xlr4gnhl1kVy/8S8UbwDZiaq1JMZ13ksKIhIZ4S
noQEDmDo9TxbOSaUMhxsgC/72yL7wfoVSFMuAuLOpD3LyB3d2hOMixZeytW3BIvb6rzsZeDuV9VI
iNN0j/C8JqaGcaV4NcLgHKz06HWEeNFZawAPAeWwlw/ly89W+YjTH9BpnBHY0WUkr8XiTRqP3dlj
6/Eh2YSSxrcV0ThiNm5M6OBkqQEAqoIGf/yAEOKoCH5rIWgDpfQIWQH2gXXNR0clA/G6KTRPTjkM
uhu7LoyBnm2QEQ7n28WEJLfwAixBkXvS28y6YCR2Be5DmfpxFR4qgZz6r5TeDSMnqBd6S5GcNGyz
p54NJ8G6MFNwEX4MjBW8/zqJB54x7/yEnO3vc8lxYsv0o7/NlvVcrGDUPd/HxoW+c33Cn2f/+PGo
rtFWJvZin2XWcM6Po7A2E1AA647X/M19Hg+lcgK5We8tAeCBhvcVLeKH+DMGxqPUQd42lL3in0QV
XLn9XpBPpBGCSw5cGrj0PvkBOBIGnYf3K/4YXIGpxn1lPNwwgbx1x3tOmIMhK9fWkZHOmtfDPXY9
zhMT4uJu+3f11LaYr16ckaOHMG+Y63RcxR27MLRX2ZxNfC6t/JSLic9nCPXL1sasQo1Bcg3p/xLv
VAY1DjcpVAKTkIbpy9jJlnJNwPhiRF7VocLwbEmRD2Dxb3T084JqRprzyLjkBHgHNZ7Atr9LIjG7
HctwjKSzJu58s2xF1EXwfe7je6Eie/Wt9WnsQn2ubQR1pfVi9DXEH5H+SP3+sLL2WxkcLhMI9JN4
4G0mXJYuL69MK/jAeF3P2UXZhui7p0RgPtI8tHJF+zGjGoAifgSkLNkAGXJQ0HzZwak5sB+4FzAS
0ynLPi7Wu5JTF7OnHjRRp9txAHkAblTU/0PcF+jo6bGbmJ523ND7TPyDheRkJvTDURzQQhFR4EVv
HMJKFJKdNnLT2nHEJTopMSDj/x4plGe19p/ueGclVPewC06q8wei7ZkI4gK2IlMJ2Snb0+6N0cm8
tgoYztZrPfmW+TqJSwF22R1CqCr1hAu5UY9YjDmDN4Qd+LDO3W9Kv8h7ubBcIh17ag16KWmOgIdw
v5p/wESdNjtpLqD9yDbMfBSO06hgPMeRCIH9G05EznAobNrdLsHukJza4vZgK2KWuX2OkqM9S1pK
+Cgd7/WaYTvHZz8Ng0VgkBJGdarc2QGDO9FFivmN7CUtkL5mvxb1s+fHoYrsapT4E+cy+STat9n9
nJ/94bl0sHgdhW7Yw0jzAmMmbiU+QIC8bW+2SsBmTRFPOTRGdyIoy8WUwRiQZsITcZRKKGr1oavc
8Cmduht80j+QoO4C4x+Wl0t0bFZ5vy+1FB8JnK8L78e9epmz2Yq/RuEHsRs4k3zSJZfH3Kpf7g0F
bPVcmJfpm+8/W1oINVGmbnsGyuptj09KHmPf2UWdtb1xhpjAVXSCLhK0SEYvTaTVM8qbNbWTLgro
MuubTTBPK/h6Ed9ZWMkoZQK6iTCUVxGZPJITJRl/GKmUSzx/TBU6Y7BRzMdASA+z91RkI+xJdEtF
9CyzZpkG0l8ROygUekbtjaxWC3F8/sd952Bsr43WmUdiN71O72ov3pxvVuxhnfndJ/tFGOe/Gjtp
0UI1DrIrs1fO1qRvuzoVC01vcHHuHjCzJRfIIfKBLjGa6a7JZDMu2jlD8EKpoXY3LUiWutEAsNzk
ZkgVfcs7G4ViMh6tOTKrfn7+2XJp12G3LciXFVpJrUi5Hu9s4lZn32bw8BcfEm4uDuBX0ZHWcX1I
S3gFhS09Cb5O2/YqEIg5AFK9NWReV9hsejHer8BYrmCGvqLgVp1n8J2dnUoQSM298YjePAQ/r9ud
US2F6jC7Tv6wnbfff8K6bukVkvgNLkG6l0h/GWO1IZI/gRdM8GAtkN+p4e3WT7XmTPHyZV/5S9GT
rGK0DjAQLgaspcJLqeBnXBxoxVWkl2xobrlDqlSan1Oe0KbqGYAaMYo5nU13mF2rQvLUJYT3ko+q
IvOPZN8wmMUiSwasAKLVQ9HkV2Yb+K/v2Laf/yDSVBnLcckj+QSJPiAcmRYxso5AW2z8hr+DP4mS
l3frSKJgGq+zDa2B/vPQojYfvAWzdsOpbkH6S8f2gpUP9iwCuzJ5WFrp2w+/QIEICzCr2gqY3u87
b73D9I3T5uZH5wsFlwxJxHWSfljaK90z3B0OVhUy6KkOWlLY5/LLaT8g1vu/rJYuVUDaT/jtWsa2
QCt65F3/MMAktpTtkZHnfnFBYoWMngwrsyWvhJKVEGS8qcjf50RG7GOck6EhKHw1cC7P4g+cb0GO
MdrODSshR1J6b2uZm5Rp4RGP02/FuMG634Gz5W2jrOlDasUB6GQoRt3SUh7XTQYAk1bQFiBfQPrP
ezbjQg0t6hCMFcG7Q1hKC3vAmo6LgaY2ZolJtm1xckY/VmmWSGF9f3PuXygc6HGSpEM+9eCrBhqF
QO6EAEPdC4Gw6GJ/ph7KCeQVAEQon0cRCOFGlobvEqzncH03yz+UrckIt6AfHAfBvLOL+8wjaNZh
eKczd6PT39ZNMskwXDSrraxj924MBRFsU8B36huqovIUgJpS5cC/5Xk3+/3nzlEOmN61EbV6kkBb
uhoMTI6A6B1P4gFx8mNeyrlF+ie6nJ7V2XIsq9eddc8DvbVEiOnmMGQyHTSx2yKZ5MVH1ru1PyuW
0BvQOpKKr2SyW89fFRxeiiSuUB81B3xPLEoLapcTUGlumJmEiHFqR8MrD90r1tFOPtA/ok+D6ypj
6ZF3YDx2MNcW5XAEGyVljOMxOOFyy3PKsAe1Ja3G+QXmShWmoNtJn2YPYghc+UzBV9eDe8OvEN1V
F2JIGjscbveh7giI/ECXfhuHLCftUTPEy0aV93zG9yhz8SeocjvjGoqMFTl2js/PK6OqhxxpSt+9
MmHyNIBqqQUoAxzgJVPId4xJ88+AY9Q88cSv0rLdvhiWDyeVPodbsCEgBCoHyRZBP/qa3RvaMMcN
uidk4jbS8AUX+ON+e2ZcHbAWePD4rF1LBAq2yHNsnfXghmG62taO+1tWmTMCBPOALc1MNUnIgbzC
E0GRe/mZ8mq4pHS9+JPjLTdtqJKtVr+0XjS7xOuZKJyFoejHQr2TJf+MfgV0r4VPS7f+9+tTKVBp
rOSOENupJczUuA4JdSMNdmdZpFJIFfAwETjSQSDf6x42JHQaZIiC2RGdpyGkwF/+KlKHcomL+X1Y
WtAIF+lkX5AAAfkvgvNMNBMhiMoxHDxJ+FlsQ3HrRsGGotHDwRYWEV8MU1HVleMraqV/xpQYdijq
UkxVV8Z6JygrF9RbWgECIASEKhwpiE0NX3AtUUuPybncRNbBZEsSJIPH1R/msWESL9Tudb6XQpVk
DEiV4RYY4unx1VeI0gbI4tsiTnPQkElMSiLk3w9AeiXqp1iWQwSr5HutXrzUaQ7Xyz0Z938pLN5p
3iBP/UoV9YUtWob2++XI6WsFgbYSzFqJSgauMl1npswVd8uuyc9GrEnp94qYEQFH/rOK/pn3K0QG
k0b9wShsHru4NdHypHdx1MJVCtVL37XEDcfGZkl8i+5Gk/SsEeminf0YvPJr+fQXgxB1wde/3fY9
ovXe2yDJ8+9WrQ6CMsCrDZX6cMSJGQ7yJ2n5iHXzP9fPqSo48Ci1q/BxYUaO3kNKB0Kg6feHL2mm
H/ohwHqTuB3uXU390j2uJVutI4ClxF7awTc+wBjgcoaoznokFGuar5nY7i9g8giUHlLrilPiV8+3
oeTmYpIfVWKF3kGp6TQps0NrQ30vx2xsqrYa/+5/JShpfodh1d9uPMDPd/P7Byzvi2/9tVF5fvDw
i1NvTG04ree+k5xQhiFXlIS/Ckp9W0FtJXFEholaO9d0nGD8WtQZvUqjSqHlEvJGFX0Pmd2d06Ug
lXfA7pp92wEPF/KBaKShsGIMmBjXVqjgtY1MooK325jmh9aqa+nPmtsqybMvrijj76IwsuS+Ge7t
dS4UUhaMZdbBNJfbvXJ1Vgg46QFhT431Uugf3PE4maAh2sLKA46oZGMifSGx08zvXCL6hG01ZkFA
Aa8zA86XD0eSBgo6pRMH15+VsYe4YnuwArDNqDruU1CcXjqBB9ZuoIF9Uk3P/SebIMlulLYBhE8o
OddxYCR6z7POruFhAdw4TvAXoK0N8oV0FiedUw//ZeZYhJDAPPru3sc4N3aGwE6sCo9FAs2RUD12
ba9ibh+rFlen2paMoXJlN0tuD/3OqC7pE/Oo8XvjEZopAQg6UDUxKImEG+gY2hFE3WGm4oNz2BVz
bYgq52FKHQJe41R1o3qr5m1zU9k1gfzMB4wJ/PgWVhveHcgG6hRXSyuKVZi8nzegOkvOYYpd70AJ
PPhFZAohs8zvA9VHZAMX3w0SaWYy40vWN/HNNrB/qLolhxabkpONa56xMLXGMUbIJZ96JxaWIN0C
agvirdyJNVejerrqLSH8P80VY4kwit5uBONxBNpHUMZcy3mRhDTPO8AKOhuVQkM7Mj5YL2S8/3lJ
SA7K+xc0DrqyQQAx2xruu3psU3Xksec76mIq3hUDd3YvONiYo6dLv82YnCZXUrh3vI5RmAWTUqSy
dS6H78L4jEjPBggUKgarenmMMN1PabD/kt6nCpKdJrDSnK3N//E2CfEkYNQ/x9j9DXKBbKEnyFx1
NikpwBtHnnUrkfJOMKF9E/O322slUjptFN/VVxyK8wCUbaHH9EnXPqo3CD48Z3K2ZmNjhZNVqI3h
ZvdyKcu5kWnYf8Mi2BwGuL5Ygoj9X3aq2rPfIr4/iNk331i6fmTfl16QRaEiXakvt4NC9SRq9QUK
q0oNnyIH/7k0Zi7qXebAUPWF9ddinq4GNgNMy/Bg0B/shJOJIhLvE9w4n2Pv0Rnv/fMjpmaSsQsg
7lWILo3u5eOduKbcgSBeIHdkPCtnTBs+y1VN0iaxBMgeKcfJgMbm+ZhIArwvly/jWfTl0FgAelAW
Ry2tLvHgJDsu1MM28J3UOri8FGUS4LpqO9GLGxOk8HCvkWIW8poEBcF1NPKY3U04n8YGmuo0/Z5a
m3IWVc9yqeQQBtgQVq4YXAFkgiA5pS7HYQj3i4Ru0artBRmbpaoUG/MrZs0qq2RDwVUiQugL4Eph
lP0kQXVzsJF7HyEuwGJ/rQfDMoezRTAE/NHuS/ANCKRo5ByBlvfZAx3Agv/LovncWPVWvGuySla7
bqaeUlp5kG+VYSvEAmWnQEhxZIpgtHPmT9NPzUAAwa8p+RqYlCbJgNDrT5COL28aC6sJJlQtSbdx
fCusnbw48/pXLlaWxHiGmnq2NyOQwaXX7Yd25vQDGeAYQpQp1wkEux8v3jizQVU1GpVF9Wm+rnYR
MhPdQaMqqFtjFFPAb33LN+KFMRCIBFv6P5iwLYBDNSHNHH473ybb389DfyZg8JxlV3ZcLV+gjzfi
lrwh6ucBIn6AFbob8D/QP4gpGaSLQxbe/57TykPOOGMubf7MIdWeLboPwBu6zhWkGkMJOJSaZz0a
qwW39xuyCw3c5X5uoCKB8Bdz7OoS6P4mGHh0RdQtCdF+boRBmaC9wIHeAGexg2u/7z0w+cepIZ4y
KexW0onoy2V+O34HUfNDvZsNYFj3/oM3A1xacNTkz/wVjDU0pT4//iO1+MHVYraxbjmuTESm71K6
BXSHkLtorXQS2Eyu/3MvGD5I4KrLhsVCFfJNl8jwaY003dNoJ4h9HNPbrMImtyGjScgyZHZN15EG
ZB9AiOZmB0vryQfPkCGe8NQ9W4vYl0r5VnMWyGDKFs0KNmI7+phLUSd7iguGU9DN8OFxnaj27rDk
fxyXASxhe3qufF46iV4J9iG0K6zWqVJEGfcx3IvAEm+JNCjbphOyiZqAeIpyFhMzjksl/fMWvBOp
rQ0MTFMREHaCRoWLODPRzBpS58ecseLYOBCgOkEqtNsU6gs6wuWTF6fEy57MlH59seDmyNs9cu15
9ohNTlLKZQBUkoM8RsNu+mCsqHdYGSM+ECMw+EgDJXVV4OiF0bcXMe9c8ehGk9u/jWtddL5vNr4e
P6gVyyWTc6z3gqlvGe/p0/1TkuBIi4dLhJRX2YV+Qb6ZQ3kMlTGaSeVQRIKEXEenfzrfARTma9oL
UCIXXcdBbZKw5pgZsaHkNSyx4D6ivzIpjut6dvFTr+8+MUKJHJNcq6RhuPiNloBAVR4PzJio6Oxj
y2AFx7mhc4p5soHOhjyGFFZC+vcwOyAmuQCoX2U4Ahg+X6qlXWAnmIZC2bvMPaTyhS5tIEMHF6r2
gH2T6AoZ/m0HuMcGsNC8EZ1wunQcSL6foJdz4FUK1lu8UgRouRz2CzhM9Z8T7JPHLQe5+us5n50u
KiH+1MxGbZrMiGwPZti72oVVPzcSRBUdO8iA+n8IUW0+vuj/hts7pFiooH5X5uLHhfNSfpXtOXG2
k1NA7GAdUaEpannNhBaxI4MizEEsi/DZ1bMhY+6cT96kiYgVBxPEsQs4WnyJn7hU/vdzHmQRcxnf
62HYZGDsam59Um9qKuOxS1qowdkdSVFuuoAUMQC4juBdE8WxozNQOBgXtVwZcDSfvAMWvvgqHaTt
/34swopx21MzGhJT2/d1I8nVfBUM7jmmjLTAoSywPYnlHz8OglpHbYdfCV59QgWKOAaIFh9Qy6Wv
v43t12rqQLS7P7hm8j6o66iXCV+ebjpYrrHa4MD6zz/L8eeDn8ThQ47DQxOW1LI0efXb2f0nmFwo
PZ7JWZ6A+JB+APDUjkZdaerZYazU+WQNvdDE0qxfV1W/cdEv0jyM/6XE7CiEer1jWcVbiFXCba1F
/1ihB+Wn5zxl3RGzQa+kPprBBzeVm70sbJztpKIkMN06r2x5qZFSzI4neO0Nddj9wypsYsjE2XO+
1OKpYlYR8RIToViOtlzXBoOSdK85dqhLEJxysddN6+x8BxYxTameWFClf2xYQEUqd7s+CFsYb6T7
owRUFRwSBvKrS9odV1gTafa8iPY4XrGRzktN/Rxpc2zvLdQk2F+nudXoTssb8RFb94MPaR0mHQpF
JBQOtwn2EE1puFdFxSMg2n/OG77txJgdNznPhDaIezOFcUK63dJfd1qnEa1Y5GH/Il08W85hQCAh
uksALbI585ce4QcjEqJ7M/DNqJIZGBl8H7U4iv/D/pjYfo3NltN66A7AhWOjGYmHiTP/TP0nVIPu
xLd80Y5EirQGf/ySMvpBQntpaBiGuR7d+uPZIVnLlJ7jsB7X/x7FTK62VGEO+d2DlftDdPforDwg
O+S6wBPlp6hNrq3zNd3+/ykp+gIzaZFCKmneV2SsMS6REr0GkOf7vHGSADvOa2z1SUS/Yhz2/fyc
1H8hSzN/Dp2dwYmB1aN0tORS34WDUCpAEnOe+1lCP9SpNZxoaJ39YYlyPP3CT17yZC8svMCItFrp
1FyMGLe25xZA7WaJPbhnYYeAf5uOYW7ZFBfJVBmmlascyUlsAX5qmaawdTauIFRDB4vA6kAnXkb7
SXi61pcAZhC/9MIDIurapR0MgR9rdhTU+zeCxh3m0ZJ3+KANrVK4ospcoztyOxy9n7UoIjX9i4Fg
14aob0zYeROmDmzQS72g+gKL9cJb/VS0ggwjU0WKG666ZDoQN3pUX0cwxBpsM6Afki9kSf8f3r5x
mFyFcEdcX+hFPuJZGsct2eWR2l2XWMzOUH39g6Szf5cZAvNVlNcK3sM2jhUmXYvZ1gOyO0jbAp2+
8lae6kF/0rnyaLzj1yM9ySOpqS3dhvQTJf2ALnatQXlMGeQp+feqKgsg5THsGZ5UiPd3uJyq8SvN
C6v4nP2calGSuJ04uHSCsNHn0ZMAr+cMy9IOZY6FFoUlwUBaZpjLUXgzSAPtdf/8hwvzxqtPVVOU
YHfkXN0u2exn7FyRAQujBEigkJy/K6/8yXNRIFdEULp12uFihNjUxZpkspNQCXvHvr9X1XlDB219
ATiHmzSC3YutqOvM74EiNZnojuW5XSIER1dnQE9Nfij1L/JJZBVkG/sNg3/Wpwh13tBEhsa11H+f
5U8yEDSuNiSo8hw1Fd9A8RT3YrUrqXeoqbM/hdh55LuBPzIr8NoRlo12Bk9ogYEMQTr8G9Go+jNV
2HOs8CiZFNPJ+jNGbLJxS6iGJtcBCb7MZoNe1GMkNCJYnqIODARhSliUy3vvHbqxVwsE55gtF1l4
b3v1TDRIjFFfmdJ1b+1TGH7S5OBkI6Wt+439lJPoVdAYAtVmSB8D05XRbMNDAT8BnMO01OFvPM+G
e74DIFYAzcAp2ukG9CZpj4CxMkLWB/14ndnUXy22wwIM7ams1I7tUsMG1qiN1auSBPLWKgKkVJgj
rzLVvk3jmLlj310M4AprAUbb18gWqfCNdHYIYR81YX+yHje2TWFWZxumKL3DyEYxQ1+u58uidkSy
pdyf5rvkp1dMZrmfbHYaBsTirWGItFOQeJq9vBjFp5wOlae9c7tC5gd/vLgZ8zAmRWmwNEU6IrtU
41MyePjL4MkEpfQvq9rUO7g1Pc5Yv2+g1Rb971jlcY5ekU7+P6cggQVb2aIqv/bZyKz/alPmtJnI
tSWowJR4uwXmJzurYsB0lM5OoCuffMMrGoG41xoJcIwfUa8Rlc4ELDspbAi9sqMixTH+DMb9bAyg
nQRrFJZ6pfm0bu4a/vy+lhq0vP8LpS6DcIGycV0Jg12XevhbxN5lONR3qf3nYbtrzGeHC+iU9wpA
eCmz85rB3GJa8FvrmlwEzvJkeFllrXSdW7SIMOusTL7FJ5xedVmbr69S7fcIQNuPYoL+1C9OXvb2
UkkDQD/66aj6aIB37srpCw1K/hXb2/QT8shUrlv0Npb6RL4pxNyKi5DCSg+anMATFL6ug0bJabDM
D4bHYk0GDcZdkgTRCf0t8g7pS6CAWuC+hPfXeKtuXct99FhuySIeAfAwOI4l2/DvtaQX+BcmGy4b
ZjrxNkWLP1GK5TLesS2cdDcRQXLXJyeZwvLpEMoqWWCBtvNietkmKqH+n6e9agQq4MXOD8gXbrgs
EBLRyqi5ES7Z2WMFtj87oMZQIcQsvaGh64PGTsZCzDG6/HFAF7Bv2oog/TFuzcbtZ+PMOICyULWX
4hNtWe9OzUzVeH5lhSbvHJEW7BtQSw6cFnvm7SfZl4vGN0TlwQ0MHEP2GIVwD0hHiWN3JJ1Z5rBS
SfXZcCksAL+HDDt9uPBvngUi72Awbf+14DSzEb649zlxZ1uJapBf4iWdJRSWWfe6QVmZExm5lW0a
8QdcyZ5x4FI7GzN/FkR4aWcqkk0A4MqSQYgCeKVVgt4kAaisu1ndAFU84en3xV5MBRT7ugapI2sk
doXQbNx1syqnN9l4k/Ca3h6VVC+OE/uhuN2CFp35drPX24852IutASkSvthFwK1Ts5zuBa7fdv3/
lpXseXNwunDQXhkRa0V9A6HurJCty6lesDfVgWrY4+nGKdpSuulEhDAg7MoWqUPFoFeSGXumLfh2
k40NJ56nR5Y6p0BcyO39jcDn+kztZLlCO54X2jV6OjFLtzNdkGQcpz0PFqJIQ+yl5jXm8w6JqeTD
XdJ8RDGPnb09JE/MMmdTPGbC6/qZ8CW+cSRArr6PIzUk1eBUUkRXYE3z+OBrmGOT/AUz75LT104u
uAZf2AT+cz7dPoHWiDfW1yVz2pLzhnfqzsbu8YiIL/MZgst0s3x6TBa/yjaqcDgdFIjamWcr7yuV
05qxvdbRPKObgUt/h0ZqiOKNrBpkwi5KCiI2LMtT4ZcWhzr/JLrIv8zKYls1MfYXTqSin0EuUcp4
gpLZrrwf+qPXyVR5R/p8OzD4MN+3MyvLolst4Xb5bPryPGi/3AikiXARHp2FrE3cvhyAXe4CwRPv
E5YM3wznm7816hC8ZkjYS1qJ+ph9wX30tbeQDntjglorlHvj/udjc4ibq8s7U2bR1VWCuqezcU6W
LvZAIc8LqeiaH07Mfx+3gKHS0e0NNlUvpCoLSjFj8UBWJ3dY82MQmP4LDAr6HNRt6GqyQz8Aqbef
tQMeWRy7os+CQ1AyF2Uq33fhIcIXfmMqcc6NPeD+0cZd0MGUcrfC282eOAjr9Y2SDDB8p+B2Wf3x
g58rWUSHHSrbCZnEnSwJ1pgUNFViuZaI5tTypThnyBwEn8+HgBxVtL+ltRXHE8g6/OUB0pYavzmt
Addze7wYPNlM3kRI9pPmzzI6hGtSbteZ9u0/gWRMUfOulUWtpP35bnt+gHZ6IAS+BOkRxwAnsUnM
tAktK7u7yxXMm7Q3G6zKmfNygfmZS/BGlGNbjoFVwWxwvoWh8T5fV9Y17bOIYEyhURrvaLzRjPUQ
VHdGyLSYLJ6SsxEREeKRmJsQWXbp4tBnfTP9QIp8f5efR6XwOmvpHbMcGlz42kVKHUInUci6JQdf
yOtd7IvQ0Ay5uTdlO+cwry0o1FqWNfJcWVt5u4EVM/cRRrQXGeAf2RPIjseC8b9YseYO0kTEv/d2
CW+KudmCqjMx3jeIcn3hbo+Jxr3rBqfsLo2CnprUa0eRR8JVkjTWow4QfwXKc2z2GkdeoMwkG3U8
GtCsOa3s5CUMnxUFFFcyizutAENopM5qgDNTAEYmJM61pD1cp6VT1ctZV0OMbDYzkBvu9aYqBXlr
nqKGwhd/v6UDslCbkbEGw8/ju7qVbJqXAkvxKP2LOwQxKVxY3n+biqa44FI84ij+sWLSJdBsfuaG
G6Ft5Yf89OTsmifjjvEN4g9U2TNvtlVkueXBM9a4tqKkpOd2y5F7PbGuQd+6akm6RFlirC9wBrJe
Gz58yCsv/JUMnr9m+UKNk0pa09LMMyhPgTCtbXMxYwbiTkzap/XaQw69++GevwhT6N+oJoflPFMm
DuK3hyFHWuZtTRG3bQzp8SbqTcrohFHnGpjBO66MISBqAazs6+mhh1Me9x+d1e2Jg6PeEs3Z401Y
B+/wnP7muDe+SzKeTCuny0Zn131esrt9AI7ohj8dOeGr2Qv20wwX+sVDZ0+2OmClzFxSZbqqiw9M
VxQSCMBaXPBk3p5YROro1XP2+24gzHX/9luU6hAfMEp99sQ3PMGbHvGEtqwFQPw0Cdo+afWIJByc
jlZg9gUd57zsFLqHaR8k9G80VXiwa9qrAkDXiMo4suKGv667FCllbO6S4VjmADBmEF1XovgFBX5S
Hr5Y/0f9tIiws6bb/3OVRhGR75tp1i4+kXBDf1//YWcBTa4XAVYt5ek3HXsci++x9qRHtvu181j6
AF+BkQADSolsWq+cjYEUOopDfLLHWfMiY+dypJsPQdrWQhH2fe4qzLk3g0CoA5YM+P7uibtpPC0o
pgdoc6tfxPlSSzSYu3bKmX+kkBDJ7ezTAK89dKdW4luQjDhew2vHwVX2U6VbHqPZrBEhxjghCH14
eUQQ0Yz1XyZgh5C7FfS3PzBmcYr9xseOM5LFYfMOQudBgHiQByH8QGNSrHcdgkjqynurHQIBnR+5
xp2+URjtfvO/6jEM9mcl7rwrBk9+u2h9LQgHsMuIeTpjwFVgZKDZImvHb9+ZMMHx+Llj8oTKQTcS
AaBihpKkAkVya82LXhvsrBLqj02zf+581Apyj3f/gGW1yIPbjtYQVyXGXmN6ouFonc3S+AIhIlz9
8vdQA0O1n6Acy/cFPrge7dIkVtYC0xE1RA6xI9WZ342IGILxlDOGVX72TJbm/lZzQO1tBg9YpST3
NnTpr5ViiZ1GRSI2tfITCPuMYfhaiZmE2EPihPDS773eFq0s/WSLQhCrw2MTNkapa+UxYTYbD54+
LQ4uFGjwY1msu7fUS0v0DT1whU/0cmZBBeLF3EDe9i9dQ2NPEF08SBzLuUTvWP9uZ94XcZ793YKp
jRdtwKWgk8kFv2npNtnNKaGJtft6O68ZRvAWWN4Dz9jmGsIFPDUKM2jyjkHtU9AdWPDNZFsdh7gK
KSeuT9HOH48Y7b+NbSYWZWrNsLzbwMiDcz5jDRh9HKJSBBpia2QC+Ascjs/5VFpne7KgAMdjCR7Q
oaOjXobgQYso1cfsbAFKVLBW2UQpleMe/+W43QmvIwjp0wBOzSHnW2KhB7mOwuU1BN9mPFd61Lyq
ymdDXkm83yH6aiQofiKYjB25r9FILeh9z9/lhVOpYbxThjmfYxOCy8LASRX1q81A2OSRLwtFATzS
rjKfYGzlULAPP3cRUwKQrsnTs6MGH7/zLg+DcBiCsvDy7BOZvMf9uORLKAZevmnYl9uusiG/2XJm
9rJYMazVLpL+ddtwVWaxvmPENsVfLi8ief2lBm8fQufjrwh3tRHjGe7NPVLb/65WEEJmuIuml/Dw
ZiHkNQWlTQ17OgPC79aKfCwAYSgmudggtlke5V1jJr7R3IQxYZiXrDB9wYGaQxo3UI8lt1qjsFGL
3XIg8KdNQntjQbbY5fCG1Xdkh4V5lkWbhbCADpYY1yOXV43e/r198f9avYKd0NE39dB1C/srCuNO
8oQeuaxTVp+HhNkjQyNEwNYIxqs30H5bFXZZ/DsOGDFAJJIUQPVtGyginfwKdsyMiL2WvvlnlbT/
DEQLXW8IQ6t2e3ThTLG/fpPb+3RMhnCqKTgXcE+zT02K+18lKfJREovJws7+jbU+ZvCOjLji2WKq
zuTFNhYOnKKX2kDlEQEvRwGFCCgZG4IsC3nfiWnBEVriNuXZWfax9y7mpPCKeMtKo4q2D03A+dj/
20UEOL0F34OZ8tFENBhFNHYbwokT8Fvg6XoAPgSY2QDkkC9VLahijluSk5Y5vh8nhnQtdtximgtl
7io7CaLosgYAWMRiP1nos8HqeVN8vke7iKfdK3Q3nVJxP4mwMsMXjWW5tcT6ZsSIvYY0NDsfwiCF
3/pDID4gH3DRWGm4MFL4de31u4WuxKQB7dckOU7Gk5ngYtQ0MJGysiiBiIcVEV/DlXq6NZTfJdW8
WyKIm+x4p1B7/g==
`protect end_protected
