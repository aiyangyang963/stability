-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TJevO5uyoq5mKuSjaVGAqlryWQJ/xCW6Qnk3DyHBK0OU8mQMrZuVxFZCiblGj/qMtdQdeq62jg3g
2H+JBtAvFGtISHJXGt3hOqp8zlbxOV3hL33I6VpGWJHWM3m/qGX+Eer36bg5lbpEC+anUXzI7KaY
CykTUSjHh4AoTSHMXiVWCGKnQGLhjxQGUsKhkRFXxcXqUQSOMNaTdE5Guifdk7WCJWBbwgC5NvPq
18weo4AD4gApJMcJ8iRyy1iLUex25p7oztzDkI0hNRcwAeFDRuagsYtK1susECSpyfD7/z285UAw
2XWo6Qpro9epDDWcnr/haN0VrzNTADWxuJ0AUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
E1GKuyPBgZulC00DxpJwigDhSBSZIKwyDIqO9csFuXfWJbCy7r8fN5/PykOUEZMEcK9pNTGCVFa/
DK6c3tNhGe29TXEdBaz5QXN6ImQe30BYKf7KNVx/aQJhv50B/FTRUXRdMa2V+LxeCuH6q1nVWu8e
QRZ27jDi/CCELvfMZ72g6i03IEfMEbYoakKGNY00MLaKiVkfhH6cN0pXn+tzzEB9Bx4CG4O0PCAL
mEKuXA7SH1uYuUbx+rTAp35eCC/C5eO0o5mcdM2orcECdDCFZf0hPnzkzt2xfbT2TitKlnZ5vuAC
Cuj0nXFlL4JnfiW4pMxOPSAVylhuB/TQscymKz5SM0uDXlXheW13glkxVHlHReGhxjX4O9J8+yw0
yvfHdYs33BGdrAzJyA1iA4WwJ89/3USZkrR9RxvaBJ8C3aDqA0aZ4FcG8i+rjAdDkT4H9sdGY8Be
qcFKR53hPnASsWsJ+sw+gPwNBeYz5Lu1SVJuKLNzYUt4FghSZ02uBvCqJKcFO5QKcyqBAuEaaaei
quX3PumjXqljCW0ip++R6WeAGMT2KQxKy/UZmOUvjcDoe6n2x9pl4sdXbAJsYNt70k6jBHmQ1oSo
McGlPKdnFgXh3/N6TmXogdiB8eiA+MhaOLnUFRzBDkXY0V6C4sxJqiq5q26K5Toa7AJCVngBjhdf
84KdMar8VSHKna5AIuZcw/7ByxPYJlB/jZoMDh7abdshI16MhDwSUVCzEFuT3DvZRi1dOqgbSdOz
OvAuZCcDq68wqpiR+u/d5lP213h/gv7XaBZ/mEvYoAf6ak6AAXeIAdtSuN7KnFFC2CUETQgTgLAo
Ov9rilMxf6HR6ANzG5dYRJ0EqKGSC2ybUdO5rloRynHzlL2XGROxGmInKwHx9GpSsuc/SXJBXTNf
qck0NclvAhZY0zyY+S2EF4SL50FSerVpCtcMS4J7EhZdCD4Ua174ZPjTXT5n/XhPa8fgqdwkBmFn
BMFLB/Ic6l89lY0mCxNbAXdBQjaF5AJEwsmjtEpRUb2K24brQ6vrORzvo5qISj2Sldk1XX85z2Tn
WOQfaqNOBz2UBLEpegVGDb2HO5RlX+xCHK37+/dpcE1ImkbugYpP/3cPqr1zbe6HocAyjDrq87KJ
zaO3mylCSWDZstfWN4kNPmcJqjQbhIJGO5SghLb1FY0J7fuX65KvFyxlCRd1mcycDGkqhm4dlmgf
VCVuOJthcMWRq2GNBzjwn+7NJ5VUSM3tDtG5vOMwKOSZZd5ql4fh5N5FTnSERlNULLdjU6dWd0Rv
Gu8rZeH6UwmO2f3u2lmBuft24XA31mPF/Ve17rk18oYWD/sYj/v7z3HQXWB72dVC/kn5tBeQMcON
fBE4ygVXhy/IlBnrRU7mt1N0gA5zAVBMaPRcek/Wm5ihlzyFg7mmsm0B6ntkmIt1rnJ2/qRM3ejO
2WaOC2rtDiwePfQftZ94E7ZYSh7MB95BqUFO7k1rI0F8fDfUNiETkJMlQEclMg6W169GGBzSbmJQ
hP7K3Yo4jmcmH9QGKeFllV0ybv+lpLshOO8kLSkR9IKPKT2GAGOo3tfXluM1XDoP53zRI/KMjWXE
ImQ77cTenJXQZbC52VBfItD+qa/58HMeqwnin6DlEdzFCkeCLapaTwyVyAHFjg3ycpO0M/uBpejB
1D6MxMYnD8syPRikWW3UjE8r7mDRbd+mb+0qrWHfUfK2kmGOYs1gH8jyP6uOH5WdWmpmA/Xaw6uk
KsZMLnzNymmtjD/x6hDSZypRTt6jTzlcmUyYOeg/xzZBIOm/E4tlbVia2y7SNCVKIZSsq+cr55LL
7A2VnLRdbHvwvLR+eXFm8a9z8TdYKHk/wn3JFrDYlgUSjBo+CwZlLpoh1kbWxCRTglhXGaHMYQ/j
qKYcrMObssVEH4GBAmB6yTl+xS4vjhXMOV884tR/+rcmwIwwgIFi7tjH8U/+QzLtGDg4Y2EDqpyW
d8DLkDhtQPGc/PzuZfBIuSIiAmLAxAknyXvWQl1ipWyKPDxYg/JqEpKzbKiLZIQlzAh05Hjfg1wA
0TcXKm7yjEckPrBIha+VrsW2hdLATnxT+erqhju3f/6uvJu66i5z9M9wKdNqiG4t+DVwNbDjDkgo
mal9Wqu7hmLG2uCWxptXfdPnLg0CCohfWNB9bgGJG0bk6eZjrk/7D3vY2rMKjar+aCTCU9q2na2Z
/QlBnYxr9l1W/M6slrGqk6fyB7IxUvZYxJ0K04buVIPvBMjPbPEqx4IsCJUeHVIzf3xZZInpwf2x
GXguLG0i4BGweiONJSI7LZc3Sq2dzhke/r1keMrjF8LBSljlJydMnFuAN6yWj6faCc59Sptmmvqj
NFV55nucGVuw4WPUTmDOJ0D4P5nFTExsu81KVjB8eBoRWzoEXdio4rpP0UH6ew9NHAdc6xr0V0ak
z4IVVgClthqnFQ9B/rSmsrUq22RrQplp/88M6T0UzL9ht8qVxJA34DEOou6KLSnEdFsaJbVAvrbk
zlZlk26bUmIIKg091YjiHzr7ZIWpu67XJnNTPQi4axDbZ65fiOo6iR0j8dQErCZp2+izJRiJjpIH
HyUDuNGCduxf/k0jSdhgGGXQVRQchOwYF2JU2kmpDKKdG1o0AHqmomHsy01MXd31spzR9lePm+Ff
MWKwO2oZXtFIdqXwFecf7RtMjJIu5sA4ff3+tVm2d/7PGWkmw2406mUNJH0k5qPmQOVgEY4+Xrny
pjDeWBPNIo/qjs8WzXhi+zMp0M8zkvrJGsGwu4CVWKcOhP7Z2r9u+CKIxbYWyWp2ZzmLFKje2djm
GjRdzeO+BzUt9rvcVAAaVaVLwKDExInMtLt1NyRHPryJsgEwPWI/LLDCF6KqT73WejfwAR58yuu3
Qv8Pl5LvPgRv/EDzjeeMl1ivlgcvUilg3n7Et/6yn5wfTQNf/a2Xiv4AWYN8/gvXP5OftJ9dQTnD
75uOAoEwp0WPLyjGCUT9NDegPKtm5wHLset+hhEtwBTEZFDNRf7PPQzRx7+paPL+l177kqsXB1BI
6x9cjU4AP/cKPBNbcbQprWyodYJaRzO0oluXsCrlxA7VX4jwTppsdQ5Qa5RiZ6bjR2bO/DILgfFf
s1Evmp8HH2k5zAJmbOQYha2WHs91DGmfh0ouemQrPdbvrOV8/7jhYi6yrG4vvbCfgCCx5HuqcfL2
6flBGYm9QniAj4n9KB2/RmpwlVh5wvkPyabdlMTMrPTnVMWxgWmqP/FRMXtqUXDuzKKl7gX+O2cQ
R3z6e+pwY7GMGuFfHo1TFOHosk8c8w/ouKyUfYyyP7+JOMawSuyrFVxYRg8F+WbFvLhNbDJ1MX8Z
sLY8QWJFXoT4xVe2pZ/e+DPDNJkzGwesnNk08DtQoIU2d9udEXdHVGPhGpn8T3Dn5+dY/SjLQKvw
gAm/IatvgCHNPdTX+dKe0jltU0iW2toRBbEAj77L2X2soTI7Npq/KPNsEcYY8C+Frf50PukKEU1m
iDp+BRxEdfic/+RpMHjQ6r5wTGpy+kmyp6N22C9mJ9g5XOXmWKjRQObX0jlVMyLEeFi3jihqY//0
EBi9iTOvjjqjdEs+Tfr8GmpkQUD90Vyfb0uLmGf014CCTBBkWIzygKvOX+NMsHue/dm/iTEtHpzy
xWgtZeQAu4Mlby9O/E8EbqUYnDxqC90IlPWxkMFnmgVFsqO2pmNm8pbUpfYULiFQP+Yb5QshxnSl
zbrXMNvnCJ9Khr1+DlzqEF7aSJMiDMMF+hoPSUdsz9P482e4cIEgM/s8os5Yh3sgu4PPiVNtzBwa
6uQMtxuMD/ueSaSEfLMmn87wk0LpZfP4ERfRmMscWUGNPQATOamJ3AnqFlgidGA8dxFKgb3hJaEi
W3XK5pKkrWNqhW+DfO7xN0r5W5wqPAc3h2D+fo0sCOnX4pVsG9y2ayiP+xhqbZlYxlSbwy2Gfie5
aRF+UgVpFbe03YOlIoeKfTTRAAJ+UCo9ErcbdiUkXg4aiCXQHaAMQMzqamcwy91aGH7+3goGOhGt
oHPXl92kozW3tjmP1iYphAAbJWCIkL+BUd9c9Rposz3PmDkIx6CKvkoORH0qjBv8o2u+2GEffM3d
uKWIeoQPZM1Whlw5nW09wUGsRqX8hxsWPt3KSFA4pQ29WGfcArnJzDSORRyrwnVk+43/IQAjss/e
ZP18Jmsd3KzIyJUbmhNRKlqyBfRTtCFJpD3uVCEasdhFuwcB3ui2lhNVNJVFfbjbok634nkXSa47
hHtefTw+QMAjgEiYYMn2c5Ytz4c+bNQUEFkwt3B5242IFIP2maivFu5Fvks6gzmrRZdFY4nZ5TVx
2iW2Xw5Suo5DGxLVSZn9C8oAAx1+SzjKsQW8IeC/NgIrxryRBcaJkRK+NMvTRlaGkuw8RN1f6VMX
U+vzSVntSJqaD2smD60JMVWLvkVDgI8is7+Qy/acvRMcUpOwx7NG116wygb0ySeCh2xOjZFMPO37
EnofnOaihKhPS9LkzbhtDXPB7bH9PnjjsjMPDXYhk4e/XuytdVyHrJnTYASzlyOrQ8Xjw3Cpa6SU
3LmPq0yqmm41HziqjIObj4eH6jyoOpdfEWUZziAFWlVvIoeshscn7DRRqmb1UREfdnnj/S6c1apw
JrgMfJ4IcUGhFQkrum/R3A3Wxs4hXRcQgitMn86CGyTKitkLo5sRFae/TOzDomd3DLey3Na8d3Dq
58+wMkXrsW55WGkaFCleTYXa6exEBHNJt8gGSrbZePJsNqCcaBsnbPMV1CtDcWgsjQErjrCwrSl6
6Jp29XAGcvRYnTOA4VGzgHz9ZDCj2yKORrFGuJWh6ir2oqwJ5T7pPCxGK48+r2FYouF1oBF2/mRs
LkxZk0YoKWXHSgeFO9+9hPCrgpbgRM0uyuv6IWbF3CUdi+DIeWsJ2BLB2MxF7EcxRF8C1fez/sp2
RPtIh4uVCnsi858hbN9dy6MzoAN4EeqZvrCSK3M4pzQ/0Y/HYsJjXt8O9yWIuHA29eQDwTpxviQG
D7qA8hgK8jIeF054XfzhL1Vb/Z74FLgnSdEctdKt06BvGRdhp0OEHE1mfDB2fm7t5IGw1QhVdYbM
pA8t82WV7YlleD6wZ2tKU1+AIQuxdgCw8agueKdT1SM0HFqdOeGHry/WSpupkht++LwT8Kang2yS
p+lzRSmIU32YIIGhiubNhYYta0TVV3+sKcsbxaRmejVQ1UNH0WpSsk2FProUiZWd0dO9FtYkZRSO
O9Nq5CaQl6CM0muzhnBSYHqWw/UNgiVPIYzgUXzeNG+Wyu1wqJqqu9ENsSLqst7oiwpNZi6D+u3v
qVxVJBTFWcmYpddSlXnLsl2/CxVDLkRRXv5mP052OqLSySH43gnexFNKEUK5GvTyAEIci/TgMY4h
mOgkUAZYoewd1wsDOFzJiEUq45sqliSZbR0iAQpKD3Yz/skG6wKOpYEkfwKdOKWSrJ7LcDAlGcew
8gPg6eWNp3MufLvZiWET7Oft0UFm0G2GZNq0YaCDL8lGro26DyQPGvwEDBwHSCRGs8ZtuUp+U8/w
Qxsh42b4mNl26uLJUgrLCZEDfGqbGX+SXfJXHbBwa3maAtDJS/Qzu8lcjL5H0K5cl0SqhhI8iogv
kMQ0e8EQzH0bsEpUFSNT2bJurgZQm9+AAe4uwDaY0v4YvK8jDRYUUtEclVp69+/2dcNyG5r8zPNT
VOIRe2qUzxmV00lmcPDCVCkbRGWvF5eSOgbyj/wgHb8nnvrfG7gdcAVnXVFwX5skRXK7zLRV0qMX
uoa8goUOLFSk/Zs/ZF+DXNCB8+OQxQuSfJJebbqCbP0HBXMelHpI1EkcamBQPa1KFUQvKJDxoutg
jPX4pto7WasRhfwDhcTm+D3gbRUsqRBFyGK2V6fqbiTVcLRxx0A/Qq6pT2txPREWl3FBOEQm/1ao
qY8PqzjSSxL1XmdYvqzMjOHLep3Dp6Tz6UeS9Qu4TG9JbTyolmlC2soBRk8egfg/8hp0LKsXNH2f
rxgel4m9Xr1aYU2fsYk2y8qlIDSozenBKFAduvNKZG3tWerv3p9GofE6Y4ovo0x39H/nW7AiHsBg
nVRmuHNaC56/6LlTS2gBGlWAdnI6rydzTcmux1Rx3uIvSOkQKI9TzGIPQvCzFx4lquaMIIWWdxET
NkAk0xmWSjGhQ1fdCbxAEQtvjVliOBI9MHZNLLhCCv9XJ7O/CHatejTB42/oRw3+NsgRuJ4gDeB1
CPF9PTRfanJTXxtFaSqQZWi/cH3+Lct8Bc4k7Ip9F+UHj1T58UKKUA/iz8T8BZpblAfGOYsZTx2q
Apnh40vBb0pL8gZiBPZwE2Xu//aT0D9Hf0A8km7e74EWm7GrkfU0hWryxVNV5eiAkW7OGmSdaNzv
BQubWOrF5ppmp4q+G4jzoXUtpUPTuPySI1EuSC1mZLdZq5AEVDLLCVFNIsPVxnlhTomsm2isflTG
qDOzATZAm/VfGhmV9T06CIzcsagfCkZKiyD6W6XqVZjQQovPJiuSDXKw+OCTf1GmuXqC43EWfAle
BrRkF/dbAtw4UqrxL9us9JEtuMdzfn1ZKAMKRxcYgi+m/QpAvYTyEYdGs7Uv5J5rw+iJwuxmBNtS
9+pis8Aw+C/S+G7MbEXPd9XYrfkbEJmn1gECiIHdVmnom7Q5cUvFzv2fu8JEuJWfL7ftf+qOrprJ
BSLBNHgwKxo3Ib0IyrmIPz19l2tBpSmBhVht+Ynr+UuH/RjovvgaJtpPURlPXgdZtY7UOs6aUXas
w/pa3jGOuP58AmZq287wEmeiKY9wDwJR4eUHB0MmRTtGqXXG/4BsNIflKmsU/6yEYX26T5FJ5YkU
Q/06APENR6HsbNJJvyk2fR7Lhi6zjnWjg+oMZLT9QMIlCpKknw01x4clTM7pBERcd90OLXlPvZ5f
zvEpMJwyesMdpm7QaUJem11fAUENygGWUkM/nybsBlULf3k+lGxpmY33WVGEy/gLlVBgn8c6LTul
U35mgim+BuVAwZLsI7DKK/vPBoabfIhWFgtMdwrSlQPbUj7F2akDj4iRFH0zxJ2nm6wkrOlz/Y96
t5eHACjiPdmMWNzx87Wlk9SNCVIWMSSlc8HstXVQmsYbNfOYFbAHS8Ch0ueNL2ZPf+Q1LO6pJ98X
cJMpzh8L5Z4TBkNXqejG/36897dEi6qsQxus+xhCby5FfbQJDyRitwAgY4D2e46T/p4c6PhRuhhU
Ylhw+r549diVlHfL2QFxuYUo/g3v6loag7CNssYAhD0foQia5LqXoKIahpc7VAxkwxkKcJTC8dj2
TdXrSNWA801hoaz1rPysAyopLx5o+ToPSRMJnZjMuqRjnMCeAaQZDlP9D0hyVV0o9taYKaa99HqN
tInSsibRgXKouQtQA3y9GRKRq9OMNYC9emUYcR/GPPABjOvPZXjN2A1SQ182OVuH4BTOeLGiqJTo
kDXBL39/vdaRQmpXM22vMlCD9JF655l8s/P5qb1G1HdoqEOihKN+o4kV4aC9pV4kfk2mECMdhFAP
dj4yi6uJP3/H+qsamBSRqQNxKg8NQ1N9Ndk3wyO+Y0UTjkGfSJPiSqI1A49cyFuKLI29yeaLHAL/
3ZqNVbvcyyVNJ+GnJ/H8q0f2wrgIEwZOOPyD29vzjBvBc/p+gUEG4Np6cbfQR+kfARGG8OdalMmp
7aLKiPiG81ETKLmFzq7Vh9VaiEu1afhvOMWYXrG7ngeirOcN3dCRZ5K9fBmKr83hcNUatlsCiz86
9RiDaSRkO/C/HJSsMQbcwP6NsGgdIoxXzGm1xcgIRt6DVHKVvSMxK1LEFtMcaAX0rA1wR03AMWRG
TpDe2sSItaudOnhjzqp5i2uFB5W8YOQGl2e4F0PB8HuHRIGzlinKBocCcxWV3k63VpbH1zY5wV7E
OkZfhidbm/a4VPBPIa7Q79lCyRBAqKwZA5dX8zqL5+deorDS01j1EDyZo6gibSJIACTn+UNCbvJB
7FYo2vEeEiFWQNKor41AJMv93MCt9TPlp0bzxGO/7mEwEqJup6GJQ1h+mJMozOEOjrodoI1JY0ZE
0tMcd5zI0QdwJL1XnWCaSXIC8AZOfWQOVjw70UiKt7wDTZOiC3fe0sczP0USzLiHvDwNPvm6HfWr
LI5taWUslFFE6wmphdWaa1eXuoXzbENTnDyb0RnLBejrXWKLdG8pDA0jc/WWNRYGFBLQGfDWTDO4
XVuHxUQeReIVmDl19ze/HJ6HC3C1AAFb8MPBdvXQsND98RmNmf3MKK7Wm+/yuB2TQpN5q7EMBU+N
w1OLjbf3DrOddWaV6e2EaDsTCaWTrSf799LqORthy/oNYy0MJ/wpY7x5I9d9JgyjNhpdWQif4IPU
e03AgJ2ioa1d2nv/dhw8UyKj0gNrjZusycjFJPA0FeSsiBd6RUTS+Vy9NcT+slZQjbCWyPk3MTKH
6f26BwHBn/mDQFP5N6qZat7Zlb5VbYYjbsAaU/fQ7zZisS3zMj+YFO57APaYm39HpzRiMN1N8gSb
v42qchiNV/evvxsOt0GW8ESe9IanBa0RxgAx/fv7UDDLW/iAA6Emi/28D8kOwpYoJfxxJ0Nt1YYq
lUJWPph/ouujb4EQxEFuBty4P0aPy1/gp+ZYo6DImJM0s9DHMSMA3uAqO+AmSfEtpPAtGjSoGxIZ
jmxM7PiVVw4IHBaFGW2isglsE7OV5QwR1vTtTE6Pod+RdX6qNF6XjNljkNSFkmt08FRshg9CxSuI
8lvlwfZpUZ1UJam5nb395ysGfBFSRre/maW6mXiw/e0YE4/rhfknEyef7Nr06nc6X7HH3qghe2nk
i4WvsoIOjT616je/ZbLzr44FCloY7yZ0/6sTVdZ300bXFDBcqm7BQqVV2sZW1O8pVLTKHofYjUND
HVAd2Vz63R2YC9X/X3YqCeTxpuRmKs58aoN/ww8V3tY3jL1kb+3GGCyCliKOugCHpt9YSkqPp9mZ
u4qxIqpMDR9FN5oFlKdy3VS24VRl4kfGNUoy7usWJVO2w6XPJoKiP2lDuJ9dK6BoKA7TFa+M21zi
6va6UxUlhfoZT7BKHSnm006Wwr/ODRwbrn6tbq98ldYlZL6eyegAOs/M5QOiZDjpctfp9AmIYdJk
sr6yA9y57QNgSHLPfnv10yDqKPfTJWH76IVYjPrUIL+SlpBG7M8KDwF3f+v7XOSA9EeK4BheG3rX
DFaEKqaY9PclfRki/4Ijyjdwj/SqZ3vQ+c+7tmS3PX9ISLzLCx7E8mlefZ5zVy41Kbsd/uYpt8UP
C+4XGRUYuertojjyCYVErP0mkRCxSjxdBmMEPPx+0gJWuBc/nioSH2MP4mv++YDtcyWxFNU3i0pL
vU8qkn8/8YfMY2UEUvauaJZUrwrs7VLZr3iZUxuudmtEFDupQfAVlEFbGQq20jFuLnHEX6k3ntP+
IcCCA6+0cj2yr9HguhbJgCmkDwlrNi4wstqXJMfaX8psvguNCsUkqSd7V1W5tPPzBK3PFo0cZAB2
HkniD74IcGHfMr4v0zZlQ72OdXdMVX33XBKaZvXGvKaPR35gSm6TyNyL0XKrqQ6kme+uR4e7FECN
wymjNpMo8R80LLIHWO8UJfFfH9d0LLxBnv48akOUjNjZlEqgOO4TS6G8LSTO04Vhcvqy7enApB9L
Mcd85jn22BP9GNoVzLq8q2FNFUnR2/Qs6bY4H6aE8GKoyv7npxbmyRgDbp02xtuWKb2sGMCGI3Jg
jq4qYSfrhFp5doKg95oqqMyPW0orJB8HJa5r56WRZiNDccd5ngpeTSXLZSSq72FtvMTrAhuA0JVV
WQYS9qkatBs9vrIXEjX9sbeALa24rlpHBL53m3OltypQvVCN80mtSEGcECigcZtEyH0olK6iIKQW
WTc7E/FepNd0R9wxhse6M1RcqHhC2xHK7znXKpcT6rzywxhFRfj9y3eu1eW+/r+EAqRg6Msow8cG
gHOzTAOeI3YGZvMPXY3qv8IS7a1+TTQYE4qlbMBkKA80YGxBvjz594AhcOAgD0BobjR116Re1qnU
87ttJrjyG9WPj/WM1V+rTQ8vOuIZTuxqlNTNm8+xDquQMgPdQu5ISYtnTE/XajEVFYepsooPE4ak
GZ0s/CfldD4oqV5mJ9ZccxSE2JAsprsJXYbCiC0I3uMXUZUyA1MGRDcMNaN4Jf++xrKqArlth75w
9VKr05km4q1bk7CWTEVJgTs2hDaHa6pqOMS/ttBPzyUS7HNm1yL57OlPZH+4f0x8ZpChmSXK4sEM
SSpLutJCFviP2dXkX5u45X3jXN96bk+3XRYAHzagqd1dgJ5lwv1u882BtXVV2zWyMbjS4xJ6+ICz
KGPTkNBE1TIOSTs0h4KaA3B3efXAG3lR8zkWg/ztppDfzEfQNe5lsz1j0eLw66uzL1012+NaBwdL
9BGe73afm6ROmmR3rmnpfjbhjyNVl93KwzVROIn5/tVZ7nVdtCiwc7yF14RdE2C4pahoc382m5b9
l9e7MroqmOntuWNQ+UYi0ztxnQ4W4u/SSobFJMQGO09gViR6258w3qg0HF9iWRXZj5Drk3ILmGLs
TYlNscvPUXnqXOzOSK5YZj1DVZe9evlphfHECCUIdnaHS2P3XA1t2Qx1xa9akC/IJ9HuXZocbzRv
aZLe8yyhk4Pse4dFjJnXASMXNPOwTtkji/LtmGQe/RBMBr/PrI81Pw55XaicuaGm6yxi+mruGAFJ
kynBs/LQIg1YzeIRgeSZ2dzLltWm7hhqLjZ0LnK9t1naU9/FB/0ZmjHf3mCv0MyKEniepUEP+pIr
7JGWrzV3uYFi2cCr/nu2lJPb6V3uOgqpvUTM0efMdg5ZbSRhfpn0aTBmG6iIQYj97YnoRGOId14a
xTYwxh9rxg11UueHyIf8mkDNSRYpgt3M5QH3nQaeYA8u/YHQgtuUT/K1Q+FtDjN1EDBl4RqoJ4oT
0W8Gfj+zG5CNjai2NmR+0cUQ5BdN4Rlpnmm9wLP2rLNr/71xT91jiN/VFIn1+dK8n6YIpimwfGAg
csj2gn2+OUcVpD6oQRmV3YhgAllbwEceD6/hblMuagB4+NInaWjrsWfmosr4upT0GIvdHaHd2kpJ
AOsj+rqGTUpd0e024nJOrUYhT2G8qZInrtMBpFdCno4J5gSs9/uC/igHH6BJAoMKogQfgZfJa7Gu
TX+HhshLeNGTH2SbBFs41e81TGUQzXth/s15qyimgYvBMGq0UJdUaEQrPZnTvFF71lif/VtKWxKK
sjItYGg7hVuxq8cclfyZHPEz1h0Ia5z0FT2mmrX1mi65pPRu7SxefG2ocxMm/SxFusOSIT+zpUvz
XJLyZW8dsfIfmhlZB92xPL1eAGIA/ZQ1ZMYJips3hoLWbOapAkG5wU1kVxzP6IRKxebIFn2HMXYI
Idhv2yetl7BoqY/XHXOnhzxBeKEinvzFsbnziX9/UsFK2M9uuFuOSwLWTLKSkCqHfjRbGr5Qe7Ml
VoX0hBaj4tBmYNhNEx5tju0KvyBWl11vYKHYCd9SoIoPIPxCuGiZcdhZlaLXMKiBfyiZ4O0IVBRb
Jd2pFtj9eARgXaOOTnzdXoJ/HWNEEOo4KnE5Vb14sDov1M8wYfz7ZxQg3xx/eqWJ4etLIp15i+Nl
4iex9Ctr5gXTEDTlKAwasEQOpSWw/gEssRB+giSN6ys0FIk6hYjR0KGIXX4a3l/uCd1vyoDwHdaa
kOjFAALHRkW5S0iwkjAcBojcF5zjguM4pWmZDoxyH7d/nnI7vnBZueGGjHDdmxiHx/u9NDbFS78v
Bc09TI70Hx+HURyJ23dDTZMFQXNiglA26AZfRf134EBI+Wp89P7H376bqoAbEMDF1kinbDj01PVY
w8JxEyb0g6br47ojvMbhFg3zUG0892iwAQQjYK3NRztjn1b3ikAjizce1taAEsuCwH3tteNU5WQC
ScwLV7W8st8Teg8kljm7V9NfivQifBdL/ULVUIYXk0kQiWHT9zfgiPYdR4Xdc/GxIbeXxgl/484t
aCTkHt/jp7XWTQINGHrSYUqLUwDyrmnu6K4OpAWqEWy5nshtKH5UV2JwaObHwXWVUTR6hu0xdcEf
3sk/BH73faknj4ieU2dmBLDnjjmh0Mfy5SxKFMNfSJbxbpcCveWrkGfRBDO5seZFPSrNBKDilpp3
TP4SaHkQsm34coDfJlILdI+pvoAljtyftnCFVqZRY7fFYmCCtFDiIf7PshpRHrOa6rUKJESEiDzS
dQqCC4xNOJGgRGWxrmVVRtsb2pVXAAqX+lXGeiA14qkV9vajgFZ7lZZY5YgOn6WymiX6Bjm+RL6t
HOi6RNOOzYPLA23RG3ibc2e2fK22SVjnUFUjxT/BIm1vZ8VxRPHl+LmD4Dp2m2m0Z8SBWon7ELxR
y6LgXGHO1Su29yTI+fggAgwXvNUZArC8DPAgRYrYN7ZpCbV5Y/cjASTxxyfPqo6e69WOZ9DGSZJO
9YV7a8x5F0R2B25GoJ5ji3NSI5bF1BAaEOsvWZbmaUBU6ygMZfYH/N1+C09wGVi9YkIk/FGCdfaF
RK76T6mD191Z6qIHoKGOlRPuDDXBMN5aY3tX0vyk0affctoz/q2mZ7ZP0NCMzB1oaCRT/LrtD8kp
EyXo3KMDKEgckC0AXwF2hBRdkwY/OVLGbUvEQPJQnmxeFLRlIAK7Ax+Pmb5VtKBjaXYZxisy3U/O
pBy4ZARDpLIXPvANtadZwldLNEJNTJw7vsDbIQCoAnVKE7fuN+JPFAR/C02Wu7wi4DqbwJEIlUeM
+YDmoyzNqKS4HcnuTjNd4qh0hbzVRK4TVypDRGXv024eBX/WtptCaqyV7FkL4mcyJyfJVEgmNEUS
LTNvPC7UvXSE2YNCswECmbHYxV4Gztfj6CkUZCqskqGte7QtsWcgCgbO93CFRk8sJsR3Yu29LYEs
O57AUmCVYjMlhlXtZRt3zgQptOSDXRMYiB5H15RjtHRG7QqsvZNT4KhStDrJyjcD2JCVINb0zw36
//Xu3YjLIFwi5Egae3cK1uJg5plYLATucMA0yaw4nGt/NEPRSTGcYAmcmYMeKup6X8DUY4da0t4Q
FFwdmUxzrQBSva57Fy4Hn+OOY55Z34eyK3oqaDJLy8mKo7qzWBOEVV+S3f2d0mxF/mrNh97JoFLG
mbAYWklRNIG4PzGZlrvcMtshga6gLYNAEacuQq4LEyciXUEyLu/sctI8nh+QZpK02TT5Wh9qVm5C
siCJKu/xhH+ZBu6zgg1FbQAu3D/NZDTHei8mMX/ZNDf+nQqi52pukyUiN+MxjRONTotlN3CRiBe4
G40buJQSti6mlyG6XpdOtfVF21+Ccy7zIoxUiYalDMcjTIKC3MbNu9LD/+2lUXJMpMUSaTqgNvm4
z5EQi7d7A2Na6ombRozAK2pwG4vc7JcgN9zp8RxzRpBSGS/REOmcwJtEoI2eqp5+m519/s7z7yK/
JCF0LIlNepPO+b4Qi+CzS998r4HcqUOZdibaKbO3YVxnNozgl+eUWqX2aXXqcgnupaBQIcnmJV/Q
TQQ8o9Ftn8CSF/Kh4QSXMC/tkqiu6I0u4hJ1wMDuwKnlJW0r6o0hKb7rG7tOdOutJAzhDf0gQd1P
TA0f+dJuz5lhtbpnIbRssiraFCNvok0mOK488i6WMan+d52l4DdA/qiMaqJdz60ce/ZGqAqLXaEo
m0Uog4lPjl+s6nUeKMjIyYguxYIeONQRUuxwBo+4u6uet5NSE1d/M5AB9uICjHzAHOv3salEj8nj
bEVbWB8xJaRxwYSCC2r6+myT2aDHbHb1WGQ6TUn5zb+ekIjksisbmYnPqdmnonumnSYOh3OgCaiH
mi4mog+bx6swOSiAuGWVq4C6+lI+hChPF5eHGWIjCTQ6uICacRqqslJqnsKGSRMajZCCKybOy+8G
P0/9mpMAO0EezLpzLHIkuPbjBjJMgoNdBCCNniM4Oqyssjwke8IQd8iweQV31zmNFUNzNwcgL1SE
CMVK14vwQjNCjYHSovyqpsiKqRbVQ0DxmtCY08yfGfgUdRXgJsalqNt7AITwbgcw4o7uwHPlgNw7
PJnU80rm551dwIpXHak8zX3Oe+JwIuCinvELJLewmJvXgjb+1PPwdT2PRApG/Lmlukqc1fZyM7DV
cuQ6Rqn09GqiRPPj6kNnLyyQQg9p347pFultvhBzPyDThQd5SlHyol0Ad/+hvDK7P2OJAkgAlnfO
o/U9aNs6IjQ2DjKYhC54YI/NlHP2ju8hpg8N7Rjk5+9XWLo/LtYXIPu5hsoZrCCf9AqmLUEDH7GS
z4g0br0L62l1ti5YurhTgNF1GSI3ijKse6JKJlWDw37pRl8ccd1UOY1C37nJyosfRyvIj0zgzTgF
LnLjtEUb/oFgdRTOm3Kp7eTE108ezeNoue83HqeJlN4aOXMUQsxwZYNqMELlqOLhHtD3s++p04+5
0BPzrfvs+UGy+e0MX8SvUDZvJ8EpQn1LXmu7dhh7mOH9K4PG2Hl5Flq+vwYjo/9iKIRw4oN3W7je
aGCGVo2e1jEFFRL8Lbbk/yxaEBqpd0lNS3hIu0zcmhNqSPoo2MiXCs4lLuWnoLPq0Oel8uOh9vKM
X3QabRbz09PK1UUsfz667u5HOmkmzDK5qXwkd45ntkn0H2MRI38grasdWxwFxQ1G/5U+q43dG79x
pABFK24Xr8hpR1HlrxpxDdK72Y17xXanW9QTjEq4ZFRIIGUmCVwd6Ps3pe/cU1v4YKH8EtZLGsHv
01HNjDCWt1mHsUdlwAdK6uixDnAHY6kfm3+3iKZ0gZfx32c2bJ/ScEYG5AaJ/TaiY759JySo8m/J
b7C5raJ06ztKfdAw74WxDj4JsCyFa7q2a/1JiUrLvreW4nGVMOSZ+DH6MTkJYu7uoPWYQ9BAlqbC
QNrjVvw/igIOq3U/YAlenyJgexiOGc+1OFP4P3OZuGePFJLky8oggBOLkVO2ulHqQJm3v8slGj9M
c5vYWscGA/okwVOTeX6qGB5jS5ar0iQEMqb2vGIFYswEd99UwrnmJbwqSOoTK9lJntoDVlkGkAxJ
vwtqskn+yEh4E8pKzUt2R5lYJMIH68o6VplXb0fF3vVr98Rr4Z2A0tF5trs/qjX//UtmRHU1TiFn
P7U4XDLLUMv0D3RF05Uy0W3GYj+QJ8Kdd9HCvj7rhKJdyOGBEsDzL9ye6N7D5/6U0ZDtBGldsDP4
xkkoPeuDZWj0okn2FQpVXQRhlWrLjKVh7gl7MZLgD8IhwuUQOTMp8o/OaP6M++Bu7vfK5Al3gtHb
mz/9PhaKzAMhEDXWOYm5RiHPMobSsIo5EVBq5Tx607U++WVHqSzhMcJkZxLiTbp8XxTTuWp6Ndnm
eNxgQxRBikpzPUjQcqWCRmszKo4GxeuYsz4s7/G2GJNHeqWBhop9dhHachr4syx7OkyfB510DFQ0
1AMyF/A47bFhaUgseGRqzpjSH90xYwu4npyGHX66ua3ryH8PHtfB3heIkcyO0FKhPjW6Lcx4vPhK
HIRCdUPBzC/DLOyF74uZJk1ynaJbsesalRmpBi7+c9Y8TQzi/HVIYchVg1KywfrXIPnexrmslXtr
oUXrabcR+IwB6W4SeVbbfqOPCXhz9Ey7XNGITBDK7k1QGCYVf+nKffm7I+XAoYtF1GofRIjzlO3Y
GgpK+fCuThh+RT+JqIWUncANXhX9Kvg4+XJiJIDUYixHxku9WlweYgDzcsF+SSWSmQmJsjS14Axy
sqS05ivtjIr2iqWPJP3r+band5uu3vh2RDNuUVHz+FV0S/g2Tli762/hO0b+jlU0xjzRSO5kz9c8
J/YuvTtdX+a6MDfmV4u0Ofg48KHAp34vQE7Wp3SQ0Caw+zbucwo0pPFfqv2ZCuDJeu2+dqs8kC8R
2UY9eVsGKn7snfAmMFHjBptH1/LT1NPeX8DnCuysFo3zpJjCpE5fyQ5EJGmig7n/h3md1fmE5Q/H
YS5a/QalBBF5nZ1KC8IZBWId9+tdQkc/Pdq1tlrqzejfD8yjfR+01qVvS+GAjF+L4eCBVlILwHmC
mpWrTa3jhAxMYNqKQQ/pdsyatwSLYsnRS9RkSjR4Pug6MDEKYyOMPwYn+bWk7M8ZwCBfnXZmZ+i2
XN8VwLdZgLpf0CvAE3CwkyjbC4nEJlZ5WMv+0AmEUlp7RgCLNGHSksjVxTIV3eU0LOG9TLSJAOT6
T3avs5mjL8gss6lJ8GySM2saivtnDgknQanqcDTz0J+48I5l6amqoL5rsdMlNa77iSs7wLIRMJF3
5C8yt7mlARRk0qfBguocD+dSv8A9xrOIlvmCs3Qu7wUf4CSByt/9pxg3bPgcNBnTU2ucclMXZTvf
WG71Ge6elVoI1n/N2yIbGGVOZlOZ4hKLfjOeVCNOi+Y2ZE2SruPUTAarob+QWDuECBe6Pz0UszNq
qIH3kJvPNq3q0WXOdEJwovYzYD49Twucn1Th7E+7EYAU5NDBmhLaVmpi7RgYckTRLzQ70LbHhqkf
ipluP13yO+9eSEMSVTexlQBHHxX5QY8d0JxDwLJWIu9RF3t2qVGpYj2zYgtEuhzUqXayR0JzX6/2
I3sYN0SAklUF2eYb20gZB/Faw/0JmFyViwQnto8mG9FR1AgFx/W+8Tgr6EMO2Mcf+Ce/UXmMwPnS
RhFjwLBZ/YQv7YIT7HcBULIK065BFxNxz9+7SCMrKxSlLPOsIHwyG6sS5WkqAix12A3CggjqbSbo
KEk4RCo1JCqNdXIRi3cWCjhBEKAyVQ6qZJaOqsPsk4DmGRcZsKxXUA3uGHRyjsdKMoN59LqhyfCg
4lsByKVRn4EEIVTBZRjlWM79cj2zjNPBQ5gCfQwBRbHCVLhNiQZcV16VMbzEJTFTy2fq/d+5+9dn
mShh1tFvAOLzXIbEUaO757ckzobwsSR7z3uWOxaKvn71hIxy3iGQciQ9CMYyBKDinNPESy4KEUUD
v1n7WLSiok/K1zhogUyszg5lAbz+28LtGZwa3960gPkmZZrbAyE0hsnTn3vP3WUmYpKqKz2MPOMY
zrANKljTqG40tsTnoFzNXZqQBDnjnlxjYNIPfmxbEMd8dgBCbeOrxCo20cZQzvtQ4i1k1hJCPs3X
5eTEIbvBd+9t7HH4/PV583oyB9KL1TLdECFEdInFsC7AuBIuINdvijV5Ek5ZZbg+Qgdt666zHhzQ
G4AQYvZJU05EifYHmCcTQsa6xo+DsYBxAR0+mQ/BEtLRdfc7UrW0VaFelB5F+4dVlKDfs9V2z1zz
b3Sgiq2SvdcTIFl6aWiExrfS8gX2YHcl5ELO5/B7OANbaYmDNQvxX3dFKW26rxsJ+qwKWb0KfZyr
Gm1UiBZqT3TPsncbN6XVYc7zR6+DowbopIhW9ErNj/GGOPYGkpFz8aq0Co4dPzfP8Ely8PFzYQ5q
wVw4RzN32IhqQohHuAw6QuAnxbe2wsFE3bxz0KhcabgNzNNpkPxOWOPaikSgphC7mx2ALZxTqW3g
mapE5LmaEtx6+0MuTeD18gZGfejpJjwGw+h9ZD67i2R9Ch1ee9gsbijKRaNqfoD2dHti5JghRI/U
5wQEVURj4x+nGwM0xswAVNZVj0azDq8Lwa6inVG4ENERpstO9NkYlco56A1I9cLg1/tH+ZulVMfx
Cq43ejCPh3FgD6rEMXM7vtnXgQmZdcsfZ7hEmCYmqI6yueAo5BhupYz0AdcA3sPY79COBYjQNBcG
yQuAUe2Y4YiiJwWFjQWYCRM/65ue22CzqotWwHyKz2yq4Tv46R+vp7vpTckmL47RjZcmHRA7JEsi
VOtrQX4Kdg8sFYVW+fGNR/toaTjEIHBIclKUqq7NPNh45YxpnUBmx1K4JNgThmqflYzSZhHwTOmK
vA5W6OVJUQPEfzus4B7jKALM0JYSs9t6p+xlx/qMgsrmH4gRbBk72E3P6aOu/j+eICuOBHiBUHAj
gdwtqVTGjSCfMV/Bwu20932K5/9TfXdwW6pDUsV9N+obAlVGwdZ8Wb0sEmVLlR5rD5MahiHgD/ga
LlBKe9peRNv11gdu1OMPaRFjxBOSeuqvBID3CKIKe2fh+vn1Z3Hv80Wwe2W9WxxKFMRkcDerJ0tw
TFS/MXXtWh3T21itbKb3b+ZbVYPtukEmX+GaTBH3gNkpcpYqZECzwheHR9ojDFlBTyG5x2/wBkiK
EQ9SI9ccY9TF2kmilch2i9qY+c7IL0A4yLmqHPsXJLiEeqL9GPu2opXzPLu+I/MRCLLD4kgjAg+f
8mTZhfIYhK5MR6W0UqbBQJhdI5SOT0ux7dHJLokqMBq7Q3++Z5FDLOfxIR3wJp+8oavW8GpbN/uq
hZ6ffD+lCFRohZCLTbZZsF5X4xy0JnIrz7NZiiO0NnEflhvy26+v+ccaywfHHHpWrzSbItGAWBEm
Rp5qzVka1unnGUTUve1J2YmQy3sAgiiRqheKdluTFoLSMAicUNPUuuM8BVHUYROjNEzoG0uQP1zN
yRfA6VFPzcSs1CNSXzvn4zzMBVS7GRoUuLUUEs+MYczVsQ/nhfmIqtZs+611aoMw/mbdpWQSti1n
/8L4p7z8HF9sy9/bjYUvCytIOuqrVg6wz/Wa3G565orivHufSxecf42H9sQoDqHitf11+xryX+wF
C+SWmPhDAwuofb72r9Q6XLEMSpjNrfRgtEnQR7ScvXcw9H6x4mcb0A3QJwSBHRa6ZihAmIMjr+vn
InvlLi00HysmThLr46uSz4tboTmvGDI16JXIxpK35fjBNt5eb8s/v+5XoXrOrlzdpDwC2bQaxeC+
DUU1HTtV2KFvtPMwQ1NRDJMn/JEc/uO1ePq0nLbfM5pEi5dyviX82dRHahZhfnr7sxcjLGf3F+0o
JxCrPN6uk5osDp/aRqlUzbZEQgD/Qh0Fw0Gpj/jBwn0XGLBfjp48DOYCKTlASqANyrXBMy5mJyh+
/z1Y6g+Zk2jFxIstZRBX7QaTpEPr97llWbAghw4wbD3G9O2wU0GtshXw7mgr1Wa2EBIfMD9K1g/3
PWK+OWLDhoS7vpwi3KOIOu+tVI9xVcNdUgSOmi72pIuv104eqafSczzO89Fsk7FSrHBupLge3fqu
tWXNHB11a24QtLBV2RCY0Rr0NvECtbwAEhqOGEmvCaX4yF2P4RQUzfRaI+QzXi/IR105VEWGbPXR
eOe1WB09/jphQQRbgLirC9+U7pCN+KbJWLIqmkuX2PxLxXjH/sY6sEETL20LTrlm2IeCLXwmF0V2
vOfXDgJeDwOCLll5WTrGvC7tgkdRcE8AW1Z3eFDcxpZAPKQ0g8XKs7AXZLZdHbHIy94CjV/p8n2W
cgvSGwnCoQAllznhv2AkRzxRwBHiWOP1+dKIxcMONCa18dmNk08e82gW+ZnabazO65nIRtEVfX4+
8onmyiqSnfy77yl7pge6rUiqYzlQMyRSilAnoFIPNnFfr/r3LVDxdrMVXUG5cphttN3C3cd+AFbR
hnpkhjHS8jrAKzOFDolbltMkt2f7865RHn2vQLVWEBwUJDp1LQgPBEyBqYjfIcXiDsoerH7R7i6P
fSNkwLhGPVZmZBe+t7kyAGDDvNX+BLDRLg77LJdVJMg7lSmyqTbl/Gi3XoWxSuSieMtBzQtl+u66
CDikB1m20rSpv+UzWxoDx3OBrUPvB2T5WhjSWuv3XNK1NlAX/fdm7JYZLY49h2uQYgZdpvxtyz6O
u4K8G9EVymk6DbPqO3dvbf9ncr4Mkt7QCCpHjVFike4T1rrcvk9vTZZptpf8p+fZR5zdYDQSA6rb
KP8AyY8N28pmzjm09qGPVTulXX/wvVBOP5M9Uc+qpUS5ytK7jbsvlu+VLYYH8AhhdFrrNM7rmDSG
HL1oH2/5KcAOm1Z1d5Lv+gRpT+o9f5W98VPGBcSpEjnwPX756IIcNVWWCr/E8rxUagaZdeXbGURV
kccg5E4RBg+hit+gcAo7qlMSlE5NZBEx63lBFQVdLf+9tbG/Bgwhf9yji3E2eZaE9CtEwf6MVBNw
DS4L8QCQxZOtL/6H7miGfVyyChONJH0i7eey+FCv2cGmAwcalpa80kTn2LNbWwkDLkIPBT+bbugE
/0xeO8AQV95wrdvzVaV4OVMLQ8zN2x23udqAh+azw+a1YABax9REzqTivxG+vI3ibOylOkgZEz36
lCqudrbcdRi7OXb3r+L+xHlPlLklcXt6xQe8+hXayLi5ZIb8eooQq82EoPUNkqtBisFULRjTMQgL
8yxf+EdaBCuGLMVEJdkordOk8j5+ZahkrfhiQt/4CW2KmGZudB1/8t/OtFQD29s73tK2JJoKxIar
ClxIMkv8i/hL7NyF6TQzonH7gE+vQx75rh3tWtkbS98FFNKMPf2JDIiUobmkPeEw1FRPkDCHboWF
BTal6dGwhNMXb9iojDP5NrIMT1TWtdPptsHmWLyb16PFLW+dzUkuvmJV4z70vYb42KdzvQCGN4dg
sMfa4o41qSZ3Ved20DTtkXVDgsilZw3hvMQzDvLc0U+ciRO6mHwzNLw5+Irocr4N5cae9O/WqIKE
zTAltG44u/NJMCoPqRpkSjQI+uGxwjbyOYs+kYFTL1TeS5LEwM2kX/4BVXm2tDMKFydvH4EPK0rm
BcPh2sSkuU9Hxrh/QLT3ocA4WmV2eiW9iDv4tvwlWzrwqncfKg0RLhkyVkVoqByuMYuZBaMhxgtw
5D0fINB1ecSSTv/CYaNRitaCi5tegqXnL33DaAEi+erS7PYeRVmE7Ya0ztuYrsUwmd1Rv/k898cS
hxGaZJbL79zanVlGY2u/cetjHi/ohdsrnAKLx473vwOwo/lG3pd/4ZKDVHxvALEB2SrNuu1ZTkuN
txvPjCbiB+gmADprpBq5q8G6O6oNciQv/5py8IZv+IztAtNx8uVwzbDW3Mi52kJVBjMdE6Ewv+kx
6HWq9OlV8GUs9KhSb+qjyF+DQfVKP5QwRtFn4/M41iTvxIOBpI5uJy/Q2NspJ1EMYsHkx6v44qrX
FWu2RuuqRXQ28ac4c9y3EdIFFeo5NPsb1dTghSXClRPGGv1U2qkt6ElBPHgkAwINenFJcSjgTnDo
IaCXCka+jQAoWmfPDWJDrK+7bpN1VKoP0DMNCup0RDr8Et5DWFukvLSMEN8YFqr93GJt24gq9OAb
nFx8WAgnwxWmhn6EDgEJfDPM+6JnosNmwJU45zbvnZqTqx9eQe5x3rJPDxM3sEugowejIlhvrbph
bi2ql6Wu8FiN3oFzQ+/mGoY9PM2AP+T7QCprs+VBugpgKKa6TBkyD6XqVL94aTwV+H/tIiWCGINB
mlklX1Fujv2qfXSCrUZUi/RWOvijDusNFLCreD4VfxjncOpQ3VUYEhuNQPd5fvz1bvStwMq/ifiT
+2daEmViv2RqH7ggRn+E3Haxptuo0epFZJ9vu6FzgLuPAprd6mlRp1BSBBSdfVcDkzOcPkrjp4Xv
dy4YF++tsehKTPIJv7mlz7DrBSZKTKKe40KoZYd3eCfcqydRbQ4iPbhA6l2xN4NUE/eW93E3F826
AVL7Xr0dvvFJxPrhIRuSyuQz+yXbKWCLf52eZ2dxgx0avwhM2WQYkA1Q+hlFhQMwIQezXsmQjtIy
h5AYUZcCp3aZJwoxwEXJZlH7I8yv/4HO+ml7XhFA7YW9kWFlbe0a5qZACggUTUQSmO2kyOGonTZm
9PwOxC4SJHJQHPrUzEWtPctYQIXv/Q9+GGZOVh2TWGLSBEqbvx3I3zgfyFEPVODX/m6cIOaKEky4
Fiw99doqwmHBiZ/oStwGm/vdBHC6jVt2XIEXPUPerwrO3pdI8Kijj23KhvScSdkMYYlvO4DR534g
ygLXbr4Af6hw6lcOYIvUSewSMeEbxzUeE2S+gPCqaOCjCTnygPdtxdtxM7OLTF5iCny2PVn6vd/L
QptlvdAEYjl6uaEGMs+k4Rhv42fKw5nsk3auf9+tFoRbgTB8+wuWwaI+jktRw/fdQLdTm+1aJAhS
DcLrWqhm2YPcemV2iqRVS8qOtIyiVEKhcF9Rf5xYGh3+vUS7yxhTNWhurtK4/e9RMA5+hpDsFvuX
44TSDgaFjmmZElP5dsUszNl8ybTEFM6WeAOftBi+MrrV5lqnNDHRHIRZ0YP5PKU/HpCTkWghtdfM
V06j29PZuvc6PwkhJwbaJKkGpvq01lMoPNsGfiEnbBDCxQOleUr3f3/UEGDjPsCnK2rZXXqPMN+T
H/T6yI/kbOcR4fxNyGwEk0wE7o26FO3JVvYLhq3uNDB14/PmEHalb9RuLMGjhbADY4g1DzqScnt0
8/DANPryGFYPIffxhnJ/OtBADqQiDowRONg9XBqmDE4kbfTAwVoJsSGOduQ3ovuAkZ09D9vS9pXn
WgbW2se5fj0wclMxUAcB2IVtICKEkRwhakOZd6yzfz7ha6VEMHncqF0JHFWMV6f96HcF9a0wAlIJ
tofqQgjb8Y3TcnVvj5Y3bOQaW/b002OAqYUJkpNhZAagSTLso2F+hhHnT2rWA+kCXLpD85NC5x2D
crEuSkXf6CcMptO0eX1bpT+Tc02p8woriWumUvj6BwHOabUDHzeYdmOBgij2uCtywJ/osIWOnwHr
f5FHZhzbv9BZrZxNwJn9rwoUTMKCZiOvJpr0EjGyhnSW4zMsUBlkXx2nGMGOZ34JhLSl/FKnrkgE
FQ4LgFbjS9rLzm08jC5AivaOLIlaAxGPSIb5olz3RFqy99HObNNn7o/dF+WsWeeJkEaZM+wGd51z
b3/tPIFyxgaepJi94rzy60T10LECBPAMrlXitffkH8hOH6kOLpQnABvD1wYn9/w12vrnECb+N/XN
fEeWLK0iLL19wOKxt30VHKWynlg5jVPIZxdUZ+XbGVzJJQroyCJzyksk9baNmvT2IPgt4lvW1xpn
SabvR6IllkuPPDcGSZe0YACYiJ9PBxY1Z9nVFE4meFUqKr8u1dSoKOlBMpWSvCQVgoNGawK4aWp2
ws1hJkNt+Amz3sfQ9UXmVyOK+X1zzJZa2ymPmgvAzx6x5Zj+HCCo8/M+NDs7Nku9SgSaKVpT1EoM
ZNZVgFag441M5sffhPFYWJRaOquyzuTlUSA/Jw2EtMebxw7P+1iQlEnskZpmwPOo3AQYWFIaIjQk
Fecjp4aNPyH//xt9mNn+0qUBOb3bw41OmVFl/QwinLncPqVfduQ/hlOGvv7q/qYof7s3PuuH24UB
sYD6RthfGAqTtvePy4IgcoYsdaTYmfHtiVO52eeIl82K6Z8vFVkzFLBIcYNGEJLv4ZoEJPpl/MR+
TN/39o46IaFt+fGv7zzXOlBElvzCY0pmITtO9VOiInu/7coTwSHfZlJFyxystX45PcUkeObKx0bA
hKSV6NdOq1dEYaqEcZMMDFVmZvqiPaqVNfW0XQenD7L66K2OZdgSVvqDp+qXcbs2Mf08uxNTQVBN
DYRi6tpHxMTN7HaDXpZkuCK7u55jkgudgsN9k3ojjnK1QIS610rwlFf/kcWsVR3KC9VVd4fUx0mz
iNzLfMQqaRzww7jlvIjOZ2ozgiqgUMWHmfjjzAM2TZIeh3sLLIyV35xF4yzoKuoK03OMHT5v3U6M
+eAV4ciq1N11cv73Vq/h30OJM3Ab5ut2zx9p4BkYoRXYpzOX+VOmPbOjDe5YXr56pr2lJbMaNtoZ
/HEf1Ei5+acn7eVyPQSQ/8UBVn00XLjguTo20OKuul9T+LfQXT+QZyVclQ9Eup9Wq6RitHKyluSB
6wP5HeRatkztg2P88E9R9D8qK0paZ4dWyqFksqY6/8CDeRttj7/kCFxze8OSRGQRLtRmVnKSSSJX
GvEp3C7nTBZ7gN43xefnc+WLAWY7Yq3ViB6DQBBqgpN0QueuXkXKABdewP6YwPn8gpbGeEd1xJIb
u9NBcg99UxISOaChzqLYl0wi772dd8ghuBuaaKPkQwXe3d/XbQw3LoGTBJppki+3YzPJqUQ4lDpu
fA5aODTE9M9nQEda1LW3UY0yAPLyCeM1RLR5L81do2EZBFl00CEbBtZA148K4SZCyOAICtlQU7dZ
Fsm3xLz6dNjEz67dkY+LUoEpOGsjMA0CwDp6AHY3m2ff9tDFy2NcbLfYe6UEfDrQbDCzqB9lvKqG
T84FMP+yP6U76UiGxWbPquVKphmQdkP4WdalBcX/vLw395bEoGt7l7UwqHpTkrSsRgrMFTwyacJb
mHgYHkpodXwIESFxLjMR4iMdwNFHKuvjfQusgnla7FCtOCFJS6o6m/0uQ5qHJHSXa6x058NtVUKm
PRTVIpL2ZDfFUdVJxmY3l63FkkkHMJnnNvWyffa276Y5lTqm4w2jt8bzRlFFnQNvCoTrn3lxmOLU
WY5TfvPH7zJuU3aGPbkyzBhpHxpLfo2utd+7Pb2aqK7UP/yqsUKKCrMoTb3FhM4T+9nqM4UqUmle
49PftafdUOks8Q0Jx9mHvH9C/V0JAac5hBfRTa/VayIP10LhV4QQQFiB9KCy3rqDcPkDfJB0phub
C3mmNK7tPF8g0utzV9A6OyDyIA9J9gK1zGX37LNuz8k1+RxxTzqGYfHGFoCSMujQO+H+9fqT+3/q
ammrrgzes84HHX/LAeUUbXjvFroQYotFmi8eHEOvNBoSItZoN/oLzA4DKieHXPPsmw9deRAsCVog
yqQqFzpjdCUvrKGEgwHSigAZkkqsMI5I17H8Ec7zpk442DR61jH4O3TwzjAmXaAD/EgFnJN4rZlr
4sPII8mYXNVFiPLyrC6mvVXmqZMFpIm1kPkYlYT4NaIyuPRSgDN5OZuUp4VzOz86LIlmljxpfHIB
vo//dEAvN/DEhT4NQL47f4orYWBQbjD0AH7OAunMblhdB2ep1gn/rK84c/UhIjUK+p6rX/jtXGLW
RSPDKhizX0IPAyDXJ4M4bbvDE7sN3VJV/rVmXpUeW75IFmO1iTBDKm8uUdYuAorTAcWFHQOOIOm/
JdvvKOlJcVpYemfOBbijm3r+dGqqQ6i83L1yo4nXKHJkD2Bf1G+dV3nhX87cT5LllwJD+3T4yFRA
iL6nf8JUDNcPyl7IZsmlIBH+Jt8+ZuBC3jzO+VazE0ta07KrAFgUQA8DIdYiTp9ge34VMyW7VqLX
XTW4QkKuhryrX6Rc/F4E2Ype82MLMQ+MnNWOV9ZRQwzKBafmvVTrDwckpuFj9gMlnGh7+D2xqEbV
lb+Xg4JDkiB6wJnVmUb6mXYQeHeUOrnZYq2oBkAmKNUg/KLXM7DNA5I/MVfadtyPw/FNzoZIg8F/
4+RM2c3gPsh/MK4oTWnYKGamRk0nlHXhM3YRj5Ic7lCn/jULWF7Si83SIBiOliUKJapl7wZgTRnw
Px7PE6ceU37LLcqi82FGkLhfaJVQeXnuJkdROO/VB36a54fbcv5iiqCmeNhOCw+EQkx1lICkdCH9
n22G02il6sW1oozMWPR1Rvc5sVQ4SFDA0YmmZ2rvRqvIcZNHrRp6XldvHVQ2t+yW4CRvW2gybI2v
gAYstXWOvTup6FgZsOJ+M58DEeli2/zJCarIBZVSkXMeGRHs6nL2Vy3IClYhVVITY0dZ8AUiDVAo
rSMt97lTADZkmg8vIt7/eDxqEy2M+DX0FwBrFZ7AMy81hO8GJU98fnAWMLkG46eomPnKiG5mNVnp
YLTX33o5Y8ny0k9LgkSFW2D1vlK6Ciyvq7VjdXU1chy1xB/7M1+lgklJokIdDJ+jP6K+v9s6Bk6o
SrrO62alFjUEiGwXWNuVTaG9TguC5I2o00jNNGNTLzdskp74fH8fSyp4u7KTzpvN+Itbtjh+/zvq
hRQzT/tM9Btzb1LBuMyw5+sIMByi7XRS0gzuLiT/OIb/W9emDy8jtR70pK/O7c3G/UnDgcJaQ6Zm
+xVjxzQKSJvGdcxdJ5gPywUt4BkAL6qncqUzLGHa794bm0+DnbrNgSfztqhckHxDhHTfOLfsetP1
LkHJJyVLHBIBVOb49hFsmXpYbX0qS+pTYK/qiXxl93LYbM9A/HGmUnRQzWWzux5MA6sL81mMg2ma
DR9sWOA8kymnabpNGKOx5fCPNnn5cBTzJRwZFXPzIjzAGI4xdIkm2DdUxOwdwhUW+90qotPvSJUi
SrFVVvmwgyu/YQ96Nch1WaRu8RrTKAU4kxJ02kif+F8ACktXqroe5owzR0M9mXSa6ex60NaySnwZ
hwVm5sy3kwU/CGfS0MrN0L3Oj9i8mWA/f0H8OI8FWJgC08FHGUOJ1vn8CslkjhYA0Cw73XOyvvyp
gbSztRrC+INvWl/AjQ0UR09851Oq51jq1sxpX8cZLjPnBYl8LcTe4ANQeirnLwnwSscr3VwXPeqE
C4WomL+R7FHKZDo1+sf9QgYUL9N03T9aipI2pNZFWHUOtUnz2XOgADkPwIJ0RJZDHkosio7/Mc5v
8mm5zM3tl4bKcqvdJfDdmWrI05HMko0Yt46vLiFUxuBRzNe2fO3/J47Bw4dB53uhCKExJBjIdsRs
YRnkcFgwVmNgYT+O0Zt/VA+h76OPnY4QBd+0gjbZRk8E3lSvH5d/I0DRyfOQi/miJC9cyLC9Xj+O
jzSyHOd1D9eRaJCGXfSC8+RVMa1l50PVkHFXNmP52yVR3r8A5hvnSTCmokPTd4zEUlBscepculqL
UeIyKP5ZILgJnCipBJZAaPHIvyyDGpB3i/eKytN4Ham98wJ9+Wc1Di+CM57AwV8H+J75xng3cD74
IOxu5OYFgsbs0zZYmPDtnKrStSZ2ekbnZU/wtHs2UBtaqhREJnpjvKGyWtViov+sECU9XqLf2Xtd
LDOln4RMtWSZlO1kkXR0dJEyIA5izVU51upx0RwOpgtpsRZqZB9dY6gwFOME+T4LRdsWeEkWWWcF
C7HrjnHorBYLmRqbjM2tF7W0QTma+XMLrHh+irwLn+pJEYdtDyMakoImWPq/wqTXH/sJwzpLQLRs
6E6xNVEhY+rsTT960Z7IAJPGECU8GPdR2f5NrWOJ0e5CN0AeyFLCTdw3/8+yOA363nxKRkB5HLTx
ivwqDKspNCPQLicRkzHIHBwonzL8kWLd0LgnuyS6YN72uOZI6BqWEENwr5PDEhovsln5d13Pq+l3
c7351S1ziMzUHULQNvU8c23V/a50MtbzUHQuVgzs2nJ+0trg6XYZPTKzJ3/FPWKn8mwzVN0h1UFy
PTikCijT0KPwLDx/LWlIXFtutey62RmjrTM52rHVytNFLl3yOijRZY6FRacMwrMROWG7UClbPmHg
2uspBO30f4EpTTaGcGAZOHeY4FFi4OkjYDsgdcERcFDULGm3mz2/PShF27ryVW+fDp2nKALoqglu
OtctIIiaO2UODT4JRY4POMFFIoGWmfKqZrY8idXrjEujKL0oR+E+Jf0rY/fux2Cjk4XsJBrSymXF
+hcuV7KzBQZBFSIp0uy1UdS7Nz1xlgw55F2iyOtunZvH7iFpMkv94kqIf6IU34g4KspriQNVgN97
39UkyfYyNZp3IxuZ+u5F3d4PiJozOikLWTYfhapwh4vNpqRRUd0BFxZOGYgco9WE/N7ka2A2vZu8
MFuC8BfPPdsS6zkXE2vhKkivwdXyzjjCoGxCEQ0+cFcskRGd/iUwo3lG73nFyeedo9HnBipNjO5d
HJFehqHeaChtSuwUrFszLhwlsEvAz+qc7YxVbCO5hdh4pZ6PGpOukBZYQJA3qoF2CGU67b3sb287
/nrQtnuRtjQVw9RHBc7kwUB+J0qqACllw2N+xRtUAM9BhxdMBJ3zefZ1xfTYA6FmTKQJpuCrBHtO
B2/RSwu+AbMk8+5DJaN5aGBvgdcnK/Zu2K+c16GeVdFw+94i4EJK395wqDRcMjSamYV4odNI7LrX
h58=
`protect end_protected
