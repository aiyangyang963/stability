-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BtbRMfIIHp1t74mi8DwZmZ3kRo6kpWlF1U9VOEE0v50sjWkZq7H0z+rtCPYfl2NsQq2lPhRaCs6H
ZaXIH/YVkzTqQ+QuYTcTCmgWD+p+dRiN0T6R0+vrVFfglPDj9e/PlEf3LOOc/k7t9uoJnSSuAd7i
gITCiJwona3E5ZY7m9oyDLfHFUoLD+vYI8k6vztLLdqxkhwvM744h4FkGblTIWGyDa+2hyuBsMUm
na7bCOfdN8KMYsx2b/Q/jp3ksTw+xalr+LA8xKIPO1Nf/VJfJwpqysVl+olI5rz4NUbLWMPKP37S
U1AMLw8/iyYrrURkLly7ILywV0R1utI9AV77EA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
SmNe+eK8mqmXyT64n13Aj7sJxMFRdLzMQYPH0KsEFYFTqctU22zYaJVOhzUd0yV0aVNx0PP9KZOG
vbJQu8UVCNaIwv03uQeqTWw1vHnX6kl6L25N4LsSVT04PUiEGK03w6sd16oxgnwsuVmy2RXMYkc/
947/TGiXB83KJUa80cvt/hwBh3TZqH2zNvV36Sx/2pJ6dwHKFL7/j5SCxHbmrNDziyS+6WXx5Zmy
b0DcxeRKb6kh5sBDH6dYBnMnzdGyleJdWLdRL5auj+4Jce8LCdinUWlO4uovODJzBkSjF8oqHKBa
KF845a1rYlUWLMYim1OL6sOABBSA9VV0GFW0d+EtOoWzrboLSLIYDQktGTKhpdOTvU4n5nzVFOAd
U7HrbCd4Fe5SbwcbGrBKrAye2KB68zcrGPwQK4WiRUxc0zEaFoMsgLSdss5fb8mNAKCtmRodn9TB
ofXoam+62kwpEafjfSi/8d5f6FESY4YHn5VVxC2WWkZOY7G/Y90AOFLSfiVme7BcX2Ci5bPf0qka
fRbtlYk/43nTQnJ977y9VImWX5MdQFI4uV+e6a9JVnAz59klot4bWxGgt5wVWTsSf5dQw3/S3W46
5Apq9+8aSiDgsDlgJHSjqGGsFfNbsS2lYC0Mz1g7HFEvj7h1nQRm0KokkpE8ZYBOxdrEAWbsFbfB
xaGufpsit1lUrUXx/EfSVBTHY5E5W3l3jC7fYLRkwyBQP8otBjhJaQyLzeQdgcHl7agspRSURzaj
nNE0TB5SOJ1KkCl+uoFrcWY/37rN1WpaTl0lpGn4d1XBWkBO79PYAkELNIVAe7mg7F6wSXcmpH+q
lesEDZmV0uF7y5ysjv2sYgbt50kmu4HRBqCR4ONv2PAXDgmQqhlF7uxLq61QZjYTF0MdWRp9bBE3
5mY+BEWA1h2oWLBvV3WwO9VmsLeswecUK9EHynsi65E2LhsZn0pYlhBUxIcND73dE91zLYnYk/Vl
txns1TlzrOAjVgb8FlqpVBjuqbHtbuL7PQEv6XiYau4nE3SEshazbfBku1w6ERqzjt9EfDyyNjKq
TC59WFJX1hYTAKxHhntMM5FTm1WerPWhKwTm9pJ5QzRaFnMDEu8idUkJmkFCalH/onAnYgfV2XF+
EiGRdWwKn3kvk4qzUOFScReVRrTWDy5JRQC/faVVKXtLr2WVTW+ajgtzRVCbNMp9P77BLTo0xfo2
bIZONnZ81GqaK/ifTE6A8B5Pu0Tbs/b2VA0d0XuFMQ3UXBF6hEF9YPSof7V0AWBLySx8TzC3tXFz
TXT2MKMKGan80Au35QcYYaYpaTZnTOQ7suR1TEWY5IGta6pcnqRcSqrQp7+TLppymuOxyoVF2BEL
Uhma8bXhRhexFa30+juUwWUQqu9g4emRzhoSBAGTpBOX2NHNfK2oH3FkwZ3053uaVY6ce7TDCQtC
pknJ6AiuD+HLa62Os/H9QKszHW1daZwsT1jOP4OIOPcMTV51GTioGuQgXxygLT4cFTiGDKSYdlf5
pK7KcQ9pefkoyzejUPHOHv2WD/ZYWph2Z1jIT3wNOhkLfuE72ngD7vsnBPwNf9rPJHcAPVo4C8+M
l4ERCCmp2GT4kIM+tfUGKV78RmqDQ5koVi+7nzKZ4DoItwldq6osjycmlxKTrbieaZFJhd0XhfCW
LUjf2I2GvzyOWf37YZs0IUE/BB69x66oT7O/XboKKH4606KhumtNbsYxNpotlO40YE2ejSr/P8fD
OBPTekZptUKk03NH0Hrq/M+2wtvJP3Ug7jlroZYiZpDK4tsX1xdTARHFS7K80oJ5H1rTtdhoqXC0
QvT8iydeNEYsk+IEzXcZcyTGP2LzaVcURylzfCLtg28ARWb+4ukjyKXPdtJESYa9/G5scvl3r9nj
bcgGBXcxmRmblsZa+abJbz+D9RWPXztGHDBUno1Ec7mhkaHRhVtMHgaJzBCBTA4UxSxLlNiNKDJU
0UgtMbgGbuNs9HkeUyLtNY5EWaTSw8Sr8drjpDZjxZmrBClndZ9zOy7E6B555zuigTNy8+OJQt4v
zLcZdZ3Jx50tvk7ZmMwejHlLyNW/JL7icAEK/SwwDZo+XJ3wXwowk3GfWKM/Ydgz8Bbxv2vBTj09
3BACLv38xN1mY6OQ8zDWKAj+YS7tFgl5mvQQhI6vqAhLJz0mbyNhxsrcxLKsSqONL5RoNrQO3bWh
zifXok/TU5bnDUczH/8SzaBA0rN7YsaTQdAfIiKg2uBiPOGq1xerdYKbQu2aWrrVh5Hfuz9BEvGF
STDrT7cYUvXyBNXk3y4rwbGTXcVaBE0iV0vNQse/PiMzbCyn0yK+Rk1qi4p1jxmlVNMSF0hbBtPc
f6UVQx5czSeTdVyH918ckOxIjEEFWD4ow6F3pAPUkfXiYerJcn6hSAhFfeakw+fZGzzQ6w/UlaC1
K3SOVaibaBrfqwzwTeZFxyJ+CSti8qS/yqSpJT8Pq5OuFWTfsHb9BnuOhRdMFVSRAkvHOr+GBgek
FzHA6xaO7zcQhDZET/YFq9BScvkuAcHjvY0nivOzttI5E+jkjxgfXMiy+dURmHhokKc/6Bpb8jvx
ZM2CG4J/Y3EnKRk1Pr95BBQtlKSslZnrukwrzU+74XuKIxaxNqtfSDe6z04Ie7CEqqYQv2LhLa/w
/EA7kz5VlxGIi6WSWE4cbFPrRURGXkWKLaCjkUvJWsroNZo0Jy7z6Je8GJcUBsGrNuIEpKg0HOoh
NAI5HnfhD+3lixopQeB2WsgFlc5ad7A1yy/yw+I7wFEW0el5bGTRB+5FtPOZiOURkIukHAmYIegA
zYcDm6g4kYSq/7dJkRmDAQiKyvimZp97XDwo9l4eEx4AJoMUTuoFYq3DqkmEHDRiDWJsmmEIP+3X
CzkcnsAPKBmsohCFBHC7v9GnQohrs7mJFTKNHb6t2IYeb29RX4nLOJSrmtXAop6cmfunSzTBwS5L
2nmEkWFzmTKPBG83QdIcRomEONwtJ2TVMMO0mj12+3LlHJqLo/GToM1IJWo4n6LrET2qtZBw8M5x
Y/d+9dRVOj2RQc7nDSr7A7UbNIgbzVgjCiR8v8WV1cAu6LFMrr/ehVITBLMGxPnpisqhUQIg2QOl
7V5jXNvwOlvd4dS3Rz9ch8xnfc+I4RqescfZUoM5FMm5/hyM1W4vtc/ytxRAsujtEW14gXnjSSfl
GVHIFOLMmbvG/C8megJ+W+7yvSTbxuD5l1E/DMPvlLOeENxTJT47Ixx4KL1pJDjXMgYhP53HRhMB
qHgq1w3ppNSMeZAKFS8ZFhZ8IbZYtV5jcW7eFtehseAX+HY1DIeu3YtbsHpom/YYONoFzmUGER84
SnPOMLl7Fop9/RrajMGs8t1shKgDTXO3hv3JngnFPALhQG/tOmCzsXK0R7MnBFUgA2D+jvYEkhWa
dhE+5Wi4EG4lxPRLzA+ly/buSpAM1HIXhidNwuCqhX8D8MCAbXqEK6PmHItjDdoFMQIP6ci487Nt
ES9RndJzwH+Rjb7CEaU1rFJHSX0T7XrjqcnYU3cAQn8Pho4pFktTjUV1iatmlDkZ3SF116z+LTkr
YGBdfj9sIVp49pGccXIzb+3tP7/HZsJTBpfUoZslygMDUx8Po94eaheG2ZjmaKKeCOCQLgQC6XW5
aqEHGQQfCTiwFR3QFQZKiR+lZfp9r6bHgOzhTy/3Ywa/wOp8MhwLly/c7unQSbNIz2jz6sG1Tmtx
uXG0iGz8A6L8rBacJ+goaD+4/GfntpDmXQZNd37cOhqLJp8CTgwTDC9MmiBRLLJz8fGYG74mBoVp
1gDYR49BxL3bPucG6wKJ334GO72e9W/IN+QunwY/VtoxkKy+jCsybvou665qSByDRB8kof7Ne0qd
5SXrHVcCJAbKXZakeSVVLgPXTgii5Gd8KOY0kOWcjMXKD4Fe6gkE03BCTawoudP+pWMMyoC1eBqn
QhptAzL5RvwdvorQNvx0Jicnh/1RF5WPSNVN8WUldNIgYhrZYCINJYbO4zS2z9HEPiurKoXOFg4a
PSMaDsr/w9XDGYDL65Wbe0u1DaTqX93F1+HDubzORTu4vrXeZsXhwTV9u8gV4eRRm4xRqouAau9u
2GNvDxGRMWmI9k01inHxZB7atBfnIoMkzWHInyYteHYAMDBIRuJi2GaetV3qGAMyVB0sXUUjMZ57
TYfeiQfkKZUHixmUVQvOvby6BsaGox435KAiw4xx22jNZdg9t+YzCcU6Mbwk4cb+70LilrUgN/kr
fz75MaPhZZWG6+R41R3QTODWf0aCfMsCCOGqBl4BJnLWxW2BzuiMTEoMA9UGn2f+3/OsMX/jtiJN
fj9sRRL/457XdRAqgvQEzlZXr5/L6n7WoWFHVCESCbeQvIDKrr5cnt6lXFqIujFNhrkf7YEZdZQI
SlCJShxyurlsw7PcOWw//tvjYUzR90+MXW5xnGY94GsE3M0sWeDzGOwNaFKb1POrG6mBscqBLwTd
10kM1EgDqxkj0OuBR9WphNH8ppMpAF2NZ6fwinZamhZb6+5naWPjztz5ZNGPo5mN4eyTTUNwZFCO
6Kwr9uesdpxTp5saRUmidgnKydm/mTodOQAKAI30zYzLZ3ItIEEU2iydeTCq+0xrsa9K+KCc2er1
MIha/6/RNjMjqYZaxfetf2zky/AQ+Fj6Y8flG1k/gVi4oyGHrMYlOJ6Iq4iqHRb8HKWajF9+yhSK
8VYQhgGn2AjwvcC2nf/ZP0nS/4HA20sGnIE1m9UtxoQVgjmng+lsRZDwMBrfYUELOKi7y9SbMX/V
FpcLFFRYO4B/tP7pAvRHFX9tDHcRHQNpX/KjT+S9mwM4tI6QkM2cMG8CMeK+jTTlzMniwFh4HInf
XLlEh1sO7bJ04IGVVd+NWURjsG+b/6BlRCNofHGcwE9yaxZvJRaVMRdWynY3n7PIWxjI7z0WLP8c
eVCCVW4jkNE16ySgY8mUdGdje5HkjVH1yee8QrKtR04sH1Uf+4xsV4ueq5iWXJbyNG0umYErlrnQ
jv3mJRFKphNQAye5UklhxrllSgWvwjGF2wgcCfyfEABNZjtgfN+Y7alQNHRjbzKl03DDK5v5Aom8
KVYTi629JTk27UycJCihaJPIscBAYwaoqwWZXAl8OR8xb1DThzVf9aA/f/hn2u3/aj0hB9R9SEGZ
EMO4SUNd83PE8Z9uIwO1kF0fxL4T3nZ5wf0e0TCOJEkBFFGxjvRP8wXuxTlWrMwaTU4SgBhyjh6O
CPHn+tuGBEBl50GbVETHXXcWjrR96RK6REXFB4SSKPICKPZOYMQ5tjNNKqR4pvWt7+n5DXKyT8SK
/+/VKC731PLM0I2aaOW+pVedYI2TSlJua47Kg6MODKEZ7tsHKBWOlptqPd0sMbfopL309epgI07H
08ozPl6iGEWs4NNJbw2UI6zPkvDr3dkFiVVG161zjFLdPtrVtYF9iZ71ouwMfkXnohNR25boJXnk
liS9Z3uhuKtlFF0l2o0fAiptVQx8K1KpL2/GaYhxrW4/22m1TVDQG2Ee/57pF9Zfmdd2eQs6kO71
LnCWryV7sOPUr1JRJ7kGT/0gnBNviKlzMEzy+IKY9y9gYYQLtoDP8lrx9L4OLL132Yxv3xWq1c9V
bYIOBQUdkJNfTAyUypD/M1/wRgDH1vIJMnozccOVVt32T8tsq5p8SzUMBYYBmcVNIins3uYiifp+
qXC89G3xk+2vAKYDlKN74N9B7XAdbfM9dog2SXvh+cPx+In0HUcttuDxClvQT607gXYS56W302Eo
n8vmwrDiKUsDvVtISNIZSYyGAhwAU4+LkdZ5J5PaZ3RZsT9TCAr66N823o8tx/nQnWxBeaIGJavk
05E3kKM3njaFDeo1oCUfZX6BcC4n0qiYcqYeJwhsoH4aZv7Ex9xJYTK1FSXhL8ailrEg9yI24gLD
QnCyiiFoG7DeM0L4M95pMlf6m1sQ2kItHfFB+mX2gWCPH/HZZsiaBbcnMmMItrqZl4YeidwvXG7o
KnSWZklp1JAoTl5X1mpE8bLRQyHDXR1gO+cyfaLwTNA5eLeHM9xN2XsZO+7ko6Xc4/cZy6W/8bh6
I/ZgVAB998nbKzyxRV/T8LviK71Oz09KOlnPjZSvjW79lmVRSadVaFvNOQwL5wZPclHxfQ2WoTaf
CSbaq8BsYfgmQPb8aLggL9XZI7SlvlDc0bsEYhdXvOsaiU6gfRDMPocg8NJYGK+m+O+UWAEYxFMA
OQV3C5UTTGMNWV6n/aT1xcxZO6C2yrnlNoov/vn4D+UHhBhPmXIwa9TSCkEja1V2R8zC3CHwSC3G
EavXlJEWITaksAGTNyWGas1xU1GgrsWnFqNOaNQlQVP2QURygWL34QwTZ9+l4By4zSG3nDAj2nMj
uVQQakdDSWi0Tz3GTE9xPgr+Col6TlmT389SFQOvPI3kM/g224Fg8sbmwkBARX15D/Ulil5aZY6Y
asfW+HVd7IVI5ciO58E4dbnuDYF2vFVVgglvmIUyfxcLDZrbW5sRQzVL67WlM7h70LEOAZ5ffVGD
V7smwYf4owMogIQVBED5G9YUMK6OghgxP/Ku0rTd2SL9LEI02b/C3LweWG5YzwS0131W78mpHpxB
95y1/Cn4cPl4njg5R0FiI5lZGp5NDqhNXkaHhvDcpT5vGnO0MKVjEfyHUwnN54ZcW5MxCAstjP5P
PjNa9sxSJEI3HiZ3piIdsLL7OHdSDNmzTWf9h0fvdNiFRSyJfroB7KAx/xfc1P0kwif8OKdzFHVc
4w1wDqKw3v4M3LjY/z1cyXxbVARm+oeB+FtlumBM/C2NsNmiPj/pz1slC+2F2g8hJf5mgSQ77W+v
wpLrKgQs+jKtjPyLB8LX5EObBvWYQNfp30uiBN6+tpMMyE1wSPH66vP/V7VjJkOP1wFxsQx6UR4Y
IxMajYVeISNQ1kTfJkO4Q/USCaof9gf3nrfB3bT86VQrx0OKXMaDfFjnXoeSkJsm9iiJjB28mazP
gqyHChBic+/X/g3SqcNTOBVfGIFyanFlBEmkPb1b9ZIHqo9PFWt0hXA6dCoTmwR58I7SL0o6SI09
kGSaEGAixc9faSLlSaR4MDL2VQeLJCl8fvmKdnrgB+oicw6srx4PHU/rD6F8kwfYyy1CMs6aD9xl
sKLeI9dJ2rymJOOlqaSPoorB/9EPomq/sOHVr1PZgXNFFUkfVQ49Xb3P4nMx8vjube5QUdYHlmdm
ZOuoPthxRFPf4mV6EMzObWTjOUEzdr3PoIUXjHgEuIYplalXUEfBqZltSxnafjdbZfXEgYVA1Wdz
h9p48A9CC4H5F9KCLZE17OygDpB0oXM0gV2aamo9OCkaPqmTGn/Su3BtJf7vlAQw0RgovrI7GMb8
t1H7qOWCubd9gHuiJVuAUXPvuWzMVajHQS2lagTjvgP4XImUTamKeiJQQOCWPoH/2pX7aVJI/uLJ
Iu+C02pe27uohVPMB5gdHlCTvn9f5kEvtE/1XUJ1b7Wc8bx8bVOrPolwco46+KeAFmK4nxMsf4Pq
coDk6xYole3CsJ60FTbsJHbkz5Z7tueo5Axt4gWj1CvK5HxVH9re9wLLYbiiQxjj6fQzS+KYJ/Kv
I5lAnVIqAAK/lonbTLYetP0pn1VhTvv5HUDd58Hp22BFej+ZN1m6Mj0KF+19vmjXCzLTnz48vJ/p
hR9iZ2Z1Qtplv4ZnbOUAFhh/6/dw1WBP1Opnq8xgwE++LQHTHaWo1grijKQBKUqBNfhF+FnZ7KY1
WqGBpNHtWsuzU/2shxcSgEgfMGY3rvsjc5ZukCM/gRqiuRMrbLaYdVZHO9r47KmIaQ+siBFMW568
WusP7/ryEa4c+ZmIXA8N3lyGupviE+hOKZthDhqS/DQIDyijf9nziQ93AsdsAz7TstjpZu5IFD0K
zEEQitzgBNLWPunnX6RYJmZT5bh9m92YYE1akf4G+jSBmlcKIVDp8RwdHIPQ+Iw+3HBtbm5Qpi13
Oq3Plzu8KBIMTzE3ZfXup0xV9Hyt3guIjqo0wQsnKT/ISfiPTEjkaseKGoubcj5NajHzzm7DWLe+
OwCN65aUvmlmb9U/3avLqSuwhTsMK8S13zlG/C7SWSiW0o+WFWVcVb5BZhB+FqJQlpLGpJqVXY1s
ApCOJsielzq5lj5vpHKsJLvu93CporOGPckV4TbNT9NqSrl1CODHHkI4RXVXvQDOrObtId8Qg8EA
GR6Q2CJRuJTYUtiNRqHiYgz0crANyLIHzdnIVqKXSeYaTQsLzbwY6gM4MshWL+09yMmO5CT9qQ8O
uUT7t7zFtLWBnnBH6aDnvcOAI76fFcq4vBl+XITSZJy56rtOkOQXgiIq9R1/pVAJBPSbtg5ynTNN
FntPEv7M7pHW4fFdOnKV9jpbEYmRuY8ZBP2uBLFxh0OFrZegF5k4m4bv9EuaZqHAi/oQD1gPdnbc
eJDkIC65FV9k+U6Ih3Ivc5Zd5K5LgTPtdVJ97P9nkvIX2PYSc/JUzCwlmJGSznNDjSX50WR7n2kk
5PN96EfJo89lTKW0RyiQP3Umcc43NKeeKXP0oftkqWi57VbZbl2nNPYOLT9zE6l8OfTCpEWliX5p
Qn2ryLanggyWoNI+ZUGJG0mj5R22cOn1DuLENTmmZYenSV3Uhf326XviFauOevRcTjb+fwHCFbzY
Ggo+342dnWr1K0LmnqaQMcIgrZKwY/SUPOfdJpZcBnrRtPNeQqsUgc5vnd1ebgy2w3DldbaLMMTl
EKOSgEsPnxsNyAWaZnMlTB2qlh/MK1Y1pFq5GgOYr1ioabTK/5v0r3CMdo5x5zdfqUxm9Gs3jbUY
kDIyz9HN5YEB9IUQ7p+QA/kFAM4uS9FiVKIQufUcnGC3n7qaaAjGjzNKcH3+cH4UjBrEhc/szRwL
/Ga+Kv6UEYB23eckWZn8wPZXYg1tryxii4EhibK7Aihbt6ucACqzTUSJWEX1+BlW2ebs1t8BcE28
ZFXY5dZPk/1SQlIoTKYsncgHEqcYA9bOsSj/AKFuegQQREbzkhx/2+2iJfCmnl7TnoPrwpakGSYE
uLtPqtJ+x5CA2UsB+TX/H7lsJF7PIX29rdYp3oQ+JDHVz17X/f1Kndd1POGbVQ/1eIOfEJne4ekO
BI4OHW/phUH5kQAWHUg0E34GL9QYvmeiPK1hfDGBSR9MS1RBqAPL0jiWh1+/2iMFZu1875yV2wJn
nmLEo/CehpaBe4VoTPNS3zV0yA9YyIIiI1kmJyEejOWftWwsnfyw/3acFvk0Ang7UwFe1Dsc/zhD
zrqL4mPqafNxv6YZygCA9r6DppdhGp+s66O32n3OsCV9mrmTSijw6BEtg0Xlr73AQWe9SFjJXcBa
moC+88T/llLhvk/6U1elXIaX2Zb9y9pIMMQOqHq0kwe5sazpyPYTvUTJ7vkhiqsQXg4TSCkdVl+Y
o9oSwTvRy6oavMH1g4fQi9cywNAzRplhxnATSgiXd2r80NC8rBVMg3VEzXE3YsiRKV3Rjoo8KICr
P9qnBYcVcIZEKFKJICt015TZ2UxHkVN4XwBA6xMx7OQCRtJxThqAhT1yMJTyTOW8OYytPambpqFl
fS2J5IEXF53IPsS4eDhFGhrY8iw5xIe7zKfssOvODYkw07PANVU8Rb0SyRNA3SBJVGaiC4sVnOnw
kepDzpe4AwhJp/BWgFrvDYIKLOWo7MS+QNCNHcRHfXQFSbsf4RkKllACEx2WVDBt51CkDtGXxPru
7YmAMNTIB6lTNYzW6dI6rAhEt9MMhXo0KPEn2SNW8J/OCSlbyAFfRpm8GMeEN+bleD55CPzGTdEe
EXUGtXabEZk1AWpEm7eFgsFZXjYwh0MJSsd2QI9D7H16puHjMddGZT1X1vhCta79awffkvasOShL
E4KL5XH42FRLlsLOpRh+vfxMPx1P9pzERuqrbxIchq3GnzDAVE+7/xNS4i3z7c/VYSZgwbPCPYwX
55omO9a3G67uXuw8eIK+TRJZ5NgtTO4dD43IrQCdUMnSFC4derKjsyXeV7u+ZGc6r4XxQDYVh3BK
4iAsMLYdCbuFL8pJyJsufywS3HiiKbHqAVm+GV5uJWWst/CLKksUikXenxzIDWxt0pUqBZNNmyOn
svedT7+Eiy2pAD22NtUvNoiamqYqbFCKRnRdfnA3S63YnDURuoQb/CwCJ8t4d4MNBPefU23QKwki
r1pb0mA2tAE2/j2h3oJ0PVoug9sYgy/DXo5VPjKZLlgj5UWtC5BuE5A/ADCJx5G1Ul4a1erobzWL
mmczj/oEp0HkYu2VL2E+1kY/y+V9uM0ZDK34YiKznI+1yT+y9+53zkAX9t8rt9uyUQ1Uvhbn0UV0
WwhGPLChib98AXtsbAk2oXTJv47KhSA6BW0wXKSPaHjcOkonc6px4j1Dq7K5ppl+i7CyiwORqq1i
ogW5dnTz6RstXLB0zPZQx1b5nsPGpgFdrtDWA2H1cWOTa9JzBw4w4d4LQ/FAqR55s6ZJNNB6397D
yD1yg3ZDkictAiuO+duKj2tVukXiD4gbSXKEB3gDfceSZhJRMc4sDGi8JiT0cs9FKiryjGMe+WL3
pKirH/J04IPOzqAtFlxOdEpxF6NC2h0Fwo3m3oqBwlbZaJcSwTQmOYY/hhQ1dJtnrgWe8kI0vg7a
F9SlSGnqK0lcm35Ofn1sYk9H6hVN8zmCiBSIRTPqRVSM34mbd+S8ZhZUJvUBpCg4bPI+rtNNdD+i
qV4ol3hoNCd2/W9vzd+gP2dkvXCRNJgytte/dY0P/NUeOEkau2knPL1Txby+iM9OnMp1czxTujkS
fxGdGbCwDxYF2a87MfCABsnqgEd4MLBWU1qmY0xQwZsoS3suB5EfaWRlKUTX9L4JBBoXkQP9DED7
eJZS1ExIyQf+ITmXw1appqMso92dVupLXtFkAyvll6REni6T/fVnAWEBquIJNqD5kCt2Vc7trVtl
NKLaLDCyoRqJSt64lZfMXOmF4LJNGEOm1rqpdAwMBf56an9IgwJyus7u6vZyK6e5Txd5qo5g3Qmg
zjHADieMo64eYIZ9Su3yozZOzSKFF/8rmi6zOM8Q+1YEYqWUHwqQGQ/NRti9NLKRzu+RbgZZXhPF
pk4976GgJavC+g6YYpbnXewoqfhmAxrZlOKhQvnzbeBbpQSCQci3dYjAVDlFK+evylLiRRbfc7V/
9eTmA+skIyyQPIgY+DGIJZbomfO+aGWYEfh+y2ytHqjYCgGmbd1vqjxmnPuDTLM6/Qjkz+gBEXt/
gIYgBvuiLeoCPuXAU3GXc/n6mJkdCeBQfMZcNpbHJlHPph6lgaroyobtroHzOcLJZEfcz8ei5lby
3bJQvOVL5fXwHFby2utCfgBmkjAWEGlrNuuxT/K7Sh9jAXSUTFs1XpoiQR1qzTrpa9m3PZTrBWU7
gfdk76+Y6N5etVgBG/7jY6b2gz79mSwrW55i7rxVqw4kXlSk6IuhOTqTvkkAHyo31anyAtRiwRf6
QJaM268lF8ytaiMGYVLPtRHnYMJzCE/o18WaUh1tlDvHZcfXinJneH2BfZOhWTa5urYtVO5hmQxo
NJsmHEn0gCCyB+hwmbwWdzOEcPrRbdNZpWWB0BaXZ515eCAE228SG42sz6SSIEzqvaAWkSCcFpov
Gl26aieolBFdvTsHMY6ciRVu8k6da1vxGaCHIXMUcGxDRE6IiGidvWOp4MPPf2exhFXM5611DSbf
95LUEshy4rm9i+Ig+RwyBsQYNSiVsj2/bgpiHdtY8nzpiazNkxMKWRh8IcXhq7dmABkY9IEBesy0
UMNY1X/8zOn9jpKgRnMS3nV+iVLI3ucX0bNlrwTakzCoVkdSbhFEYE3OPEsrP/H6uIEDEmeniFtx
O6THmFL50cwIGMJEF7Om4QJlxJ5T2OF9bMgp+g6YXoCAYT7qbtNy74Zqq+wzLsq4E1hkkP6rvJSu
TX8cTgLlJNLsA27fNLT84AqNUi8p0nfnZsU2lR4cLyZvJTtxJxfjkNaT8NlPrQ3fOnSA4gYMutwe
2wLK+5tNdPgVFEwqS+tp4byxCzVFtjtPDH+0orOSLfM/1Sw15hsFqzbc4+rmOQOk0tLxOkUT+5MF
PGxhZOeKMqQd0kxb7wQV5nbysj50GGLYNYovvrJz4hcNkCTZl6rMVN/USEKFTEiFmzEESyisdb18
PAQ6m/WGVbUxkImYpG5wT5sXd2PyhtQrxnNzZ9flEFBtxkp8g62yYvqaxAULhaUKfABmTAEckTix
suEeOekYHVS6IBlQ2w+zy8REbvkWegMIlWcKqyswHR6KTocFzsH2YfG/oXAPEw8hj+EMZTnJZOGk
GPBefJYL9YPsr3M8xBNUk+IWCXA5fNYi6PqOKlCgUee5B60sHZnf4YQpGBjp3IAJXQt2rOQzVpkz
1boQcW+KqY26jpFKSdmtFFrm68qJSBRV46lZLRDKGcvITBfcE3RlocSnq0OiPbIL3k7ZPh5wNCpU
ejwI98eUSI5uevyfpDK8aPC2H0xpof3oWGYKmXydQyTjdDgEkIdXR1QfCpWIJDgoudFfNSJOfH5W
7jryG5RDdcghGRKWoJ8wZkarWpLx5r5xp3Gsf0tT1l7cj33vyUoyM++s2phIqqwT4C7DiLqpJYU6
JsUWUeTpNI9EPCIS2JgLXPnVmBy2LDZ9LyykoOi+DCyn66/beWOEut56WRKZZWmSZZXm1lN7FwrT
W7KjJYvdEJSw20Z1q4QANCC/t3uTIAsk8LTjqS+M4lSobuLluUyFWYfyz4lorILQ4uKOjztvRJWt
ue0XN6WxkgOSfOmwX72wsIS1yNnTvSHMVyO3Gj7MYHolstq/AYX2NPwjglLh5WqiV244C4/jm017
CnAMvH3+2E7NwXPqrPwriJKHM0hPkxtFv9mR+9Kg8wNa5eTQlAqdStjpI0CC7vs75uXoSZPFOtCP
2qONdJV04wbwgpP3TjwqfjyhpXoGG2QgIfUhjAKZYXVsF6wZy26hqw4FSQgvkDLiumuvN57KE1Gn
M+Px3kYLmF4P3Vqfer4N0GU8lp5RExhkyoIlNsHyMqePxOq0WLbpkdBgA27eCDS9xyqE9wSR63S0
kaECcK7E0pgIHPbdBFyzdpBXFbMcS62dKTUQWaYu+UC92MKG+RV/HwhGM1b14er8I1h8625AAss7
GuKwZ4hwt9+or/L66mcz/1WZbUnzvv2kUa3uXyir/H7GqpiquMx1Qe4K2tAGtw3pGZ70P8H6p8lH
QYDQXo3u25EG3m2hVVo9VmAsWuC+jShSurWEbycTuXsBcQxp+ClINZvGdhqs8BwlJ9rwsYgJmZgy
1FaxNRpbZ4pUHbHvt0jur4vU5sW6SH54obhJ+h71T7EwxvvaSQzOGZpkNhw/EXXQqSCgjn3w0vjn
OHewbR/ToeA0SpNZ+mmGbaFOsx0I6wlgQhSJ519fsMFZS4V6EK6z5rTvnzMrJnkq03egMddPy9lG
4PIt0+lyRidjWi53wqCyeuQl2H1CTKgB4AtQT2lWw6Vt5MbrAcpaYexGHV7uxYxWiYJ9YZfle0X/
zGwMunZP9BXbp9pWtZQvPvDRT5HdKM0Tvk6RUW8KS34wlmvsIgzCnbglawTkp1pedokf7D855HCw
2SOn6QVafUd92uOGH0YpMpJww7MQ4ihPmtvKdaZV0NoUr0tKfzSMUzoO/n2IYsvByXM8CHm0vcyq
sJ+cB2yIiJ2EKMsIaxyCenY24p0X8batemX3vkPDaMxNJfuHwjKffSlCLnWoAdsPgN81LucOiDI3
oIpf4mJmQZeLBzdgPNrR/bphICJJPLNLgFu0X8XGCH1oBWwQzmtJd/LPKFCGog43HK+7VKTS2nJL
sxOiRwQehmhfivrvYjJyBQyZ9irtOHrboe+fyxm6QBODGu+VSChxLqoUDerS+63CPTEZFzoUwGGl
V3mVXiIQ5hQxz5/9+ManWiMg6+5maJPWxeqnUo/4Xu6e2FWMwAnabzZnyhzHeezahIvgHTci5LRs
91U7jNUuYgpI6Gm/OybRAEbUnHDJi/hoYqmnBhp1wqPOUXPBVzvsy+UKQJUOJhDtuANjm+DDIF+5
TXMnO1WijrX8rvYRoXtIG9xHef/4dJay1K3otVAkTgmdX4DBqRsdKDMd9CL7f51B1MWQDXBVDrLY
cwpobBRewjigG+0pxS06u5q8sczzz/MPgifpLC3AySxsJ7mhoBonwjTwnfePShFjpSxIVacDB7mM
7YC9bhBD5thCbny61hEenvUQH6wYV3u7gU3k7/Cflh6oK7/XmpKE+hO+bcd9+D4d+gD/6+VQhzVO
WFd29eGN0TdZOj99HvpCLOs+yI+9p5GQuseWwpbzpSfA2L6Fldd7tJWFTW+cLNr1WhGJ9b2s1vN+
iqo5gEjeJAmFYyRTwCD0NioPb1jX9pMNNwIVxnmxUql7y1OJXdGhdwFO7mUZsfgNo4XzaKO5dNaJ
R5qTvbS8lhAfdC3YO7c+BTVch21IVN1VPjOutNpkLSE2Id4VmhxWa9nBa/SKWRh6sm9Pyi6OeLe/
yceHMY0b7YOWiQvplAdktKbsTlSbb+GyVmlombrfq1eog/qxzwYrCMsVV5FsU14CM8kgZNJBZU/O
56JmuO+pMUoG+kW0jrZ6OyiWHmYON3sOzHD54VXyqXfRYYRMLz8F9gY50kTki4jXAML57KTSCy7z
n6g/pIycgL0XB7OEo6H34edP+3dXdwGpJscu+n3hv3d3/wu9kgxWgKQuwrMmA2HhPSaGSyaQHWam
SE+JAxakvkY5/r9T3UOwH6Wu39+MOMLrQmZDsoGVLwWvvCrLBnsYCMvyYu1YqTck8bjdjOb7HPGJ
pwNV7eyFpwmyQe665wLHrMu1+lhJZTaprfwSa9f3DDKOkaNS1ozhmEmnTAyZNnwhA10b4WC83LoE
uJGCtYacJj9wvZGk1cPZZaNY54Ze+J1/01mUrpTQ2tmv+SEL9mExUGV/b/KtyG3D3iUv/i7IqLXq
rCC5WEOdcfOktwXTyfzFWixyu9zAzkOFBy2lcFnvugTzluUlA7m8/E6DQNuMh5/OplfSOGRV957C
+BtSxBFD1p1pU+F164tv7BFyMqPYq6rCpL2gjaDyyzcZVJsnvDVrOYygSrtHjZGvOWy/5EkA3wp1
oNpJzH/TSO0ZsTvNzB/f4UjjHxuFybe82zh3ez+uruJM9Mq8jNKbXD1GdeDpg6dQ7VApHkUp6icb
YOBL/H73vI9cnthYXJS42oC9vwBw3x1XV4GVZXUIKEL6Pgyp5ahQkb5fP8hZcW5qIqh0lYg0iEkq
rN8ckkJITNDEHXJ9eRxWkWdwqC/Rjy1e+gdk67jzX//qHO6Fvtpf37Yc9aZLvWOfW1nyP3DlOPuO
FajafX+J01h5Y/BtsG+if9M9DYYDbxajD0d7u4SUHgIw71ypGG2PAic8tgQGifUMedV+KaCkK6a6
i6dA0LZzS/zacRy3ImHQfOAf1lukG6+9EeKkoXDGlrBAfwchtHFCpc5U9VAkG+xpog4YYMaD5MEq
w1aeFw4PoJTlPrgnYQlkBifb94+2kWXFHg1vkyZfXKgax4aNC1P0qShxYRPjAKI1wAjgxRb/TTLY
Niqlh6ky3hvVmDKGipdVoTVgP3+wCQA4kTVcCg6ACw48sA0JI31hrsxUZ96ZscFZpORFMZi5nKCy
xVtrjWUYf+KmdhUoXJ2lRoBJt+GlV8TIyKg+JQxJHYRnCb5xR1Vkqd0MONxrqaMyXAnCTqrCRoF2
ehl6WKpBWBK5WbST3n15ENfOoay0fG4ag3RvEwatrpxEbfIV82T+yoWOm7m1di4REpWvdoSSNQnP
vkXchudpYvO/j7FklY8LzH2n27H28sB0rVm7X5a+8uO1hXfS4QZe5xMrvMXUyGTPl65E6zlu56Ls
Fb8lkRISNb7/rJn15pLhhNRLJg5BGSbDrBMWls3fr2v0jWNRSLr8lCbMhwWL0ETWLHqopMMxaR/Q
t5i7J4PAEDlVIh2W0wOR/Y3K9UMJ+Yd5Xu7rNRsSaT/rSv+LrDFIYwyJwy0nXk/GASMzN9ZIbLs9
aI9EAJXO9vpXP3PoMVj9qtrMhswZiWEg2br4G8QhFNErf5H5c/h6fLcMo6R7s7Peu8IgmpFD2gWf
7BMQyW60egrJqVN42BOhRuyFS9D35QfE0tHRjVFwP5DoD7cotMbm4i4514thcNiLsnKabWnkTwhA
x2bJNV+Mcmyntqi9e/Ur+geaGbIm/eXV0AA2syObDXYXWUElJ04w/yGLX35d5sD2bIcQcVjQUmcN
5KdnDRQm/XUyDew2izAyVkn0pJFwuXGcpW9ukfADzF35ixtHFP4PolqPEFBuUOzWc1zkkzWnIlMq
P9l6N0au+hRiV5KV8JGM+2qjnXjPaSoePRUXVfZNwq3aoF9oUc0b2VlwBTngNmt2C/Ph60EdWE9s
Bs2OlfH59zw/jqOB3LpIteEDf9hcgp6LcxiGgK9rcm+n70YrgPPOIsWkme2dy72VzhG1omJ7/F+8
gslrVX8CPCupMTgww2syrTdFef7QITvABKU1fEvEyp7yuiysWw/96kpt7AlwSFnqxkSfq8RBoN8M
CkqsrfeIksFAcEwhT1hJjEnVmEj2QaNY1uBNp/GetWDbbICLOri4Zq6Et0KaXWGW6ouIaUL0u5hG
zy9/BUuiTQHarV8Rw3kTQhskM4Ep8DZJ7NroH4TfWcyT3CfzkBQKb3ayZRjZkh+IK7vn79OL+McO
lXtmyive9bVP4R1UCtsClZWHp5upyPsl0kVFK+YQnwKB6Dw7hHXKh/DX1dPwVjfKU/3alOzsB1Va
rYPQ6bQ7X38VZPISUbF/AE5LfhGBQgxlokWlbNkBLQNFSsjVkYhugiEjhxQlJjIcrKY3jLjn00Q0
4fLMoqtvg6sUEL0N4wkO81EpbvpZKtMWww2f4gqv65mYasmmrJ7dEKEMHafMh+ZQTJdq6N4C9Uor
9yune+Gt2VcBV6TUsphs/orwQQQtWPgDkiAzB7SNxAJjIYCd8FtEJKgtJbKZ6bBqFKY6yanRPwKd
4x3+eMSKPFlgwdwFnGVIKfC6n7yxjYUqqFy3MqzNa5eSlHQ6KKOFy8zdWIVcUrZWDEHD2/TKzkki
rdXfQTlM0vOPbFTvAZ+s9H370p2ys1MnZ4ShBnrtYOlc1lJhNn5TgCg2bivdrlXsFDLWO0+LXsEn
AuNLe8EuzF+lbnAecazFyGnqGLy3kbsQPM5rxBbWbMLNNnwOw0oawZENBG6OY6RdI3cW1nRosSK2
JkVBonxzx7sDlKUe6EAEp/d91xW6PEUHWMc/F14mViWMqwW3h3P0/U1otfelFmgSoNb7Y/Q5lOLg
WFNoGFWy2nsVmyk1Zs+/9Xt07ooJX/D4i3GO6K8HGm4TxeVUbn5A7ZaMDO+Kt7lKMl3ni1FgHUKq
goghtzSgVVJm9loNAdZA03fcsKkgCg7o615NVJqXhzV11+cwoUoeFB4e3zOqm0BqniL0LBl1P69u
Jk23StzRY4XNcTZuyzWCsiBvqZv1P6EZy0tp4BE2QdHyJqB+4bJ8N5xKHbJn8ZKnBCMhnpksbY+g
ili+pA6KSq6Bk3IHIVFC21Ss2XT1t89YDgHu0ZEfok2B2byHtlcscctW5q+XMJmXUiNqSyUYWNTg
t1b6oY6Iu5Du8RPUKjvkNhVq+zTA9yV2PnpS3Fw5Ov/Dp29hlPcQRqhVZrvVuyMLHAJqzFPl4QmM
1nxxzqnDqMLLo8CXQkbYvh9Ujg+sLZsbXaUTUBUt4lNImF83eFw2AxS8U31r3SVTkPIxBnTaxs9k
kKmOK0YJxPJBE/M7wWBUIrkDLzBFuzgogpPem3TnaMTqN/KzWPZbZxd9MkuScn/krCUV2SxGYmH6
uvtQTl0+C/vcPUPMGfL9Qb7ou6qeZnryjnb6BtU3AG9PaWCqD2/ywS6eNQMQLNMw2THUZ6x2t2lA
s+xGktrmkPqCkClQmj5OK509qdU7pwxRPRpHO4qlmxyPGiJmV+X0gWoMBSwqfeMZLcUVERzXq8Qf
Nh/DRIxZ0b5Rkf/wIyccaKUjBWszgSJmoFtkkw8UKnBQHdEGp5q6GfNWN3+RO+CG36BOgWqq7ujR
8B3xduhqBvWlDLmXY7+msQlf2R59jOgNuPgnwYiYCJ+uafH7NLkyP/WE2c74Myj2nO3G2xOHjy7P
G5Hl4QFqaVWuCG/oCfJL20QD5Lc03+XVOxd69vanctURYaE7uEelvKOhMeSy24iyKkwyv93xAUm2
fRg19nKxq5JpzEuzEEnMC9doizglnKhtOfuAb9CyYmgBYWVzo/IBm9zc8/kq7xnZ98/I+uj20ZSl
juHLKRkqLoWpL1UeId/Yal0x//+Sl243EMrm7IpomZcfEm+r3VHHhdsIZwiSZyvamAliqXWyOWqV
YCY1AIco2PO0uUbYNurdvEYKWaY64H5z8mDnTybp+ImZuHX9WMBnHlvkFjW8CLL/6h3fZSgHKVI6
objIKBVBSFtT+lbx4TzBcPwNQcoiieAZPZNhB/UbIn5C3PN/uCLp7fvVhoOfx6deyYf1jEjlbP5/
IvEjW+sVCcPeJ9E2Ny88FdJNH/0T8/ZZkdDfYCf7oizdOm+dzpSYSMveM7OD6TTUim0k/MmJZ+5e
9r+cX9KIMI/k6GjfS/FzG/KYHiJC9XZ/dLliiqnH5oYyF33qMT8FagF3V9XJE5DZob643RWnxgV7
Xh/ajcCB+9iy4loVGl8w1BiazSdkNH/YPnK00P1xfY8RD2JXrFglE03WPoX20KpeM5q1u8UCWM5D
Jh5YX1oJB7RHGOPKvKGuROYIrE8NX3028HeteL9DcWeR5gEj9EVs3XslX2QUaFgld5ZwmBkE9n2c
TRSHPx0jO83PUB41cOW0geTRe92Z+qGJEOba37dBWlNzFNRibG8M6oIjTRNMq6np/ALbyiemH8da
OOAfCvFT/TWDYfzmI7rSujMOfxwmsynMA0+/PghOb5JdY5RrBC34+WZhQJtxGjenCqn4PqvbAFD1
/uQM+x9F4wBuWMPF3+CYQy26QZ3YoJ5RDpwNE0vv5fR3tIgXoDSvUUgFPxGeNVXGALr3pyJVRvYb
EeC8nQthobsBqWxDgPLseLELFaPuEaFiSlYq/p+aO9WEQUEGv5ngX+yWcj8fxyGw/N+YbjKT0GK3
DG5T+t7+YPNtQnYzn+7ZdPmNfOLpIK+RteIhCSLfrhgd1FSWtjHiPEi3wLsTtN338vXijlxjaqTx
Hyt6yCajCGQ6FTSzrLGQrvcKmtkAJpT/w3v5JyCNVBixA6COtVrVywqDrjyejEQLy8s6n6BSoFty
gS75htJIoBVaZ5hhwRNA92FxqE5XYu+gA13nSZmVaMdkvSmAtVV/s2x1MfOvrxjnKDY7+9Fqt/HW
Fl5ofuSyiApePymQ2IA3i9qfb6ybhQT+C71L+nKlLYzc41yr1lUGhlPvZXpwkkvEy8Up7ZgzlCX/
4oYPv4pCu8Fhdo7dzz9bnfPjB5yft9bx2xi1IkO3pAt5FAP8eZTSFjAU+es97f5OfgjX+QO9d3P/
YxWA9F+bT8AfjcvOYUnn1+R1KCk9lS/Zvwk3gcysJzQk+m7vz+tovrisFRxaUX6fGml75X68ROdl
8dOuuhaAx/m+uemLdDrPVWI+cY/84jWz+rpuXYFMr09bJMOpeo7RIc5kFYxEJGv1Ci6moIiEj1pw
4M+bhzTpwnZbNFjhug7cw8Z5+V97x/JkCUvbXMSTnVaRRtugHKxB8dzQYw3luYUBusyGgtWkVUET
xUhP0QBkkE9IExPe99BvL3yNbxBJMutys17zFgEttrRARiOWKJh/Im3RlXVLsomXSe37b0/iq2mv
YJhRYgpzV8PgOk2yrBLcRu0Ox5FDUSMxmxpUSpX6TUHJ6QB7VjtmNlz3dqpjYy5LEtgI7meXfKK7
4iSCBuauFFXDBDd5QO0ZgeNLzWlmoeZ3Hb9uY7P5Yva+vcDZ31v6sVeuE1zGX6Jq7erypq4nNxUM
xUxjt87srxAb20yso2N5AJfBzn2Q5b47QKDpK9P3SBk/xgesWiZudpORhaWsGYZbvxjZngUCnX0R
myUSRyXf4Yu5a9miulyIzEEw5XUs1my6VVEQrOWO3adkRL3Bm2YHMP3ENeNBTqYZyMuDej2axAMN
pyy/Mnkn8ZJREvJ1y/pNZ92PSBMEE69N5AWtXlNdoV5h7sifSKiDn5p+n1F6sv/0JKp8H02h6EFd
dlcSzytmz820KxukxgsC8kMLYm6lVYubgDoAc9QKkXAP4XMLgYQNPBp+6yfNkXNi+lI1YUVsNgoZ
095tVAvPAT82TYXgxR+poq0AO8dQGE4l05IHFnEVDAOaUzY4xC3i0yIiZ9FYnyeaNaeJ4zNAHXSZ
yj0g2JNgCGyM+m6fzwXInxT4Qny5D9a0oDrHgsptN+i9NwmLhMsdOtT7+ryYotIfBljBoCvWczqf
av9ZpJaWSVYEPWaqdRRHNss0tocJBKiAjQcFyf+EdgTbUDBcSlIvmQoTaxDDk6jhiH7xoe57/yfm
5w3Fjn0PIzok/56aAEEOcoGhC4hmznmjtSyebNOQDQ3l4LRywFztQgp8XlGajhpEPm012O+XhUfK
pr+I2Yi0zvQGVPnA/Qqgxyn+y0oAVo2epAgR+4dIZdp+/gx4cUmUCHgOB0qn2eolOyEhtNaaIunY
eSVOQ0cjPGE0YFFANRQQocLIcYzXWMrlvpoE0MqDZ2YtAL0iwGtX65XmO/icS+oH32VYoXQyhe9E
/kihrmjqHEY1Ifxn0H0K3JpaM6YsFcHcxCxu57baC7pspmHU+TtAgfIPZa60Op1GogWxfSNNjIDy
Yup8mMUrAeep8jeQUb1k1NUav5oHrTbh7N2DKqHw9Qd4ABgt98yagEg7X5ME1+WSCQxSTffQj8H+
XPZS14rhDApZ0cFd0tmQYkiXcD8xKOLRhJZQ/vcT2zrSSUu9e1OCPS/vtAuHQ/Vo1dpLdlKMfRGI
eORENMyXwWme8kJJH/mbUsn0m2VcleIEPg5soPJJNqHRt12ufuYF0u8c850nl6+U8VctI8OVvKbz
pkA161C2CIA08/N/r/K8DIx6L+jRGYOt/GtBQz5esRn0og313epHD/uioqb7I1lAZnUVmYbtVUxo
3spxNeZPI/g5mT/H1+bgZk/YO68X2YTVLc8iZ8iC4L6TkwCYh6fdl5+xcSfTlhdKi5HHotWnuiNp
tTr620ko6lsWArxVTcEcnCLyBa8xSc2iQfBL2Xj7AJkI49sDIkFEgxKZN2oMI9jqJV5gevv/4G/X
7Um4wPHy6ippIK8/IYf2jRmLQzvzLtzoX8ZPnjE1vG3njgO03fhMx2KEdT+96lTvlFSzdburZsx7
+e84FU/wds24XTltHaj5tofGD5/8zblyjOaHKD3GTXUhJ0FrJcOZUmQiy09WedhhlnC/bJKu0+60
ldz63HHMUNGZqONEc0EUzoysdzkVsZFtyXgKSxuQutEq/5hlThPPAqPBoJ1hvpe/NoRJhcVBe654
o+m66KTAPra/LRQRC0+E3eNI5OR6Pt8wczOJ7ojWDfWaKQ1XcgGeV12f2vm7kLVz5GPJc8IMVu3G
hyUwoZ2HqjWK+g8gk277jq+PLcHAOpgH/gSzMz7qfyvJekpttjdVcIp4j8x/rDGsuAktYUdg7OtE
OgPCZr22TZrt50KUXQd4jZ+6XlkJEvB09DVESBhANQ0JA1F84mCWWy8TyTcUFa8fQn11KuV7o2Uv
rPrG4EUEu3NmcBE3TCtZ1nW303laMoiHP566g0HaUvPI412mR6FdiqeAXXy+PWX5tESs/+PqNIqx
mLute/oNEMjEYwIgVgonuEN3XSd6J+DTP0LUaD6vNqmfgnTMHNI8lTsUbb81C/XcHdLN55MyLScW
Cb6ivGp706LA1CmwPWCQ0EZWMLSM2n6dsRI2IkDEy+akNTY+d0m28hLW4rdJB3BXVORzbD9l2FPV
IwCHyLhtyamZn8YFr/1dY3ekhgfYet8xqPZK8dt6MEN6xObWZIpH+b3/jhVqBOI4yUVzdGVk4fE3
I4fiRtL+o58csRbcat3tXM+Ssp+IohdexlntNt73KWfKBepwbyBTB7iVI2e7hai3Alv3uWNG5uRc
t8pkraqvD3CEHqORjM+dCRhwwdX8PAP/rHGp4zTZ1g0pQjwA+Ns7Kte5QUZgSxxipZDJ9DQNJT/D
b8NASsRsm38Rs9POZPBT+GaOkPAnsgrdjN4epls5E7T+ewnYu0WAubyCKvPscqr1C8vGs7X0/70L
OdWQFM0ba6q+I2yyAYuxuNEFyDjV4n7XLSXzplirZvkYYKxLEtZcA9tstoueicNel7BH74eWgWUd
FrfObDFycWdEcdP4DFZc850n+i3B19+Yuw4tmgzH2AV59IgUq+JR7eR4/XX++3FOKubDFu3ELQK7
G8DOVmHcWhvY1nzAdm4Z1oYTSHOnsRfM9VpdzTVCx/QWeVtiG2fzuz5rC55bYp7B83q1M0/6XVME
0mZo412ksaThFh0gDcrg8iTcVexVSB5iBwoxLtlFufXZTNH0JWP0fifLmiF/I4yDoFL7amN4h7D0
7CLIF8lBYhNVagx/d/xZP/Wjbi+pYCK8UwtJu+znwBq44FHZqsYZ4iaS34GxFlx1KahoAFaHm0ka
7TzfQX3BzpcJ0g1VcV4AT6eet64QZ3ERHJmCy9Wk/zfCF0HnNTrm2gA0tZA2c4i1IYLuaPlGAq2V
Y67C2boGOsAsRQLnUJWYggGga0vIAhjfKhiBBWtw9SK9/d/Lno8xI3PPkDBvtsXvScBo1R0weAIL
hxN4nvn247Jp4VUI8Uria1sUTsid57A6KtmOpeyWFRTn/me5O3xnK91E730MfFAkes+8OUxrxxfv
Q49TJOtdshvub88k6ZVl3t29ed3s84QunKlECSoAzr4FnRHFZEPUZ+1I1dmyfC1RkbANvFF62GuU
+f6v4qZ2jd86vVbkWh6BkMdz8B5fkaqinhB50CN6nK1qPpNSwJZeos/WD0UixTmNjRxdrSXQhQ2z
hsRDSGn3WQ6CWygb4/SLDrvsWopL+10GuxlRt3ZR2IfbxoatJQjqloRvUgzOTXyG9CcEWT7o4unV
fF0X7sq/GwYCTym3YiGLR/orC4UUHe9jS5Jg4ZxJKeBwFR4ij9R6fUTdngg1PFFkSlCQm5pt93QV
idB8punOEIQSLhjw7Vjw71OXxeE3gGygCTKxAl17LW9Ts4HVbKXnoR2lJUkJgilJ0RJ1V4hND7c5
vz2rfET1bM9laMNeQy1VkrD87TM5Lgn5zKCz3H4B4/SQW2CxK7n+j3TGZIJTJTllBMCatFOFWRwD
SvxY+1qPaBJVZuUTgviv0wg842Nzhr5clmoyBObcTI4uuk0ir3l9TEV6iTRNkYlGf+O43mBwEMNy
xS45998JE1Y6BC3L//sZaNwa0uu3k1A0voaeKNWSYlLnc7xt+taT7z4LIOkGGaS0V5raRBiwhyqv
iB8pXJEKcSs5tyX07ANL1mo/x2BZSIf2YIG+O98kGI0I4KkiNol5A8XW15EnU4W+Rta+Q7F82eb2
c58HcEFrfAi3G2aFhEK4FZ97wJ9B7v/110j+pfsizbdZ8VA7Gv8d7lgUlS3PObqm649zWwxWzvQr
nRGDT+LWlRvjMllufyiwYDko1LPORe9gAWGjWF5NCd0inu4tcClc6Lda8nQMYAmBHIs4rnrg0KNG
x49Ef+o7GBT4L1AfaBfFOW37eyBXuzrWKbanvYfBXHn32L0iiHaDzNezj95sR3dVm1HNqLTjgtIZ
HfBxxfItUY34Z8cImwHfIq3sRYRDUeBkb759PYwm+ogbx4J1oRBYOMX1xZun4NPPwstByazQRymG
oV+x05wfvt3unxNQUg7ohjazSiNgXjTfshcXTz5ZYs/bUI2y4lLND5udPqsg9efvDorCN1h8gJ0y
/uQWj3yEVMzwNIEWZGMWtlbH48AYXDX235t8cwWDA4Uw++IhwECZV7QEHyqzrjrGRG5LRjpoQuIw
HipytG9FE4hRwEpgMP9x03pjMEPjY5rPaJbWmZ4e7PbMdf703FzAPvo5tamUjjEjA0nkcjS7xA/w
jp2OiktOswDJhnxBqAjHDOlnxvw67g1xhJt4Ac+ZofQsB64tjEMgBz7PC3MIC8OCX0aQlwyPJJ4V
6xYdmbB64SGRd3H7sbIiWBRzRRQQ4LC0rkSVhgYh98x+S5NoIUukO1yh+JZwSBTTbqCqYwZ9hRuY
DP6nGbF9lRObSbenKq3BB0pf1gNqdq24deRE/aqJ9nUeDrvby/dy0EBvBcSn7eKUKAfRhsMLAuzY
3SxIKrtCPZqyvK4oTrOQWprZbut1fXHPv2bXOUv1M8d5WiJ6CgIzC9z6VU8/T0Ojr4SkJ/2oI10g
jauLaPAsmQwgRf8Wu6Bq28S4L0PegqEVdSLyQ9zfDvweMXaEwlw+PpTNSMcH4V0Hzd6EA/Q1fSAw
UAidc93pENVVOBNBf/ujw+0FlYfz3ijuielg2oe5JqmHQkz1tDVq4XIp2riuzgmvAQJgMeRg0BJh
m5z8IvqlH/U1JLe5esEks9K9SdK8jBQqLbJxuR0LFhjG6ve1MQcGyYJa5o8twMDkFtW0ylAfzvQq
B+JzJ64amfk/IpwvpS+0PCBtP2ux/qKHTmASMpP6dm3Vz9CJmVSPw66ynfMDh/aG5Dvt+3dR3Sxt
tZW85sal29DohFU189iDHPJWkABVIlK8reuJV1+x/O9b4dOBj6T1iEqicvqEg8w5Re4R1JnhiK8y
B0/D3fGemp4gtxABVslXPC0+ROq0tNfNwSAly0UEQ7JOYXSa197Co7wdXFdUBFVmv0uzMMtWMThq
yM7Ruf/BN8q3WTEI61MtPp+fL5PcWNfkIoSoTf3Y2lIRyqfpppXEAZkIQ6TrqNRNwpjtPDXFCU0T
l6pDv2J/rvNx0HFJxSg1IRBD2EfKgsW1hz5aTl0mXBNIpLGPw9LaYFQynWOGoprmoDuzOUqjgzc5
zlDOL4X1JKPjvNpicCAHQ7XuWwDm3LMAIjyKGmyWYvi6OjMjQw2GYpdtTsLxclqXx2dsyaX/P1rc
bahek3n6JYgrxlJV6g7YT+imSi9qdcs/dfS+lYoBSYHyNz4N3kTl54Upr9Lbx5cUuED1Q4tsOB/P
o5XEC3NXj/CAIaWgglNpbke1QMuZJFZpjJ8Srwf3kXocvocm/KCd+415N53mtLjZSSc9n2CG8Log
cLFbx2OKFBFFLEvKcGxmojHRhNvppSOb1UNtMq3p2AQM8jyUhPiQTJnHGtPbXFgyHpky7XnEs9Je
QKXEtJcRbterm4JPcUZXjuOi0WAUFf/cO1QrXzV0qi6Ylt77UiYzwCu5zmvUr7FFfpQQrWkW32kb
Ox+OPAOHOAD0UBRMGYVw7xaYWv7aWT8byy3TafAdjtZpucITGEH+rc2h2VgFA4U9FFSkR40Tek8+
nz6iOstIokNEMOr4uocsPqI1qof0kia2iOWqwcMLiJEXQulARmfXakctD5zKUetTa8DuqmhmTYq5
O4rMri32KoGydBB4brSa1GwXFpYtUTWtkkNLN8q4KeFWSnxMWSe6fK5qZULYYS7GkZY8N85K63QO
pf7RNs31WykJG/+BotbCzBBGfXxqX0TlNiurCRGc+Y6aLOq4dIRnve55dvIJcNjiNZKfn1YejAZX
gDrv2giJj5foK1TMLJxg3r3S8sBBq1ZjTLygujRxsj58TnQK8nBBrLsnZ5t4JvT/LTPVnV6wuFQ/
HXi1azGcpET8iDnpBQHo2IfEVnCKX2rgnTJGgaYtOUBdszclTPrGI42/maTWwdZW+uxwX5ka2EHN
A7pgSthOC43yfhOGlGcfNPZ8/aS8XmF2m2EUpwSmaS2sUlj9E9c87SGKUVQahjUKgYPFvb0OUe86
5dfvjaEgaSwdGg/pBLdeYBRu6YSwpAlHbtQEyQlZZR9lnCuYDq6Ra0/kna6NTZ8EAYITnUu0ENpy
XOjh9Y4MWlC3/2HhihZ2aZoP4Pn/EkGejgGvfsOOtDZVqvOfYdJssHrefYK6fHqYgDBVRiTAwKWB
D0pTB9GK2n3pRk/7+ctbL+swVsnU/Mv2FGdza+OkcWNwYpYCFHDNkSNIfKV/2hwxEay8gAy6KJCp
9Zj3PUfv3wSMf9mC7i4uQHjfbyX3WZd9U8qQCe8XU7rd1RsTbPLUcvUk1osp+g5A0EP5S3nqMnAl
FFLVb6whVZL4obeAB95Vtnl3Uxo2xh5gTleWYhGKLA899psBeCCSmLtIezi5Scll3PwJDTt4nRdk
F5FrVmpbtOHLRpyux/bNbb3NBrd2agtPw1RETy+LnsLW0fmE9YxQbHblt+Zklhnp7q1rKOkqxl7S
htGE8s+9J4MRKFYg5rEBicia7ERiKhyMuwV/fcnhNQtrJlLkR59u2A8GvVkV1gqM6hLhhF73dqwr
mJ/xzpmVIimlLDO3bmqa5pU58ZhhoLynqGGIUeK/eW854es6yhWbx2/0hdeTpy5tVM9eQKEb2QK2
16yjkhAeYSQpc/pqPMHs0NXFzxHD9+MWsas9RBMPEafm7oewZ3Oxy0vtE/Te90k8lkNfa5Jnud22
7gEE8+FHKZIk8c/3UF7IhIh8uE9MDIMh8SdUJCn83Xag+WUMBDAq93V+GQG2xzDb2/CEO5NZ+YIN
G7C6tlUOQFtFV3uB5p6Es6VzRcWNk0vkSufxrmNMIwKX/dHgijy4BTksxBI8iH347rkn4IN6CX3E
TSevAjd/Tc3ETZ0jlkQLLCzAKXT1plhdq8WDZrKP8HTJZNFQ7SnQh8DEgNqoZLKX8MCge4HCIBSS
PeXVfGe+qVGUAAe9L28/yD/mC3rVA6CqgHY/zz8d2sDoCmCoyrC8jSe751w1FLhxQIG4txeF3HGe
DsrOmVkl3LcGuyKP2Ki2GGzN88AXa/Fne2UjbYaKOVdq9oISZWX8eaPtwwvoiawo/GvGb2qKZg8O
m6PfpXE1Hjawp7tZ+InZ6hr7JRFP2YtWyvQaeMxd4twRPQXUr0j9f5eajUwwh0NvpASVIU7zVECo
uso8TXgtLFJsWHejc2dJ/ZhIFUGZ1wUyAcoFsX+y9QXrGmVtCzobECOLzEW2XTjiKa1y0jYZ5XVE
9uBPyOKNPANNZ+c46TbZl/qiPBskCJ63A52yxODCR5sDlrFmexkHlPPn7C/YWJuNve2gJDbhhN1x
O0gVYqjoIX4BMAHgkaCr5CU2ItDTAkjFXwN5IhWq21ZrIf5fIwwmf6nfg8zXEyZgOzl0+OANkm1U
Q6/WEvaG8Xqym9DVeEXwL5EQF197C00jZHKgWmcQ9BZ1sN/mvrenjnl0DVHcU/WbU5hDNM8mw0vq
oyJJvBCMZxImkFwiH014f3dJOuaYD2jYnu/5xLd3hOtapzUkcZj2TqbSxRMb6tbRhwBd5MJfFvrr
w+oaLLijpUYabNGC5V7/7A4+GInj6X/pi6notKnONqkr4N2Sn1hnaadHj+heYrFEjuDU46VNBWeF
MhQvF/JMxjii5ZYamQpVVNppN4he9Q/JLE6oG7jcALNcBsHcXCj7dJyXy8qvq9TYV+DrqDvlfudV
HNznxJ3AeSMFVxCvKyfSciYN58bJO/0C4dLm7UdeGSYJqwo8Z4BEG3Z3sP+vnaofDRPuI2K4L4sU
D9c1dfhMOuINPMYwwWQytb4LqibQXhgIbVQ79dQhRy0V6t1eIzHGo3cCIK+WMX1UCExxXnW72kio
FYOeJmre+qtdV3gLdwsGZuSE+w9nYgn6wpDYfYZ4JlLMDiIGpO0zBL50fkiZYhMqxNTqvL0Oupjh
ULeF9xTNGEWJ+OjwK+b7z5cgoHgJd+K2Oly0ctReF5N8Yx9OUKPUIN2r/pxhLffHA+Y/d6QaAFtw
xyhfHj4WYnYDEMPIYpLjWjKQ9Ft8/nF90utRj3isiqwXwBXF1mkNQeF4gSLiGiwvX/VZUcYVUkiS
9BoA8dK7+ypdhbKb+E6h5w0akJfSJEQqEYSt51opEw+SSxe7JhqVm9sOcBmnWUra8zZBJM0ZCSMt
+d3yJykBZZrB/r4LotJ2D9py9xRjiqIhN0e7XWRIXT7gL3ko9MkdaLVGpCQhxTzAonZyyqdzMq1O
88grjE8WE5MG1yoIkemFl93m+/bcjndS9rF/jRf/YGehfeoLlud52MJ9U+Ve9v7igThuUbXUmA+/
R6phbvJ4EZbmpurLJN9b9dgPlGbvCjiK84N7wT34uTl1BMgiHGAA0wO7hzoVGHasQZhhue3Ri9GR
JGd7TkVGiJeQP5K83PWyzsgNN0+h48F5caNTJCsC4UOgyFIujpbJ7zp2tr2sNXoFIS57uPtFcE8n
PuJNEymdY1QxwJKORB3ffmWeaRGXdeJFp+DixCnQSiVNhi0MOP6i+/Sk/MLoZH1qBfmjZ3s62tfV
vZMMt6MwYsSgcLOm7zDq1EIwUTdTCmLkG+VemJwg0nljwfhW5R1eZGKkkUJyUhgodMNzMM0EAfcR
l0A+2ld+KQsBqhAOKFo4m5N1+miLxqXhQQegBSvgfM1wW+HYigEU0orKJZyr6h8p3zdVegefLNUu
Jw+YuF2ducZVGlsmHJUpsyFyWdWvzMqEUXlubtojvCRaKv7V+fgHFpc5BJhnbg+umZn5pqgQ0Y+x
DiB4lQiFEXDK7XPch7Q657gL1su7FHiIMKeCamSWhOBgeSTKhezgz6Ah24Yv6w4kbSxbnR/pJzzK
9Lu2pGuK8JQwEZgKGRznc89iE75menqAwRuFTPFKcx4f6fQ6MsvuH8t53RrdLiBjP3mCcZPemyIY
7dxXhJA44WXubfE7iAiZrKzTebD+HyMmaGxtf0MEwuV7ywxs9cOfB1SRSaq5pBCHbU2L7gnU3DYq
A+YWO11il02zjzsmLARDc30l1JuiyPLYHA2lZvNbMk946v4DaQvwDlSFdE4NzOJwbqTWSJDODWct
Ay2Mk0RXgII08xh7YzFHCvj4xHiJ7qc98Ia3s+a/+0Oz/fIXpDeszE7HW7ZfEamMlF898TfvM1sw
RBiGCWZLUKdoq5MkKbnh5IBK3Hy4fD0vcndWvwEgJ2+N/TTlBE/0wapavGGbQGD8xKs7SAOztqZZ
ohh5CDod9CmmSD3vxSYaqVvY6Yw+JZsNutGV+rNtdSiLhBDu+lwbRgAlWPo+aKWBa8SjcydKPxWe
Q2nSSp7kUXey3G3c8d+RSirgkKHclrG1q+ZfvHNJCaU3MD1gU4aS34sLmuH11tQrspMmLHIrcnus
lRBEXKyFtuPJ1fRxasp+PqQQXdgCWICpPHLZalC70J9QakwlC4F551HyqdfFG4v94lqUIuHotD1h
Tseum/LOa4NkOowBduuFx72K57FOf5BREKIuKgX2IYSky89xSRKkFQJeh/rDklZLmlz1NdGh4Y3d
eIdGvtaR0+E4VS74yjvCmSmO+idpauxPRZf1ehYS4r9oQWPKMpTGVzoFBeBFZoybK7gv2BseSvZD
wSo4npINFmvAsf0T6OAvwNgYYlP2L78x/potnhu+gqLztFiCWGrmyAoZS6v1Wp8oyfaqkBC1AVcS
lCtrfroYd2Qf/S2wlBOf7zB7/w5WNyITnwET7Q1oYZ7XKrp4H/B+E8kRN6WhOJSpvaYKdER8v1FL
mU8ZafobbaJ5I7FDVtPyDedW1xQArbQmS6yXTripAOHZhCQMtiUdDV6fuBx0krrh53awnHnWcSDG
QFtvdlC5XS29YD4iw823c6Z6ZuKwSCtnNgqs6IrLMIwGktpcJ7HvivaEuDUQ/Fl7xbvJP78LUO8L
euR4Cmo3SzikG736K4ytr3kR9ENv7hCpAdBuWVIEw7jMoNRplRUB2S54OCqbi1fPfly/AizD4QCg
VvYBzjncJCsaO2G3INT98qOAlExjYsmlk87fy+kF5x6lBo1EaynIlI1OGPXgIY8tst41ZyFYHfQz
othMCAzqpD3LYGJC8xuer1svr5tbKX1ewPoFn9FBPAxxsuC0/kUkBOgyEyMt5cL6vIf4U0hADHBW
6W3j5IuOlJOKVTVSjUfN/BLNFb++lDfyhFdrzD5xebTb3ip2YAtAmYhQotdUCV9H4RQgdP37BKnp
M1Q4u/9hcOjQxPGCTPKg9TOyCRNmWiUP8jJVelx3ZLa1SJ3rxz431/2kqgIJBjZjIaIlhucYDeqn
6dxYKVcuqyZHapbWmc+LucFe+wBGmy+2nIo/niD1BEhmOEJfE7Xme/MzNPiZ5mdDtoGaw7lcyqmN
v0cwOd3kqAb37b/NOYKFyixgVEFfjo45ZQCFnzQUAFn5Q57xhGirQZy8s3+Bl5jSHb/q8VvAnsCC
MXbjKQknXEkHUxZ8CgqO3iUzBJoA1AezaHMPVBwRVooHC6I8KJRUR/SaP/NPd3U03xzdmE3oDY2c
oV8hN9q9uEihpKfjxjqeMG7V0tWIiusFGu6p6V5PEmB2E5Ri+cqGQNqPNipDwfSMYHXkbB/kyJZ4
YMhdgZR/GrZmGnXf4H1EP5X+HJkpdvfmml6Ysw2IBzpIoSOqD+igU0r9usaT478zWorM4+/TxZ3B
d2Bfd4IODOR+PQAvPqEnTHYikvAznrfnYjs7tsaTKkCuw9HuoHAASR56KPujq9yHmZ2Q+UTnfdxk
aYZIOlRLoFrBET0TQhxgTiWpTd9Sw0gjbh9748RRZinilw3hZVyJlCu4wcDlutMv/BiuvKCriY2k
QZ/Swxpt6F9BRBry00UBfKBIPPBgSguYykTArQPOsIbDCMd78GWYzsFMsNAbighlj1DFIPS8DAYy
TDlcJAVfclJyucNidMIvyJDlq6U+KK53wpZjE0TW9zGxyWwTbJrxj1uQ6kHuawFavJtVX4y4C92K
kbvXfQETf8wjzUk6V0nP9IYM8+bhVTo4bVdro34hYfGlxd526/T7kr8QQvbMJ95TdkoQ2pSx88hG
qY3UDQn7nqE4U5NzfROdzdl1rQN5nWFG/w1qrNfEmlbkW3GzJhpdlW8Yq7J93aClKrvRN11Sdmq7
guA4e3/bvDS6KX+LO30IE/C/eUFIVKUzavXXvFPSR4Yot34ZXLdJpql0hW0bUrcXl0kWNqC0U6jC
Rhz1cnwv4gcB3s+QW6mkrz2PP52vO+EOZ9M8igl149B8McQdGK/R5HtpUyFrgK9EUvZzuvuWrTX9
XOWRWHbYIuwdZPc2C5q17MXo7UcU612xL4VBQschkHnBPjvj4UjCMv6LyEuK0atiasz7crZdk7zW
GL8SNN0bksD9j9p0y7ugUHNRR98dvKkkSW0ZUyW92fujKHhH3ZCpzcxdJMG2r7Vv7kb4jlu4es/o
lYrBizAnsTICOJSgK4WjLyJWH63K4Dde4xLjQW4+5EbyoUNuVW6DSoYZFyobf08T4t/NocssAWvx
1lvEYjGmVMyse3+pJttiTpyijVBdC3uNkQVbQyFYY7NKuJfv5O3fhHDjtaLEjrcAjmEaoPnbltFF
w0XI6LfYDMjQ3S5SotjQw0WBUM0sq1WPpZqnmxPPPcOH95hnyC0v81fuIf5PegXsOz2UdVOo5eiX
IeQIvfXD59PNjSczgYCUNhEQ12nZ6TKdld/hAhia2LH8xUWfOJPFAR17nKX3TPwMkPFB2Maa5n7W
OAmlM+det+Z//h4VkoejA09ABxKOtb5ZjA+XxJ6Mg/rlTr9hwhCBW7xxns5vZ1ZMI89qfPVLFjA3
WlhhdBRTer8YcaJZZLe44wJDx9IwBkxzVhE/J4Esb4vUiR5lWZqnm9omb2joe+COhpCAxHqac97j
V0SmpHqlrSU5pIy45ExMLln+xn9egMxtZWkwqHdbZB6jwGJ3XT8IcilRcA/urlAzHBQepNP2aNyE
a4jtB7vvoh/yobFU2d9/lbSJ2zTivJ9R0FdApDAPh0OogYnkLRm3QIVogtNG8uDyOp/xNIS9Jp7V
F9nBFd97EiHNKouFR50vQP7+vpQGtCoiU3o+/2lrcH6KcQ04QXJBS0Rfm+MqO8aHVakEZ6A0sA1L
0ZLbAmWM8KlR8qXxw2hzYAzRhyAQ1sbgNb/PMhU3eZXswvpaIs7J6rB+qOBdy7JwCUFszcn1bEA3
jBrI0fSFccxQ/9EeZ3QL3w/2sA+m4r8gGUlgddFEGCgZQcWzkbhuCmmxWoNyPFNg1QGct2rMuFaD
rRpbkZyuWBri/8OqhfoVrvbM2ATtJHpXNV2zXDlc/uow+ZpSY/ZmMe3xHZCIdLDL02VEQduYkD1s
wU2rEAJyZDLGcAA0OtKZIN8vz1fgxRTgY3gcuwYeSlbpGVFBbZjGyk1u/AMDK4sUSRyeUPfnppZ3
LJOYZ5u2TdylxAqb4vFoHDFDFR5Ng0a750syZFuPHrqYUd5HNU6uJJx0ak4Cr0DW05sfeRa5LU9F
pkE1FeSScSLoYxjgIUMvtZc7T0v5aSaPIRw+fNKUuvv0alvnwXq6mvwrGu3m9BuzOqb/YkgxRa2B
iWlQYNd408lwVT1jHzqSkkXAFXZqDdkvXxaxrGH+gPh6m3sWz6wQhF0dxpdHO2SQyRjxJWTB5nOZ
/Wa2bzyy5+UFPJSKc7lJyzPE+RX5RV58b3RfYSEGtOh4V6sQJ76tglWytkAvDthzh9YahtZS+hHl
fZzJVKBY4qzQY0oOJx/iXnVXmSwA6+XlriRoHr1JJ5eDLSI5GyOPiZiT0+PfJt4ZkM19Bqj+XMHD
rBJxYZLfuCZA0dQctEJYvZ6PKuSnTY8n19XY97TzC66NKmgTVDpwjLehFcpCSgR6AyIWQwoGELfL
R+FJQ4uzhHMToQ9R7BnYpINPVvRb4Vg9g1f+EeFUrnhRs6fLa8va357IoCBjvWhNVpF/djs8LlQv
V93LfFxXKvbPGl+4o7ifTAJlvzKw7xaNksmhraYNOjYFTr+6NXMoODXnMZgzoT0zERKUYd5RM4I+
AYa1CQYKZpzn96LLCOw8jiVxyM60+uAv92fd9ND1zS4bAwFc4MymosIkiopQ+M62avycgHcX4lTK
B3RUuUVrsDJh+1fK+hgcvB6ucajTX+3SHhB0onFuy3oHfnpO5I+6B/8JrT5WgBM6d88o7vdCJaGc
dh0b3XZbx2FZ96nmxh5LJ7ysxWIh72O6Jj0UO6/hlw0ccu8krW3R2LhGiPp/cy/HgpdWhom5Sqr/
JBk98flJQsOKgTIdRjO3Y9eSEOV9CVPTCd/plLLUc96ahyjCbjjvtHL/+cHkei6J2dDZGEDm30lj
fbXrGNkR91WEFUfjo9pBmxfUvJzB3l8UW3bZmTbjJ7Zl8SW7W0P2H9EOCAniQnm9ATORou+IMaL3
RMT3QrafLx2ADHMzeLuNqtoM7M5kcLIGuISBSQzhXLIszXDYDgNoABPu9BkB2Wy/EosRTzzZeF71
zKFOpxR7Ags3cYOYe06tAVr244rcKoPrzqmOR5nXzeyK3gNCCMGqvZo2zoyBlFcGZsxLOKTTwlT+
0oq1LtLefZsVurdknOlmbCN6GoHtRdZ+Rs/vmAbvjd1qkd6Qvyp6fF/ngrJ9PudmjpeOVPZztutV
Rhaz/fi/9mIDWgBUcouQ0V8jloJF7Hco9d7htfLErVFo7M+E5OGfM+QKPvK0B8uywuV0XorVXuQa
2I+s7/RH4q7dwxI71LGu044RTIq6rjlBBgq/2RaIISQz6Fa5YRG8tlII9a4we8X59B5fdeHkVo6L
KkqeoDLElA5KVdT72Hcy7Djngv5+a1xLyEZBo8jFmVBPda5g/oaOVVSNG9Rl7ORV53J70L/HEaOl
30qgThhDV0L7gGDgEq8myao+X6UCD7c4MXPdDshVBYfeWyDF3ijHOTgvx/wYQSdJzJuyyDc8sN0R
5Vi+taaDoF+ilXjPhjtmTtgxQp/cxxLG2IMPl8KU74ePOEG7dA2ILiAYGTGypsaYBUQbc1JkZWD7
LPiTZO8qk9T7a2DgeDahdlmZ4YLDbJRGUJ/alx078H2enK/NhRmdRO57Aia7Lp3jRyoFBATlLUM5
Kbw28yvggQRWicHcGjCt36zZSV7ApAtrmYT/ufxZUvdQ1hzzZPMoDD2RvLhFv/kmII8+w7AUrNvD
aYhYQLEjeUxhbtq07vnNy8raIRhRaGM9WHQuPnyxADwk7Dpg2Fq8bLioXLgYU3sNB+5PCpR2tKKb
r9EgExo2jv3pU61bqPc6L4DIOZBG1rVA3iCGxGEtvWAxPxtBvS/AnYVinUkGz1oO2ZoAwlHSrCzs
seuS46meY5wu+6Z25/dVLkZobp9VvZah6O19+NB6Pn57SnX92/AXV9A/LuOqN80B7I97y/W0bIaz
SKuw2XK2ZBieTV5OJBq/uTEnB0oRlmLShcWWRGnCxNsoLkGrY38jvkbRN6Eb4akLGsAKeU6Uyj+e
+X5tJJ8MZ34Pxaa0k+KSr7TlQ33Ebx2igWqJF0R0/8FTQhrWaPcNosEMGhVp8NKyMaKeBebVDJw5
Ahy6hMju+wUtIlUuevT+lodpmg89ZEkGz1yFCW1M5K0BV4YWzYNSynavSI1kqoleCgdYbNwpFk9r
LCHThtU6Zg1oVkObhOClDNT8HntSVK1IUzp+lcAWnWa5XZEBtaB7TlH1KMpXETI2rcZdHaDvzk2w
pO9uEIb9pbLLcB0n2tmkyvCOu7XhHCvl1GR3vakwR2okOfWrGpOiOpK8QEzFMNvvGklLgvNOkc9F
+32hl2F0TnitbpGAQIDrkyCZ8FO29i1SxPRK08IZ5VKugWvpSYp9OBZnSS4743ZZDuLaO0kOKbo0
DL1zg5U2aQ/pzad/oGCA037EKAOhDthXSk722DtXfzGH30ggzaqApoLBw4Z0KlED0Wa8WKz6K3dI
ykPe3aeE/SdTPmQPOeeFHrqC2PkQXqJGhxffJ7/rqwlZ4yyBtEjimps4BIB87+2yzjS9jKETXoyr
wSwM0Y2zjBzkBTxGWPEbD6th7Ig3ZBsbXge0qItR3OQobWwnC5luelhRFQdymn29fO0pOHGnng9U
e2DR4DsMoQ6qYPI/3ovszOD+bD8RmFZld3dbJ77gFKp3CqujM+Ou7cDcgxgt/Xm31+mAY9aC0jGC
w4ELo1K9YZUvTb3Wz6Jdd3XuVCiRPgMnj2Z9hOaDLh2gpoQM2zKPMc8/ZR9G/4i8Lek9J+ouOveL
R/XlZWxcxlIdhzjdzyJMbqAN83RGQO9nIZQOe6RSvwy+Ap1EtdifmSSL0NjZs0yqp3ShZLjyF0lo
O+GzHJsyK/aQBlMvY+6OVvNfdoJ3pJBGvVDDZIGhIbZZQUl6eyo/bcVkmtujW5ELb+varGdxm23E
B4cSSeAqJRj/HtR81ZkFCWcOsC4f86zkFrt6bQy60bc/e6TI3bcZvWaiXXpX1x3eRMWLXUN+rfGd
choRILpLYANKZQK1dd268rCyVsqU90pNoinI8cjGZetS1IGsGp2FYKe4s2CVRdBkuWsnN0dI8GXw
2CbIq3D+MvE7sSIw4uKpcBPZnShG17psDSQ21GgGI0rmA3B6Pc2agAIYXU0ueuRDKvzmVf6rep+j
NG+jMe4g0Knm7B6bE9k5IhmpLIkQIg5GUbMJ+riYrtE6o/4TuL0/cThiVKqymKHOHcKclwZjsrKY
Ftz4EzwAxK/koRBbdEgLQtx+xI/Bhh5W2codbbPRzE4EzS+GldEkytB8ZVaIYqhfoK/UrJQ0CWKN
PGvg4HNm0O96FfR6YIVhe9o3l5XlwuhwVgRc/dwMZgVE3i1F3Wce983tCpcBE+egTshbF7T/wGiv
wu+8dJqUCrTp+mqvNKmjLQe5ffbGzt3828ai9mMmms0MaVg+ZmxdZh/A2+qkQ4Yj6C2XH2oB9uij
fTWatnX0xNz8YZXxj6TXom1LeB8WGX7bw1+2FmXkDl4KvN8+qnIEFLpAWoz57Vg39xM9OMPk/kCC
g997MhV+i4qO+pU4G/OoHfneXrIwnas3PF62nL1zgGycGwM5PqtT2I5Hp9BlQgkCm07pJrRuLxIK
C1FpMk2ULDmJvPcE2VZq/4cDEm84tDuTxUhoL6oczYb27hKcT6GCnJ599gPTgiB+T2HY0RGpuZKy
3s2mH/Jw5dRYKhDT3Y3PGBoiJIDW2LOfckU1zaLNWW+zIN/2uPH9J40bMPhYe1XTsWWSTh27l8Xs
olQn1DcdWHV9wD08yToWG28y9XmRtz5SG6K1UrSXBNRdZ/ss+3qN3PLKuI/Az3WO7sIrWNmbeNnn
qVnOedJtz9ld37CCicCXlrs6L3Yefh3mUn7bgKIDUd3NZc0BdXEIkGO9u2xkXbmP0IxgzpgF9Uqc
oj83BXWJXBRv7jqPsoqZiaATVRSDqmUNRcfBA5k4tIPLBpakBVagK2E3oZHrj6eTn5xcRAwV0FSo
idI6TiPzVcGGFdZSlkvDE9FV4BJelXzs03biRhJNSwXT2ll2ae7ppwHifiPNRM+0Zn+6L9OpjWo4
ocOKABbIBdOY8AAQGk16F7T3STnqBAG0ZSn+8HVPcRMWCyYfW1S+6zTXrdOHik18Yd9RWF2fzVbn
xrv/jsO4tSHh7vLVGct6D4uvFfaHP43chwWpDsMt6kRYukzOfz60tWncdhI0L+vS4MHH1QdH0k+z
J5K+a3Jp/Wrfe01Xne74rSdkbJVsSk6zWgflKx9dmXc3A8TTnTcikHO0+ucV/IpAARJpJTIaOhX7
tzTqQwNRLPPWkF/G+ZV6Xrn0OZbd/CU9xKkKJiTkKNuAH8Vufc5FJJF7x2Yah3OE/SVIjypCmLXo
2qJ8oeo01R6D8usNqTQLh2OUYzxIY8/nj4jlqtdvUkg98GEhy2hTlRfoLdp/uHLUriOzULEyuEim
1XJfhRYSJgif47GM5gbvwc3pAAbf9XZXNxJ+LqNCy1+cppOV/rHrYf2rje3AGjs6IQDPZlUt5Bre
7gIseI5QBph6/2XrNYGR3FK36QEexhijhGLOjZ4RbmOfBJ9/GZ/lBZildoSReDMzNzL+bF2JzLRQ
2hfvdiVFSza+8GGXux/P/04sOjCW1ISSnq+jbQuntqtZUmp2Y9ZeQipIzl5L/ep1iQ8SJw7HLsmt
H3g1xo/SBqRXg4L4B2gdU1xx+2tM5XAMoIvHBrlRAFw9ruSSSfaFXEQc/nzHl0pLmT+HrvBWCB32
+07dTpA4+rZUKo1gC6MLK82iIdZ5QHp1mY4JM20Us9Ge5Fiesz6/jXvgZm65JTGLt7p+4Yo3SZhn
NCIyBZCCvOB4HqYxZEBSmsPn00qNPN3CLJElNCFW86HCas7sazOYCoeDRQkX0EzTJFMhVEi9d5Bk
Xv35BjRFz0fPerm5bLQsGVQDzkW4hC9JtiFui0UDUFPpjah9yKyH+z8oeUSavjF7LI+WcVGuoYa+
ufYBrntbKdA24rMOPi3fXJ99wEKxipCcChdCDI5G+D5rv4pBvbzra1VaXXSFXvpjHx1TgB01Ai8S
ndjJNAEm46p48OGhEwA1Hh0HgIVvYV1nP4lJGQiKuuSKuyFt1rIkREBp+KCu7cF9O/fvR8ipwEU1
MP/JeEMsmCqgP6YJdImMtgDavhXrQkwSS+Kz9oL/hCbRVci450QJC7dxXSX3ocFJW5qbouPLmQlO
O61Ky+uJDPej89NCdiHyzlKDqUxiAtZzBjvm22RLfOCcltQlBfmUJ3MtHGZK199F7i/q7aeaXpOG
QhuQhFZ1rhoG1UJQ+wzlMI4T/qAJ1UXpyYl17rDKDKoYoaI3nqjvbAMawaYk7LMPTdu9X41HcDwm
HQCVrQmMTKz/IUjtP0u24Zpece2PXsT7GX8f135ZdvHHLOYzbcoy2SbML7n3Yn4qa32lnK0FrtgZ
pRrf2TUvc0mMlrnL8oRPTfn2XQoPysIf8+di3PQbH3G+gG0I/J9mB9VnoGa8oWSqm5yozuvWGj1v
Q/j0iEi8kjFbKAmmEL39lhafG+BeX5Movx6TqprulxK3BhA5W5D26tiFwlzWFludIaZu1XyWtfit
Yw2he+uksE8cAAwuZcNzWUhpoSgXsYHd8Ec7zOsjpqG0pJYUbqbNzbIhAp8ilqkJZSa4EeGlhcsq
7pZSt28yZ1Bvw0DDkZemWWVfzTqMby+Ex1UoYMIDqw1optOltxoMCytJL/mVDjnNkpyyz+/aO57+
CLWxp7Exs6qzVraIf3K/alEjSZSl/1f2djTxvsAJ4SUXAEhgGy3uq1fivPCquHpCJDAFTgqJ4Bbl
tVb1kLQ4T7bAWgxNiuNd8CLr4TPI8IF8HL4sGZ6IKPvH4W03kfDPfuzKxvxiDFaArlZK54LSB2ry
JHwFIZfolQDxHwNYGsOs0ieodLfyNzQfLgU2aqPG4sJTkV7/q93Ild0zXDCgqOlLgqQMGuxrE5eQ
6BgvsdK8jLeY2Q/qGU0HN+eL7Yn/PSNX5LGJHQ9ixAQAp5zjd0TwCZBX3dCtTs78Iyb/UXaWL5rw
QdCNG3+vSCbzvnvqBE+VLirLcUklUoXycPq+LQ+p8Ymr1DM19+BHRG1jY/3j5Is29TepR8A6ufzQ
+wPYweC42FgC4r/c/cOt5Y4a4D7sOVD88++HGShi1/A8wGNox4oQgyl2ZwP5ywyV7y3U3aNUCtDM
20+juFWTbnoNjS0kznHxiui77f04KaPEMvnPgXfoC9kAA025nKpkIvZKb68oq01hjsgNBYJzR/ns
F4uc51X1mI0yGhsAtob+KgL/yggZ6mU/cDXfr+lqS/OosytQKhNaRkP27uHqRjD5vxZ8aoHgQOQ8
6bDFZsznsTmvCZotLLrfmulX/FrwiFufYGhkWV2qe/kknuQKz9vIo+AdpT7tJifrsPsIY9YLkR3d
2jgs/484gkTJPiHIOqVWWOAElcJ01903OeRKqlMu7qmD+8TP2erJ+KqG0ejaq0l/uKi3IsgmXn8G
ODTqwhsq2y66O/PvZ2F4pzNIb2kCYCvly2/tP/BlM1RYhWm5z5luo5YaQGK71gW4a5QlE+IW1jSu
uMJIl9jk7fMZT6YTeVLSpqzDB36k2fu44jAaz15IcwDsHDCMBUHDSgSRvUDbTvGg2Fw5FlzEQ6ys
5MiR+XiX1m9QxaR9aJgdHZKmK/kwKNQ7lHQLMRJfF4do/cc/v6wEGMGbH5XGbNKn3M3yN/R3G6v+
l08L0dyBPUcYofU4LsNKT1bo4dW1cHpuxPOAHHRR4ExY55cNfKpUGuH3wzTEcfLm2a49mdiKsKHB
jjwY/lu/1H7Rd7HhPppZg5U6D1/JfP1IulaMaX+Ad1vxKgElno7I7CgGh4bUwAEabTjdD3m5XiJJ
DdXFNWpCpFOaW+X5xBRq9qQmAechEs+pxrGG4lMwsOc/esDNLplh4HfNYSEccO2gSkdzheSlZb26
gt6r2nYiAACIQJDdgi+Pj0e9S1PB2wUwExbhhrsK1b77O5SJJkqOJ0avXhhQXpNUxzasfHB7jUpw
wjXqHqpz+DQtbzxy79BQy4cb/buabXwSNEzfyrqQKvK/MC/6LXJHNRDshDRw35EuG8j3DyV31scT
Bjh4Ul40sayJpnAnIaAq+x0YtRqrtKgRwgCS2Rar8bTVQ3b3DeoORanVsuU55xyNL86Q9vkAAhVt
v7E1mfFzhYjMs+AY+p7xWG2Vsm/uGY+BuD0T7PB7/TMAvOqxUFkVPAY9uy0MEPaTGspszJVZ4P+D
V6zvdH4EEOWet0l5caesOmVC107S/cSJrXNmDIPev3LluH7EiKp38fLUFtIFSykclrLcYsaq6Ea7
NtTpvP1AfxGBXkth/jSHXsW7favwrNG4h6VvdBk1vBE+/hQ9LiLboE8VErBnFagMDT0VjQn8aDfN
xt72YYnDsE33IhUc7kO5kwx1qvF/qRyXiqgkYMQura4WeJPliLjCqJONMk48ILKnD7nSI89675A1
Srursvn8PxB6++DiFd1Od9qAKaLgfSvc23qAPdsPSnj0JXmHq9r9VED0keY6wIKrCzbadHuJWWTO
HNsefEhnaUPFoYSCDJZlGjT8//87MTwCTXhRvaZxw0phUz+PpPLh5ptMwPLJRr9iJWUyvoAtssLa
M+kPq8s3CyJnG818vcW42HLx72bY8jWIP2CFGOq3+us+FDnMB+btag59TDUJRDmeCPTbbYi0qLom
jTbtGOjCN+HnnR+U2Zh6sXzYZJzEsaZ6ZJZu3nthTqdfLP3LVlvAgUuh+i98gLYFy9TsIcxKnFGR
486xKbh0IqCutrBXqL4Qn3a7gmcx41LPuJ3Sf1xADXToTkI6K4z3UndSKmpDyjQCX8kcPvAIjEl3
71CBIkmP35D0feaUZ/WKli7h2aO4kJlvampVfe04KbmluehhnRDtTyyUP4GUqNqzqSTawyl1WYMI
CwV5bgG/9ztwY09Z/4k+XVyV4a9YOwYPGRKPVwVeP9P6sceojH/En/nH6odyTGFItIM0IeSy2Gjn
ShqEoChmcaVhnYt9qnTmFl8BIp+gKcZWQiXvMJAtHGqGAKrmPy9pmUjONL159hVpSqsKMiTQ1y0U
aHZ+baN6OvWvSNe+/952D4wVfUkXhSO7JAZFKvqQCLmAMuwMzlVNQEoHf9f+R3jU797MBwo/A6ry
R9fa3lk9K3rGg4Tol2t26yfzRjQ9femSm7i5lVuVvKdNKvE+411tvLdILZQ07XRU2a27llUj6AD8
n3DPkv9P8itizHLosC1ibpEeudY7O5dwqCwA/i60C0AP6McxoFcDiaBKy54CG42/IJ1WKIa1qq4Y
uE54jDFnSqyC2QOBm2L+QtT2BSCYyufswBCV2BP67zB0+VgWV7tpmzc74KHLrawNzXt1wBpeds62
BuJpdx/VQrEHKaiiNGBLJ2mN/AH//mav22aRskhjxrd35oTu9glld9LokGNiFeYGKpocwRnUSmEK
y371fMGi5ThjuAV60+xxrZlgXLCUU7ChRk7bRM+pvIXo1tRsPmDNAXxr5XqB81zSWRXpJXECPfCe
D8E/5s5RzyGLgRysyHs4ZltwTktVsxqrWCr4rno5jBnqrV/nNP9Y7K9LO+BizqsTZJNgwV5Wz8r4
OJLuVSDpgAC7AdI9GxUMhZ4cNkiLk5ir27UArzVQW+D48pTY1vG/ByH2pHPFf85hq+sBcKNk0F18
mhoB9Fjgy04d3pY1M8d3WCTToUkbwIW4TTIye2svTy5zRv9CPbq/9p6UUqaOCzFyErtessTAdWsD
8mE1oMO8xkzBt5Ui+EXnYK0zCZpOEG/b6hiJ65HWqM2YLq5fMKFW7iAA3YuBcxMGy2yoCW19v5f2
irymyy7sD21piWb/vRVFs4Ws2RL+hutRqforxFbnRttHWz/rZPHujygE3KET4N+YQD1/zYCM9KkN
Ix4AzPoU6mTVshPw57ug9TosoNPWDL4nhHFjJkz70uoktpf1cMBsNCueORxHANJpZbooWw2r4yzQ
7cI4zjtu2DnuhwBD/QAytnu+6cqiwckzIG3Dy27d8rVzQgDmYvaZ2a3VCEtNjb4jmKtuusTKlp0h
NoR8sgsKw8s7w0Ui1hXW3yI7rkEkYs05D93kFM25MtJDonZWrYPdAuhvKn8ZgVCuLsaACOo7dQLJ
EoXQAvRKCroBUSg/tC7F7m0+F9q0MO8pTovECR7sGUi4pjAV7gBzCCZlvJsmrbxPBXes8DwaBgNP
kmKBCPIYj7EwgicORUR5EqOc5ZcAFIOnpuOUgLhQTd84eTSMKbNtD7LNWHEiADusMhE49UiaqaWd
PaP2w4VEavcggsXkMIvZhdTqZPI62jk/hr0HZHABqaCtMMQG/OnUNkgeEoZ1cSCN29ThUPkpgnR2
8fUdIQb2GW66rLY14xc0I9PPYKE0IpomdPKltrFoIzj7ihfncocnwdHw5vh/fqu4u8yUvdBNZGT6
Zbe+sZpKcdLP6FgNLCoc0iUkDP2VySBLTtzFYABmkSVqFv25MqwLM8iipY6BPGJuD+7n/cYaXKzk
8qRCm6oTHtsIuGBcevlqiX7kX0Hw9L043ZHeAJ0DjEMgdF3+Kz3mkQgDF8S0rIsquCIrXekXfdlN
pTsS60uEtquKjrobdLvEiRAR7MZcpiTIiFvjeYqbeEOZJULYkEqrqm9vcsk07FA4SqfzNx8q2ChX
oT4w4KvWok4wCCjKs+hQC+r7e+VgoyvuJ8silnO7IsKWNc9YKUCIX4PPIz5Bmnls1SPurhpohpyX
PCZ8SsDBYznF9MzilfW74xerCUzVx8uDysXApWCqL8Z4DQKM+rMwk6KgPE+AbO9u9SsfvfGvgNPo
m+8lBn+ry/Ma7ql1czxVtGFToXdPh3d+rRbWEPfn+jvVrVjUT6DxLlI5WkqkDFEFiZSMTt5rXSrr
lLPVzkepyCiNgK2phBcu8dqTih8u1tCkK9ldiaqW4MbDemFbXuslnNd39I83QYwnXhNxTHxI1YFd
ruwkGHmU3o/MkM+AUOPLk1oNGTZTxBtRmTU6yE3UMeYqetXH7RvAuuw/dOxtposkuad9h+BjcINy
3yT4lWL/favQRJPvDwjCs4Te+D1fbH/2Zep5khRrJIi7GYEQU8X2A6JpUfsjIkBOMy2/htnjNPYl
Lymx7iWRcm2tgAs2qSMfTmIwhp83mhAi1VjXGS6eYFtdTGAjtg0T7vU211N02cjZl6gHLgOHFIBK
8tVEgj8ffepGYxVIp3CR4Sc1ICM+xziz+7EGujGB5LpGh1IGHgaAXo+apuzBegxN7zBIQpJeBUlb
hA1dTLNOnnr0N3KZe2p1uUO2DcDZomhkdYuuzbJy8bMc+Wt9ucZEzDQaFT08dDKtrnsQO6nHwkk1
EiyWRHfdgOtcXev9vHPHL1amyluqZM5BOx9wOFUNI6/KTNoGy1eoit69XJLxjTrJe9k0BNcUGziP
upgrhHKxKPZ+IDEA1HJJXHfIS+pXHrmT88IcPNPSKFduGAc6rL+J8wuMgnmVqhvSnWzCcxDgwbCF
4eIXXsx+7DZ1eIMuY301/eHaswZAMly1b+prOv7jdTUHU4v17J7GCu1IJHCZVu1X0veBpfZ0Q6RR
aNEGbHK3vs7bDCbW5QAztx4VhjQ7UoYcse8cyjVKyjZ2Et509+QsKWeRHB79afjFKSrHqlHPs+OF
lW2zGEThpWxO+5KI2eoa5SWuK/5aGg9+TcFuOP6wTeeWodyaOcVm591htNuQifFuHUe/5Cbnc/67
l0r8oMFgEb/5E7ND0Zi3/5S5SlpQKOjEkJcCV2TaJeRhhmpQa6kfhBjmR7Bm4DLi1Mg+MkXu0Q3O
AhCpyrlBsS3BeDJfWJPknQ8Tr7rYyThmiNEJPIuX56izLmHM/yd7mQjNZ7LBGjSThOQtdUDSuJG4
ZNJBesE1gLN11d/ar6bbtBi+9f3qAn9otMiKCOteM5v9TP7u6wvBIyAiHFtqfriKgalhoabvX/ZU
Ipxf6yoA6ttsspNDBuAizojocw0YD8VdpMXW5OsrrWqQyYac+iyBnyXTyx6vEdX3AdeP+fgo/ZYy
UEeP5nyBF2I4ztLm9yiau4AO1qGS6VbAeghy9XhlXiRB43X5eVpdge8H8ONA5Cf6/+6PgEXJl4Mm
78i6+g7GudABOgmO2z1ILqAkbZoZnD70v38raV+b5l9mrkKLQBeLXsPwlWWZ1GJz+o3tULOAbLFF
ShTpy5FJdTe8v9YEylpiSqwG/tl3boWtytmfbAskFyI5t8cjDxnR3eCITiE+PKDaGH4tTgkhcZer
iDh9UEdBLePtbknHmX9HUwK+dnyKRJimVJJzGLydY8wAggerhlf3kwFKxYFg5VwEqu8Q0xQqnW5S
bS3Hl/4xeHB94fVy+hKT7qnqxvTy7p+TP5iu2AqQqc5wJ7CaTSz659zwEm3Boj2VqKmrCSIwwFUu
C/H+YA3NKC4+MMBBKsKcQwb8M+9sOo2jnWrbzSgV2b7FnSpu2DWf38hgCaS64exbVhJ3lMyQaYTk
WlMbNjqXWY/8DUNa6Yqts+7sPROmcnspZ+TojDxP3PtDHzl7RlLTGGgEW0NM56jxxSqi7Ib/YyCZ
sjAJ/zX/2PAAg5ejIHUViBUPuGJ6HfpDV9arl2HtiZrDu6mCdK+EhZd/Vtmh5bFMnJvMhZM3r0ct
2PCmZahQvd7hPyCGkjM28pQ6DdC+dRl5kAUI+/jKbwlranKYHuU2QcLQjvHjq/uNLnILXaiQ+ndD
kIh2uXNedqDLoEqCqYrsT/ozReaLq4HEbG0RwGgnROfrsZK9vnYLho97Xi8Ut3LfInQ1B+dNv9Pe
5ld9tBjMK5RY3ICsAcGA2hsmF6T7sUdPhxnKAObFRUp79QGOs4/OpxLLhTvokbAwklQfTc7n7oN9
x8Xp5XTFEHrR3+ZUSnB0dOnoQ7JoHhLt+C8sG1rw7PPoz0mY0Vi+E1LiI5/0t5o5Use02Cod7EfO
9UAJkXsPmy5klizz0+98H6uuIEC5YtvEBg86YQO6SBIzRqJXYf3PbKt5/Z4VMspqYnca1KP2swry
+CuUkjguf9uwqTdHaDdN6DT+HZTQOMepXpXzinF1itoxUoMm+RGcsyhdErBTbOMyyyKulwixoWuE
aFnco7xVSPFQu5LvwFxRtwrLcvA/M+zy5CAl2eJvs4K6cMtcoJ6mztu6yczN5/HqX1Qs/2rnRaGB
NS5+cJMhjiy2bqNQMsIQmDbWwESGNVs9SRfdZx+eccqzipwgfHcQkfyRb/WZUpVufta/DyqOpDlM
jEhsw9r/LML9DNk88qrvvbpWlBVWpW3bVb+24aUJBXyonokZbEfLP+F8uLKYCC6Y9UFnXcf3JVfd
rUlM2laWXy8GDzEwrqPh+yTwd8wQGFvpQpguZOVqr5kjk5Vxgl6pasjcqpZFspJc1fmBNTaBzjH4
LZ58O4L53jD3XrJNUZ4mF+w0miGUaSbDNowK+AiBfXzl6KebiOcJUk9jANbAnx+T1PA8IQW297B0
opn9ayOhfUtauqoZVFrci59d/dCYLIXGkhPRQOiVHmA8Y5qkkzyVmYhzobF68tX1gDFsF6WZFCmK
RLIVWXiMRjwxesO7BR4yg85/lRiUky5iJcWtpsW+MIa2x1sdP8TPaHDgFrMSgI3euWJ826U9GY/s
/cE+8sD70ATKPiu+g0m3zqhKuy/FFq8n6SLCvxMFNx8XBADTyDtINOZdWvy7huEU2a+Fjy3VOk0i
hVG/UD0goAB1KWNVYewdYzZJqgQE45lunqd82uHyGd0CpCkUupnMkCuc8/mB0NGMrrXnBfBYr/E4
8PZXPCZtoPmecR37ibAwgyKwNdykFMwfmXRh3p8Kri/X7tONXu2sH2uqiht2ksBLfRmzof330hib
NPyuc1vcXrYFZsKW7XFRzMrO46YYipZK7g5uFl1sMLmvVH/QGo52puyj1e8gcox9tFMV5WzSI4kc
4bfGf6NG/P+ne3a1bri+qLMiWYkMAKHafhkBYJ6vq0zisKApKZRSU1gBuZ6hOCnrN3Q/gsC2CgVI
iYtKl2XHdS99mK3xuqLl1vz2kXVriR1r8dguJQCkemQWNYK83xUsckfF8JOmwCkBw3en64EWdLHq
pAb0VThGag7FasmekZ9m7UwbkjCfKSHutBCOeIxP0USISM+lzE4I3UeGN2Efd68lC0fi+AID2qgH
oUrAHusi1TZiuSS+LXNqVDaD423sy6P1WvKhzftQIcr3lK0TaHRkknvNoNtzaef8qZfoOBcAWlQC
1h/ah/e6oeupYQ1ySN0vPKZQR+Nushj9I1vW2J6BwnpODVZRusXeccSZJa2pCJ2j5G8Rv6NFlUiH
iKAH/64Nwsy2l0l93Sil0W3mlzo7PNS2+ADiB0s3DHbbrXU8EDcbEiVlP1GHSu0qdBO2QpvUe7QH
YnPipyUOERveOy1dShEgbbBFou3aaIhu8ilm+rKHgMKwORESmczK/4WSa3kiyITBv578pElgZzhX
EeCDNaQNM/q+fWXU3mgu0apWSAE/uPMw4/7kk+5CIMw720dzGH7IfI16Dzki8DeYvrtCPyE4u253
WAxQQkgWuEIozjhZMx2Ar4X03oj584vhCaO8X8yxNFSa7geZTwSVPIXlXI75FUUGbGj/5QhLuYYP
GzEN6w8c+YZqtY5FSU9+RX4mfZPmhANH5Cl11v5VEBSyoYFzOsRal5IrsZgVLUZGL+FbQRgEaY7C
ZjkQBssFqrgujP1Bp+YmRFzn2+HXdFrV640JBxVytC8w5xSglF8pJcK1qdoQwmyCTFjYLcSMNPM4
q2LoKQ3kH63AuAwBmSqJHtBjHuv1cQoBAbbx4wra/x+pOlY8UlNcRSyKM6eLnC5gUKP4KFodyg/Z
KJYyEdL5r7m3nRQPk4q+QIMUdxRQMYjycqIVVvLQa6YDeecXY33ZiQk6NrT0wFquLyf2iHMeJpNC
VYtm+YVkOxV89vuhm+vkCEWqd1knByZFR3JqD7dv7qVtiVd387iBiMw0I2GsFpEzEDoLqIn+nFG+
mFMutZsOp/WvptCWlsEA1z9qfXUkxXUUI1sEm5pAZyt4gs6PRVdLGCmpSPJWjDVMEDaSBBTnrz9Y
/nhU6HJ7G8yy9XMMEgTv+7DKG+W0HDIcXPMbwdXpQ+SdW39N0U13pBKfwtjcCXVmb8YoXXcWsa1j
M1NyWhYwrn1F0K5BoElEDrmhkRm7+NIQzWFvkMCOefRK61JEYcWjpHLIvfPYYP5qTSIAXk2yytTt
YylW3zDpVG4jOuVhHokwExYUGL1qQPQTkfPr/SQ1OhxooR1yztgTEJZursoLjquDE+/hgziqPcyl
vaAMl0VR74ElMFmDqJNUS9Og0GccBmvnftkzB5GVp56nvIhVeZ8zZDKBtpXZhR0xnjZUnDvZ2Wwp
DsPaAwrSnXLEPu/bARCxmfNHHVBIw6Sjg9lnDRtu1KV2hZfwNpuY3XN3H+LmahLuQi9/oFgvZzpB
CQDanTiIQ8vHvmD4kNofalocY+bm1KT6oaZW5gJMit9sd3RP09PIfkYTWvfocLqUqVCloveqvi+d
m7ckVHzrnIxcMdM6O7igTp1Scc2DXxCjURjuy5dFEP89+ZiNELULvjCEjmJ8gmcPNOeE1A+X3vbd
H/sU+PZmpFmyFGBqTOMus9kaqqqP2LOYjDVWwDsJ/WxqdbJq/EcXuDd0SRXMsyCnqNISXxFnGdNQ
FT+WEkx3axVJm7QBo3f/FSpn2fQ5rCkjIYwJDUyAGUiWgOkJngAkSxUaStw/YfIEr88e7SYpc1/i
RWAUiloEv/wDK5nYbqbe/HEKscxWUIGxbCdnUARrOfgrNraE0f8hU8ceDw3wWc0Oek/ZXyL5susu
Dot5BZevEf7GIJzAu2+z/gN38e2Rj2h48JM5wNRSKFM3CAzeWJi9y5IIozjkZFhNgStdmB1e+bXt
evrqQZzmfUAZhULPgguSWYMFecRPR5kcSKRehqMRixt9TJGzyLfAKb3m9ORKeV71IqW0ps4Wx7El
xXI0vKXgUEy8jruB2xTBN8K7/hR0x9Bjg5UQVTyDIDnezX3AFbxN67ZUwyLCwMqg5p53LF4uU6Oo
RADdzOwpsLTy6Vf3BDmwhjxBinYaCSqATu2tka89j+G0uVQqLbvwsMuWfbl2cFWpAQFqbqcIPBh9
RLwB1O41mVpLk1uhObpvaYfIzsFbVwt3lKa5jnirohXCwQk/sjylJuLqj/9vm9XV15t6hxuaaq/t
8ytlhTq2M/kTPr767I4SiK1kdwnZ78QJKCvgmdM+TK3mNcp2Vam8BIxqE1Q9CyeXPJkFZDKw6rvc
mztthIQqNEsLspEelOp6TX1x1h2BfrfKT7voEQdqd8sUn9YFNClye19D2ZNgVJbuK11DGrzK4udl
44jeaWxsmyamx7hfw+PFxjbC+/+P++r80chx2Ltwj1Ny+C8GUtHnAONuhWCDrNXobXB53JhHRb+4
NX+eJrlD4tNM0MROQupnORHn/aDaB67LjuAVb1fHHXK3dsUkslScwnZTZh2I0gORR/+/jzTt8LxN
3Vt1171X2qIGzMak1FGnhIFEC01ZabWOHy7YhfT9JAd+HpotS8u7exm/lGjgP05N6RbBHZCAfCXq
N3c9rJQOerPW3QNP5BEn+xHhDls35cncmu3TVDt7RRsweMIZNuhl2MBm6ulURDxrS4kFzI0IkpzG
f/VPCZxV79wyDstH/Wf42OfzaF4e9FuKAiHK6i94iWIUhBDfEqE4H83TbtyRgktDPhelO7DivHXm
vr/2A024+jzulxmlstrOg/nxadwM76Jh7DmstfBdvHsVfjKS+LpEEUt24xkzwC4M+Oj3gDNvylus
7hGZq/qJ6PpGESwlmq78yHuL207mb5MYAwEEZATSV7PT014QAaf0xb9UeAIRryBDUqZYLEDObnXD
wwrHlxE0+FlJAJg7IT2CfYuZ6yigB74cedx9E6BP6W2pbH1mv9kVy2qzlTYdcYRAU6lmSPLFEH59
d5ARaOkW0IGfDk9JLFFGKhUgGOig1vSDqPj2vjxWshD2JHgPaUO0NVjIDgqlwq/PDV9aTsSd+0Km
q3C5nSXuLHaLWN/NE8GJauWsEvkp3Iq39fBC+BPaRR4ipuPFgXvuhtSW4bXQ60NVnP3v9Vk97VUj
DlYDvQ0rKCE2Qz3Q3VQI/+NQX4bXG3ahL7FimGd0i0eultsyzsRf2oVCdNMx29TY0/VxuFli/pwz
dRX0PHUzBMTrsMks2vOJ73jD2mEhWypZuwzqTu9Vq5dVSWYBcJFk0YYJvf5C8Hp2tN4MZ4QPa+EM
xEk9wB9rtgvcRrSZPCDNs945zxNSEcXObpdPzAdoZ2eJ9KKcbzXpHt22fdVsTlUiZ1T7jNzbzTn1
3ImQOoGluYnuwkoPKPYPgcoosCuQJJwT7tcS+qVvEfahYZ+m2/JkljXpCY13igrTHcbOU5ytmRzE
UfwURSAXdj3JHwj6EsJNgLu0QiHfXhFCJcaIKS3ACpwLxH42o5LUI1aRk1PnX4doxmbRg9POf1rb
D4iJDbXwEgLFYkhWteSaQhMFLe8SsRWLOf9Xuh2KSJoinpsN2TUJv6/cZPhyJjOxI76Lh24cnIp8
Pp4sBoBwrsQjcFE9+vMTX3TAC6JP7758KljfqG9t8xMUgKzjkfaX7vAi3hAEbI1iEQuPa4g1+MlC
nFd953kOGJertokwS3GhK4TpNF94nDx1Hp1yxCNfo9WpM0h1VK1hi4AXm5hHgoHVJNmzmmGlGHAm
28j6aClCjWLifGWIqOmFgZS/m0Dkzhe8fJ4NNc277uk5F6HoDFXxgdm+XuFbaRfeJdpzf3qTocKG
l0FLkcLXZQLk5D7pcD8TQsVxjy49q/QRDjQpnPdMII2V6d1iIO5UTf7i84XpHApMctk2ESmYfio4
zGAxaNJ3qU+Tq1voyP786qfHa+E6NGTJMULWQKGpLV0UJGxfT80IAlhmMQN3SlyIbNiLvd1kCbj7
SgJ2cz148hIlYXgtVtSS3v4/JFQwXy4zpnAx++TgOiSXE4fP7eTf6aQPDw3gUEQzZlr+VazVf9Dm
86thKwFiFtwZ5ySLKJ2j82soXiQRUim2ktemHxY29mw4CbSG4w88QRqVjg0iV5RiVQhTjLrLWpTW
18NaFSa4rzMRssca5Q9LiiEshlgfFUR9FIdl2f/OcOKxn+4Fd4oeYxgnOThCJP6VrX8s6wLtK91S
voWkRNn++82Gxu78SJblNREPKpBigssrCzbIccE3f/AZ/Wg6s5stqjtTOiXE4hjhcAI1TdTtmdzZ
sr1+bM0/waSHN9KgGXZYPASEccdH8ANKJQkUG/uMNsn0TgORdAlEjjojD0Y05Hwu9c5geCUbR76j
dVRHi3kZ6bYQFetw87wVMAD047ZrOJYxMInrpPKrEhKwAvKS2VDTVH3+vsPJzSR+ba08Bkzrku0o
N/UYfU28RD/giCtVTmTmH9+AyrrJQAzLqUnQdSHQDOFDz8l/4HkrO7NVX188rPzgVtIAwPoIRjlX
oIvAlOoi1V/dqSKlXK0z1IOkDM7JV/+HBd9evUYpYSzSPazb510HubF2br/b8cBhgtVb+P1KxxBQ
H5xw7dhFwv5wLjLv9mVjMet9jo1xvb2Lf1ap2pj/EzmVMuYbRHPJN41m5xL6CKGjxoSX0EPVZv1y
XW4sIYEWNudb/ViOGGEddrVSX5+sZM/6Cj9tSXH+VizSGiRbstg2cHUhuNctAFADktgDOV8MylAa
GkRbwNDMcxi6jcycW5PDcYWIJTWgKdXORd4u1i5/oVs+GaKc8V8J+9To4Y0xU8lqqLv1tjJMyNpp
/piMLzpyk5I1Z0DlZ/o5Rh31VKYLbpVTe+J8FbwE0QYR0l5DBVrR+lBYqZr0mDpzJ9ddknJ9GjfN
d8zZveW09xlZ5fOdSdc5GoSQqUxuCcBJXYAlygIP8pTTO4hlMi43/Uj9GnlviSo2dxAXrlZ5S3TF
W8Wsr0FQPqMUGd/XGux46dO6UbFPRXczaIsviLVv5qfarAutmJmrmoRc5TKbMdasHnWQ2UrVGkuc
EX8k/4+Urr9o+Lbk1FfAVbgREznxk92qG/QoaF7G/bfofkG6m7f2vSbzYO6l8XICqAdWccGHs3ut
WvxYp6VCiVQdWDcYNcoceojNLlcw2A+OA6JaPqxg2r/T9UVkviNeFcJkDnT90tqKKrs2wd7Ntdfq
JGGCDMar6BlHB51Ja4KTZPVPAnmo4Wr7sden79FojqGy1tY8xQuh8UFU3H3BtQIvsGV+ajqeSkV2
e501UFQMY3dDuLCa/F98Fnr9C+dxVi8j84/PwjEcv3LuAq18veEugpmFI9SfvCEFBAQ+nJEkpKs1
sSm0K9VDtl1jcGUctxM5zM7qgg1YHjuRnZTEe8ZpfAbCe9t4PsDyVXYimE9CU0DxUnb0vk4jMCIY
KfELx+Ku72T3ckrH7XBR0M3cK2XYQNGR3YLBdAA/FvzSIOFsAQsK8ihYsdQOso8BwPV8uO40K/q9
vTwbVYt27oomOAfQxJWQ+IZ7J8IlpD5G69iTalL1xeMFudka4p7+kSNHiNtumHZH0ydRyx+QL3iA
FRjMSyHdSCL2eAXqrqqf0GIzCFHNC5JZwIoIYOudzqcD6qfAN3vHpoVD2NT/9qHZiEm8ONX8N/mp
1FQdWALM1p9ZuniwqV46CBI3qSQMWnKFnONvRrWKWHIwYhc1eL7RKywdVsxHhKmjF+JBnVVrbFce
yHABON9+pEDFKDti5rCQgmeLhizUq3VeON2lVz9BQ0wQpQS1sX9iWbSO7uD+zBuvrJMtQazlZKqK
eog/Z8akvBYPcQXO+xdhQF2MpcA+/fEqajqu6AmnO9vF8/Ckx5XBkgW7kAHhnhe0a4agTD4/PMiZ
qEwg0PbZaVMja+TKu3wMYmZUb/kDJPWkhgNF0wi07Va2c05wP10eOSudwmgWW4LVDL5Rso0misni
hYClzhss15BoO/8E3eBJwztvxg1F32q6T9W3LjibstjB7FQ1tdhliwhbKI2erl+Rd8bojxOdVFg1
iubhE8BspGBbomqJ4YSWHGAs7H/Gk49j98eQM792xvh6KXzrjnN/ik5hcG63/MbIEOrQKQ4ec69Y
Uc9JOxZ6QoSOuKyDjjaqlPVYQ5bdjB08hdC9d3IlyH1bJ+D+EAy0U90CtY8TVRIZa32sOau2CREf
T7i44LWHDduvU4mGHYHlEGLm9ngvYyzaZBn+R8lEb3nzrwRzjJKrc1+6MJoNUYw8y990/N62MMAT
gviVdzsOa/vYekUI/aiVVEEfpH+3/Qvu9FQsdZFZjSBPfNgeWfEJuqMwPWa8nNJ6YSabEf7baMu+
MOTT3l0RQPfpnaqMVYP7EEy3Wfw/lQBcjA0NbRu7E4tnnmoUPvY1f5/iUyHe6FBmBai6seBG4byN
Eg+w+dJgSZqTeZIDcPhDRrffollPLq28JFMi6xFewsB46GSmJf5vJ5FZjGnez1bgGSVyFXobEDYx
xyQeKssoa/P3iK3iA4wYDbppwCjLJsPhbalJk02T5YJdzoOjOLnV4NpBM2IcTNArY1b34XBI2IYd
mrHs57iIuwa9biA587q1wwdO71KRR5fSHiZW1u21DbxL3ThusJP7pckIRO0yCPUODMLJuFKY0uPD
8Db/inrCy5cwG2Q8r2mqPutAk//nywhrNXaGPQazAoXqw51sE+/Wa5Rw3+joTB2rlnU2LlMYIdQx
fa079X2gzIlnvs1PJDPTiaf45q9z428uSYlUPa27LrRo0d0zPGJkCkAbqDtHTIv1KZ5pBl6jl2C6
bokz4W+v0IBX49qFzXccj+2cVvnQQn/js8FpwfKKO0GgUzYleqdm0Tu/v1/vAxxzBT5pZqadZEyF
ibdFjsgtXaf2cuBXKsmCKdjUcd5R2HDUmIArTTpwUQ7dDzq5/LYAhnQEqW2f0rHOn6VJWrnhGWLx
lYkBO8kCQTLtai8Lr57NcRa4Q4CCKZuvYadY4mXVTzkAFIBz4l/uMweq3Fx0Cu2AWZqqHhETzJS9
p5/jqXuXd0WSzQIFSgt0ihRQe2aklwETHHhI7/hjcjYTG56u/XN2qAJSHzVxEqlnczNtuH7vioHy
fSBE+a+bEyG+SWBEHyWqdD/9t+06s3lRFyW0A8s+Z4MS5B0/kWUHFvuyepos9k0dP6lvZ1ZASI3D
/N02Z1NpwTLiHTWBhVmOSvmepXni2oEjoWiqd4WHY8yF4Q2UvWySGlxAcI/g5kGiGqoOOk8Hffab
1iAiqvrBvW/QmmqWPc24Y9H0EsjCzgA6ANl4SXzxPXMziHzv78+pWdH9iQdOuW/D2yeNrTG1bK5s
BtEVcUlT0U3tObLMY2WPU8KK25hmgBWyDoYTq1a4vdkUDAsVVvPISEWp6PYTNoZHDnb6U8/qM+Lk
q8XqktP0PfSdygFzGUHrUrNiPqJy8AHiWgXB9uy0It/UJqgroImtg1w1H14nv7iR6FI9PPIlAERv
BArrlsEmGqe1A9RJDjRaiW9Ee6r+X4IuvONHSEan8T3oJfUHr/D6MHCct4lQ6qU5YaVZ+X/r3r31
Lv7mvz78vyNp2SzaEtjLY6kVa8GNLuXpluTNrs8S7ryahufZWZvzVbhLkp2by2urTycK0KcDlHHl
JBhwbXyIMrNZV1aHJgS2eBoMtXtWoAT2gIHGhkt7+zjZNj7PUvj9UAfIkAOA1Pup5c9tsMAz34z8
JzVfEiPZ/IOl3hVy6+9NTJ2jM6rFvlcLUYQAosvmU8oQ+dj7mCaIlUKLJzax8HH9uqo18G4jEpLD
E0NTTWGUV2az+OatyEWLGJBEjPayZNcekK26aqfuK3qY9Jmq2zptwkufzlkIvTaiuQw9X7GilYs8
5BI7+KoCtZSdCfMM/G27OGMRhnUZqd1cQRlkQc9zpj9CzzlKo/6PJxkh6Aq7lCw0WMcHr+nujdKc
fkEpFBJlrtIviPeWX/qg5TFQrSNTEUZyXLvAMI1o3D9IOaLGpY+tCj7/NEUpsdi0PLjoDX9RPmvL
HnY+67QP5YPWRnFumdgEy+r075XLFD4FzrBEvOMo131HUPWIIFTxnqIebZFWNrfaqP6meizO+kOY
rELoEbPdPkBSHCMIXo5VKKx0tR53Ta9q0yJurNLh9WAcKDfaAzuFT4XmDvF9U4jFyZEJKKFoCqyz
0JhRDqPX9+F/OSRBSgC02t9RnDj68mLk3ajc94R3sn4KePnlmj8lxNdGyaoVgyYs2rl0rmPFWmJO
edXy9IBmb82W9uIcBejQoPnOYW57Uq6BuyDRlxxWIuRbQq/Jtt301eAjOEEXISrpu0ZYX04ETdNx
/D5xdZQHxv4caOyHty9WktF+hc2nGwxL2JS5LdWyFJoUjNb7QoTmQXU1UIWIRiiQ60QWGF73oKe7
vliyXv9qdSUcUSAhnCgTDiKoezWrrGDTvcaxWX1+Os5k6k0vZFNhD6aZ0HZ1NAvfUQRv+PmrZ0lb
YpPJFHdkHdXQMQ07Kt1bFo6axkbzircCKM07bxAeXMdAjLQDPxVN2Z8zO/aEkzKGT2sY9MEW3IUw
w6935O2e1wai4NzVll+wd5sYTNG15aZUeYNDoPdzhooZ/nj8dUXhPg5090TUuQA04ewpzxlU/Ri4
kEXMKaEPzRQAndv5jGP1N0LWUFFG7ot35BZOOH7kIjbxvY8J9eXZFiTOB1+augWupmzcqdf7pG7e
4QCiWJ162yfYIoGclu32MK0if996suxTwqrDvp4aVi+Ar6Qjg64JpbWHRRBXYBgJZDJbXQd+mhAb
CXEvOZLXuZXdnJGBpu5hUOCxUY2cSD03nxuUC7jIscrJLztV8puDRuNNXms+qK1Pi9P/3GiYp9cl
wWxPrK7vBItRwGB4TKzCRldPkA8gB00lWKdgZt3gQqYyY9TzuJAmjPgb3fvGNw6sjre6oHPw/QBM
2WtOzlCMJNVVKgmDvwVLX/xiLIRgrpQeQ7D1sUAs945bNad+op6xRLpUMOxMHTVuyjnGkmtvTZsz
hB6Gj2MYX12ug396oHL4IP+gt6+2eMvwZmuH9qvRCeO4bPIFc6mwkDDGWeVFjjNiDfVOvpb2s4ze
UKuxV2AF0SHg1pH9PJkqPqw4TEDof0HapAvba/RXwRAoTy48IUBOKRLyeF4L8srcQLyQXdmNcgrQ
33gGWRcKOtLFvyfdUR9DxEzSa79TsfJ+6N+NxRUIHck2O4X2KwiBLRQtuUc+9Me/wwQYPP1061oX
L+adn5b9qhHYnIYkF55KvLu8QdZgcLf4IT8iCqWB32SrpbqBZPv+f1taUoPR7qYkIGV6HRBWFfYY
VOeEIAXDUBj0DrN4ULroP0O8IIw/GyR82Z1bcqx/68qoQUGZFmTCLzolDrpeKPiLBiO/5Tv65WZP
Q3QEFSOpU28n5ZNoAajbcFQATpRwt6jX6SqbsKQtItr1Mr2USmB0MqlNpDWAI1lSMyLbKSeDE/iU
9L3WILjnEUkMrtlgbMEc63jkCBz0E+9PwRbr1oiA5WkPhEkkDyMns/54fzN3fRT0SkV/am6AMxCc
BxNhUiKHPs9F8R/7WryAx9Zz77AoAMOPy8zlFHo6/254kkTFr4vKQrN7FBpCCLV+WUbT2ISM5md4
uIutkWuhKlARBtWOrc7ixJUIyl9sSFLJcoCqGHiWJxEeRR+k1ZB/zY91quKk0c6Q4cjxEokrgLWu
4/0aB+cxooDG0YHm1MOtmnD2w+M7btQJ/b4zEZEpjBuSE3i58bFxchb46kDPjG15Ip8JDGcD9hQS
AT1QO2eiq9DtaXjX8toSomHdrn/3zCHtHLfKUmRbn9yBG15OO75haOOI8YrnKUKC+NC4K3jNcU8L
rSgTNdA+T0gh+9hl0rm3HBYdp89RC+1UilW/bzCiJkAK8rb5CV+UWL9AIaGHnEFVQm7hAN/AE0Xg
zQh5MDfPILa2Kb0sL9vV9LbLgvknCPV2/p6rRKfIBNVLORjuS3UxicSCqoncesQ9mNvi49CNLOT3
3Ni3CGelRTs2KG9gIGZ4JTM0GzRVzsYgWoeBfZG9q+ozLTJ02U9P9AvBavD8uBSm2swK/FXoPL78
rGIfplRzQt5NAu5t/7Xu9I53UdSPc065QOXSt1Sw4gcgaAzNarYKB54bCqmQKSl07CaaZGsfgZRx
cxIAQs4+EP8E6V7aSvOnmr9YReoC24A7SgT7seLcd6HV2EUv0LZmDNM0PSKBQUP7UFBlBOaP3SqM
S0J8jjTRQOB7jxlPaaoBMuY4bB+BvfoGPqWrFmImRXogrrQQoOPqHy/xsl3CpwZd/az17VVzdAMC
AEIonwt0vJ8imMk0LwTzt3sR8zx8Z3f8zmr74S/KVxY80O+MKUFNFwRBXfJsVP89E6ekn7vpcGmL
FMw+j6lOEc9+zT02dAQZNympYQqNQJzAhX1OuWjpmoiKpBgW6TnswTAQMCeC5Q8dOSnqwJJrqf/d
yTZROptBP7Uih0IY+nm5fWtW7DbI48Wwl9t/X4VYfryy0m4rUwad5gMnUFVg2aIr2SZZ0xcNEvKd
42ztVcNj0ZQodvGSb3De00DQG5J+FXlq5pDyQ0uREN4xhtnKNDMlcQ0qgTAakBPfqc72UBLdNMIf
qseWh7WFrz9CMjt0bWRMETwPrpvLlk9N9T+ARxUwPYJZkkgalMikwL7b+YbiE8JjG3spSJPEmodu
a/nzGYUTdYLuUXVUISZvFAECqHLjo8nN5QejiOD8sdpfAHQHQK6GUpFyrbOtcPucUckgSDQUhSKX
OifQA6P8sswTNYERLZw+tMRapXsG+4e7QeJH3iFHWw4doj4CnKPlwguvt0EyNxoM6K0e5M1wrfeR
iGtWcEDj0Ai8IUextUET6ErxlsYnyAlh/Ur2Qw/e9wk9zAhOl5+7aTt9/wMmLjiJ6fGlOx1yvcaB
jAqjQrbsUD2xnCaasoYbFqCyLtEomdfppesT4dkG8ozZ4EmIPGG2ivBetJCuds9tPLnHYpNlfWbO
l10vE9RdADu/vmDzt3jNbKMfBty738fMw1Ep2tfX7RvXntU6LkE1o+A33wkaZBKmrRutj1x18Uvq
23FgbtyKqTyZ4mlpPrXcnB3/9nNHwTutD3YRS9MZkJkVMwqTxrbGUQCcNO7WOXC66dFSAiKm3FWw
Y1mIV2AJCWpTVX6kBJNYRijNHR+Q+3lcFgnLdSnK28gnwu7WspMSOi3IvwmyayEhUY83ynZAHEYx
djRFctYJFDeN/YOOWdvzNFcQw0KXB+l+uZtxGKSwPCwexgsBGY4BmGYA00YQm/PsZ7M3SGTz+g+J
uhCT+yzTskDNIEU3UiBP074f/ygnpNrWWdhy7KP4/G9sqfHHcNReVRq9vT4wv/oqBdvI6C0jDZlQ
GSV7zlwm8FXtqxxBPazIuUZEY3cMILqhDrwheZZHuyoUL4LGdpiHp7wo8n9WNilaBp00McHZZllD
bMDATRnBRPwC9utWv28N5qly0CWDRnBYo/IssvxxSmuUWAcv0rmgDjlCgp+88PU09tqROLoI9gLD
ggyzzDHC+Kl+k1Xqf/gUxRS9qfnFipeepX9WyhREQm3MxvzBw89rE82kESnf0l8fB3JU82fZwQ7e
xMj/hijqKKgIEDXn5vWiOhVn/aKcQTBRB2s6GI+f7eP4hZejtkmz7WcUb5XcffMwz+iib8EOSDX7
x3GfpjrF45rkchqGNhxjwN3GCyQAZaFewMWXmmG/bs2u7EP4f9n5oAU+3WOB6+gqtKypkIJRCRk1
qITbjPH/GoZU/wq1QKRetBPvQYlMuBR9kRzD5Ew6K21gMuLNOd6mnJv6hJ76m9Zb88bur3JStmYX
Tj/lpD/8zMXO/qsPD+IK/eePqZedKA2NgDF4zKV+XRbHq9TS9utb+BrEV66tIS3rMpCnJ5Ma8N2x
DKilP5rDHUfAY8PJkIR4f5MjXq4s/seDmaY1ypafLJxYE9mCGM45yrP9K03upSzo8zCU4Q00Y3DF
FU9zytUdNhrqEjbc1PRh8n0DY/8jKj2QMsgvwmrxvkX9S1r9gX5+SlJYhKvUe8fGGTRba3bUB8cQ
9PIznZBu8qpT1I8Pt4uedDNeHkSgsL2CtDUHVMMCkCmVcHq7MyedNvsyxN/mFoCl9O3ghzV6jW1T
jJPnu1lk9oaoVzDuLr6GVZL+O2tVkw41q2PFDtCToqD/Q2VZ6Q/YIsGaIxcCuRcrO+T7tWsc7Ipv
FA/2r4TwfpaojdO5oyB/LeTUYdJjnreZ2Re4otZXT0u3bX8pmJyf413y6uFcynlAVchLXTlV73ks
J6/+/9ghkGfex0W7MVElkRFBNfJfY3iecvmn8H1VaYZL3t3ZpGa6IN9sGvVetMN2nIE3mIHuA1nd
sdUEBLKKIZ2dLORydjC5A2kxEupUSEaevvLDmrh/ZSgxtkIY0sARIHQzIZnXyUoJFMJKyn4t+7qL
V0Ogsz1pEgjtAEAzEmCUSTZ24/G+LfR4vc4Uj8W9YM4ulMmeVxzUDafPf7jjoCbM/0RV17PFM2QB
uO14lEEu419uxHW2zS8PY6OnroCXGVQFPh3Hq2y5zb8YRPoY2dOXgzXi9zIEqPUc+SWKeL6tCfQx
0tjZN38Rft23qKVSH2hy9p6RcOs+hL/aj/tXRIMO1uN3WOB/hAADluQGsUHSjo8GjsYILgQUC8Yn
x1cbvbEARnSdef40TxwBowSLfS4TSaMd9DlBwh8wAWsPqcACBo1b47kt3fm18C6AZ1YIi00zZPaZ
KCl29m555Qu9YYBKC/ROcm2c8GWjnmSaeJ+IHbPl0Us7cCO762S7WexMmGJQI2MbGRxRGoi5XPfT
z6OW9LCIML2dbsSWOwq/MSwHEM0RvNLNMaUrty8iN9NhN8mO/CR8E4OQ0olvlxsQzBsfjbjYXy1X
Ub4DJU+WSOQNQLOqTiiogVHeAI3rzv5JOLIJoSFDtHvAUB+pkf1MmEnyQYy4oa9rLHHdTrIix9kF
bUTeqFMq0+SSvbWNadTryF8xf+5jWlA8eVQ4KFoY4O0jM7VCkWQUkVqLpapYdBzrj/dVOPeHOMoH
QUz63hkqQsXip6D5eppwGhRziyxxJhtcdhyWYXECoHh1NVp4N0JjVR63im41mhXXbd6YqLdk9mnL
vrxyWKNpVfKCdcAXelC25VR9p9jSD09qceQA5XbOHfIgFaaJifp3MyidLHh/WqJU4ng055cKLji4
QHBgJ90xxeCmQIEpzJz0BKH1Tj/cJGey/eai3BvoUmimQaC0mJy2Dsuv/omzsJzNqM/hL7yGpykc
CPPudlGvQ4XTIJcoLi9ycxtzYgJ0/8ymUXgLC41QrJSisfBT8bH8E5lJjwbDEFmnqRzAzd7E5mLK
3d4/GhKP9Qx3ErZzzqXqmaDqNgDqnW5ZYvN1H/KhDIfrSKwz9dRFqSixRLRBZP2as3g2+LYEXztr
4BwTY9ouurmVxxY9eQt+eiRlalpXSHMZTckhpNESWJowFQ/ViQMiktrvUIWHguMtLnS65jRV7W3f
mS+K2qpmPohHYfWPCLJDKzh1Do9cQmInuflFgiw5OsA9N8dY6V0eIDpHvOrNBlW2rSHgrN0qc3tg
K0zHrbVAAa/H/o7/J6upSrqDzlR3H1RJYzlHAG6Es92OX+KsszyKsOBuG14zRMGc4nrmKA+ApZ7T
2U01wK39R1JgXoIbymzTHGz9FvCpV0IX9Z34WrBX/AkuCJmRyBQhStGJ47sH8m+LEBOuzmjpJunY
CzTHwD5FyL1c0v5aJXZ+h8/JfUC1HglhCG3vFZvY3K40R12T2akoAFRvESKxEKpNpdQAUL9dv8r7
vItFkxFiaNAJywDDkF/Bxc/TP0c7Ngs1qfmrry4IjnXV8Q4SN8TOxr/uH+HDDH75iH9t3OlNAdBn
EU+DypNb2zyYd1H3VfzVCOt7ob0h/Mkkf7sKoQeD8CbpugVqnf6oR+HBfsZCdnY/GV6z45O4cZfd
6p8BVeR/b4zrMBuyXxuoejXT54aUJ3bvnhOWLZuVkhDTN/zAw4CAEM2feMvQw4Kayx8cK9NDS1Mh
NtE+FQttp3AthKUrxdQYR4CTgppADlhUILnH6nyJ4nqKiZ3CkzT6/0jPNhA5FEBQmYrSzWIKQrTm
sXa5+3SvsPVsexrssNBMD9cQGt2nloPs1YfCnkIcchC9u/kXJVbT+mTFd751ZXDeOsgh0c9c9kAG
nFjnDxVIiAvUIly0NxRsBjewpG8pfN0qTgQZMaQnWGU8MfaYN1ChaEyfH0VK9557h7zNHyn9Bfdo
bmWhwQlgm7legRYlSjMtmUPw+TyEkIY2fIj56v4yJGJq7SPz5kAKSD25CYpeTNFZ7Ow60wlVjHH8
Xnod4m+6R4vJHLttalxRTTprxfBs8DDYfm2JFzsE35GTQdOH91b7/spGGtBY0DHUCTbdeMdbly95
8zPPw7RoY17d6CDma7LsDFtsRyZL/gW5wutEh2uTU6Fi8qRZtSy+jASvDt+OfucLPnDd04xy1NPC
LwEfo1puXH8SMcO/a2/U8IenopK5+cIX8kN8GvEw4ppFKmytpVa7J7MB2T04E8GT+DwO9AO8oHKG
yef8JLshT4Xq6bkUkY3Y9d1b7qSqvpRdHHaTKgCfz3+91lqPJJJ6Xyk7YLADd+WyynpfbBhdPMWB
8gLBb4nXuQjBOf6YaGxO34gHknl0nVkaHTfikGZJSP8GpislZc4cwfqoS1JbVX7FrmfhGkwqY5cg
Q/7tdGNeY49C7pTSJvLxzhF81cW8iy06++3EigvcgfiaUmeM1tvYd6uHXYMeLjlCJ2obbJYQgNV4
A5g3jSvLCqFkpH9qIOdtlhDnSiB/OUleKfHt8C5lawnaR34OFw878M4YdioulThI0A6uMLJ6zpq4
UIbv/RMNX3R+DUf4BwH5k3YvW97MEL5KigM9ymwrTUWqCBvkJB7wESWX6oHDJcxya+C8qPhVsHKK
ORH0iq3H9I56BXv8Wstp5mmOyeIhqEjSRubwbA9RTbu5P2CfftajhCEBkj9J3q22EPPtA81nnW4O
dPZVptoUo/W7qdVZk+rLT03OGuwOG2eYIulLSEbd5o6KFaOCc5N69k43WFyhqd4TlpKtB56nphVI
g1VfNRWmcvcI1u7AWUPxVfaQ4zI/mW5+Zz4Z12kIzDfQ6joI0jqkgdIWBk3MnNGcVLThAHmJBL/b
ZY2Rl2O0W4IBmPtUJGp4FvkgN0eKck8ek+jteDko/6X7VjortD8mVPnNjxxmqDvXGoKk6cJldtH0
RhxyuUI4Z3IXDR2GKFXJwNUO866BGex+ifmOBPGmJbRT8AydbJGO0NpmYH7Rw5pLGWZJDEa1Emkt
qEW/6oA3B7ywJFMl6mNFUb5mgP5lPoG0a98xWnNzYfH3oufG9aUmMk6o766a6pCQxD+4y4o7rjL+
7FP383vkXj/Kkt9omc5U74DBIa+BA1HpypC+ZaqEVsP4yN/jS77uKKGBhlHTExtHkL0zZtA6FI2M
fQrUEGh3CZJIYDRG2RTdMiVgvIIecP3NjSHBjE/NmeVVNC+5J782D9NtdmkSmSc732G+I4i6zJlO
q3/DbVLbq2s7XJvhWxO90yRw7ZRdqCjGz6GrHrtHWG74j6gYU70HvvL2mP2hmtKoy4h1j0AYot81
VGS59uf1hh1y5Y/sJ45Iq1PCbGbs+WBfYVT3SoieydVx/V91pYZY7M0P/VTcDxG88Y+Abg6ekJ4Q
NWKswudOgbTKXknW+p567e0ZUv2J4ZA+xild9eJM74DYqk7l8fqXErgSWQxfGyn/RUtRRLWcpoT2
t/Tv7RO7YijuFNXznOnP6Ejr3+PSWvNMh1pbE2/QvIbm/KsYmpJHqmfX+NYTThG2VK/oOjVucwJT
PAVg7pl4WeJD6m7X10I7yJGM3Ev/nrIL9TCaLu8ifNxknbpWBTcB7PUnSkYOBfmYJfxMbSJdJVDF
ZqVMbZSb7uYrBnUosvmt1A3AvIUSJTke9P/3tzvEycv3ZH83032/T/9oQmaPW03rY3hHTAeDM1aM
Cq33qwvqKgMcs6TquYWNVf+K83C8f+o27Mb5cNpu+QUrILqVAVsQl+29GJq66Af+4vD/r+J9GVsk
FzSEd+wa2nDeQrKbKret7B7FWWCp4vnoOIleYyBKn77lSI/1Q+33zZkfZwdiVM70dsPCMwal/GK4
NNoLo777DYnSLnu1YiLwbVQsG0Qcixs/8cg92CMMvDNH3Oc+j/VE939mVbhxafNN3d9qSy/z89iH
gcN7OEzMDJ8ehH4SY/0xEYcAb9XqlZJ3EP05LsdYB081jY/0v2ZCRhUrCKuYkN+pCFDjtumujept
or8nK83YXuSlVi3M74OlTFKwWQ1cZWG0Y8Nb7RnhQLnVe/B+paDsr5rdX1RAc82wJUl5bRhHa2/V
9nR5eINTD0DdK66KQgv+9gJYq/exCLiCAqc0ukHLI69cdga0ztbxS/zpGKJyz4YLtE7TXAoEs+WR
aGOkqQXEwGGaB1rzRff2ZrU3mzhgBf7qyr3B1Q1RUEm+FYw8ehDzQNCXdTlu6NPJhv5jT6JvCIxe
036tiSG09nwerpyj5OST4/AmUaWwJ3vR069ymTTjWqTF1MGtFcEzP+oDG/xy19RiK3/eXfi5Io4E
bNz8eYmQGga7eWiLTz3NVVzUtci8LHFIv0Uc5jdOM48ephakZmnvxGK9I5aGBTRyEIO3xf26nK4e
QYOS363DP4LkILk4aO6+xjlThJ9MbSemqEsam7Exxc3XQKjaFNcW+iedTMKNs66y2mNJ/Lhgn1/p
66UxgTfDsIYuvb3X2Q0HIFfORY1rZQqVRFUawdzSXal7puJ1FZLR7aKqTel72K3ECtBPxLpKhpPG
R2Y1g5BultB8+84v1NuTgFh26qM8G21Id/bbtph0ToAVpRqMB5Fdl3wj78XHZAjSDO+3g7WyyXz2
unn5TnjsFTYtEV48xKZcEboIA4BnOfedmYvrO2g9uDx8cGZ76qp9LTZTXRQ7tBzsksq7gJ62H6HY
pp6L7yYsjZZlqBOvvuTX0wQS737hJoG96hWLxNYCRBRLISMysRqhLoOBi3y2GChBkSI9LALzn+NM
TEMJg3txrDEzgTnUK7CuvGsMndWqINlR/A+LOebZPWsAoaNsEGumqfNjvO7QeenStFoV+4KYWgkD
NmFhxPwg6K9d0hCjPrDzPhNKvuB6Bp2x1XM7SnvVI90zNwgqpEolshNAqRJmoiO0dUJFy4Uj9sRN
U2+1QigZhCFl82VRr2x9kmC3lSh+gJaas8UDpFE6a9oxfjVeut1bBmBhwlu3Mohz70oms+JhYRa0
kRgzKeErVgj88ibBcPCCaNyoba9thLSx/rjNIZ0yyz+jSdN8Tb+I4thw+cj8IflB1ZXAX9XiLeHM
s4YnroUPhT1NGvneDiCmxoEX1l+xGrdmEFnwU8WNY+lxYLwNvqn+bgRdOpDSMboRk8pE3IF/u8mF
Sf4s/RLY4dQdV9nR/T5aFWQywdzVKmVK+E5gvYqnc414p4g+JJlzzV005Xai67mYq3WRfAoA8fJu
QxgfrXC730iCPbjbaNfClDMiPcQX22iCkfVR+tG/JJ3bbY13l03YKrZvV/SDVBOFn11jO/Al/4To
YLtaK8WUPkM+UIPYTl+FAJpOTanG46IBHZpFbWsU47IyENXMC+N4o6W2Ova0y89UCv0+n1Ohn+b2
Qy/LpEvCEOaTqB0nTiz2cdBbFob9g/8ryEJoin5PMmqHIGapa5u3sSIY8lsU+7/+gVX4yajZJtMu
vCXtQb5hHvQcKL8T6H/h3bA9g9+LetlIobZUTc4yCJCdyP4hWa/IpOEdBtRgYMG3k5ClGprFb/ty
akiqlNBJ8ZNyCUSaYVuA9tRy7iQxnQHvcEyWCbW8d77S4dBjLCnC0D5UsKPjy0DM5Jxqa0rlolzT
rprjeHv30aAVkzAOSWhXdAud2PcSGHFb/IQiWxttiiQjYoeQTTuLecV+1vIZpHrSi8cIF3JhQ/Xa
JE8wBpkqaRSwayVsoIzz7qjKS7Cq9223aOe7uMtm/rnCZWSaD4ACmh3U5QUAXdYx2Cj7SYHOJUAL
cxygnvVQUXxGF5bdw8r7qcSyN3hkc+TpC5I4zEMuNeVpenO4cyHXkfE1DgtntRg99OeV+7RNicai
ERyEEZyWfljNQ33CRrK+vixeg+WWC9ITQUkfhuwpAlXumI2aKOnS/jm2QO3C74JR25Pi0qHgg6RR
rLp2rOS+DbY4zsLH/6JXaolcjLWEgOnDHlhz1w/TXItngDaHNo8DDVreA7sDrTfr8Dqu5YhXCL6S
nWB+OOLhyjQOc7lpBnaRj2GSXrcpqrBIDSWDtpwfILCwk+J5WYWm7LSPlTK75d4nUgCNpDCg7CdV
WHdJ7JVLEpNruXAMSIyW8W28INXKrDDin3PksZp/JjyxDvRMEt444/MyO6YUvKh6rYnVShW7/ws/
BOUbBjj/SVXY82YDpcz1d+NpabGPdd2YNeq1tQbhfneLGymEd18RMeAU1TkyxshfQgpae9xSD45y
cjQdXjl1Zun7inUzKtE1SIijU3eEg+6/wiJxN7iRt9wk6YqthBnRK0MV0gAGaxwVj8272Y61kQrY
5I3vMsXNMdxq9etQH5soDAtergI1pyvpPFgu9W6RWXUYr2ooGO4ceP8fGrTx43ktjTOrmHuj2JPe
7jv4y2P9X3aoKecjjaCMs14wGvBpZ1ns2gR3Jfc/DtuUTlOeyGN28aHue/6JIiIGGL0gv3HnaI04
/j8J3XSrEJSWlvutEGnnkQDBJ31qsnkF4xraLOUHov7d4gO7bYuJE1lrolalpNZ23anui7khXnIa
FFoYejFI/0mkv5inmJvEIEulRBPhtah/5fCXlNiN0GRqHGhvb6r2JVNxLFF354AGvZNaGRCbHtcQ
J3hvb6ubsWjqfsRsn9p//eDH8Z/ZOXtsF0INwJBLpVMxOrccH4MuzH8SlW0njNx3zIThlnjPlEFz
UlAJ5+ChvruaiZlKZAEz67EdH+WCoOVunjoxJk2BkPUQjWc6n8RF9KRbBO8eSWsaNRL728/fixU5
+s+hVnOIycPVD4wfRQa0/4qSLmSkHmEfQJ/7JxqxN+4AWQPQ0YhAO/wSbD08qV6sy2fz2soCqhVP
PSjL2rctZR1806F0QXJGOfNLyCZMIhrvRYVczT4Jhsr6lKcDYAS8NTnJLW8tLB2S21fCb29Ri9M+
H9YbjIONmrJZgmmR46C1hLvrkVTZIKGPElcu8y6Qbr/jJkso6eW+t8qVPrEUxrAXDYqHhJkYzFpT
W1afNB7Z/8NOM3OMbRh5/lY6Ou9RPsthQvMIYm5c2IuAvJLcNw2CWqedguLnIwJaDlVDbxAugJZC
DUvS6pW+8Apq5vsIMKd7bbck7U5Ep/mjgsrXmC6vWIVdPHA5p+oAYINz6hhr5GYqM8CXDSoNC6zy
7nZFuMEhR93Gge0u6Nl8syeSqa+EPrF9+WSw0NsOcvGuP3FVLoQ8fcX3cNnRvwo/EjLo128UbUBJ
O2xqd7XPWFH4cZSnS1WeNmVGWWa8SGOAbDN8pud6YqvY79D5T52L/caWafK4YGMH18G0WwoKmYE7
t5uyIdx29O1OoxXZiRNYW3EOkfhhbQLaMlQ1t0Js5PsIpzGOd/SEQbPGln9qKFRnwDqDJ9HykWPC
q5zA1FpLQM0H/fsCpL5RJFCgUw1jXJ07u9aXJAzEDn/82B3krlh8K0oNDE/b0xn8qgQ5whn+M3QA
TW/4cUNoyw1o5sHC9zIrVS9RPQ8oc5TyQnnLtaM3veMqBhEpK/gaupntiQa4blWkFexpvxbeAuYH
5ikgD8QSNe9eBSG8QS4PsHSwGJYcV2ZfgFUu4WiEMvMfhbVR7dpxBrzSm7GYfn3zOTtCOulLRq/O
GLKWclC9blUQ599ElzTzEFgJJY8uf2TiCLn4fIGflz/h1oC4Th+upn0nKKwDaFF/9OaTEmwSP57T
xWz818gjBbyvs1qRhb7bAi8/FiyaUMBp8HKoQcdL97vO+OU/VJVOt6JJWlTLVNLwqpbqe1Te4rPY
xZKIEmjWbOKw3Jmm9/X3EK0phebXJk5vHJCvao+9Sko67IitDgcU9ng+79pgCumdotwJkB2whhQ9
3Eixu9K0XZGbIHA3wTCIUvgeBWhKu9ysGtR1Xij8Bo4B9xa0kbyrf1NKptQKd3D7Tr557i/GYTh7
+qrwuwHV+nXSbgTmrsLCQXfo25zY/swtj+d7g5SzoMPgiWRhWb05pmlhmTIEBisQox8HHhHdUIk3
HzxWrXNaTj+TIoVB6/E8odrIz+Mul3yTz3duZnSjbQbQt6alKPLTOgrThNJXpQ5Iphm+ea6Uwnmw
oEwwzMblGhbq7C3RFox/JeCIOMJw48aCth9cX6ckk9hB+gZ9LOm5nBqG0VmjQX8cPrpDMm5TX+Qf
zpBNYisbpkdn1E1ibj3/HLnwcdcIH+z3ju50iZNMJcphzwR1yD+BIWKV+WNFEC/FPGeFZ2gpRmD/
auD2s9VQqNm0V6KSJMZ/lSgIYG6HU2E6Zky0EFGqnCM+irsXsifh1XZhrOAicLW5cLOOomfKv/CZ
RUicMv4km3Lo2M0cNx9Jet2uJuKw5eIXbgllB8/gyrp6WcEDUoSuXDUbZ4n4Dmj/QxlBXKyhIVZu
DECh3i1ck3KKJbA/fvutOWVsUeN5WxApYQKd5dPxHnc1uUycITUQPXnQvcO1HsjrJPm7+LPhWPdu
7EdtlqWVai5ANhY3OsT8H6L/oTr2x3DJM5rJz5QSIn75ZJ+pFcmyRtaCQUp2NjLyAFhHgKVazFya
xe3Yk7IWbuIEr2o+fISffkXGZFmnnapmthNkMQ0GLkYBoWLn+xDLAQ+1trFVX99ufl8hQ3ziOKH7
CDXsECuuNHIoisVAQ2MMDaLWseoh7YjUbudMR+HpwMQPT8mvxKKU1sbT1ekx71Mha05rrdl7+5tT
7D8mEpOX9w6NQjdDPq+qecgHoJzjxiFWueF3KWYSeS4QiucprtY2kML42bRe7354+s5xNxerXjG8
yC7vzWA+RtwKIZ66ntaovKpPl/fVX/sbGFg5BYLPm4uRVre0pWOnyyUpp101TUHIe198NP3KEW8A
wU4gF0NuGGTDlsgLbVqCE2uHrGvodNM3yNoyIjKg4PJOjeiC+B7U63EeHz/OC9Fm6UqJjuSoLoog
kbulgpfIEMw6vxVcFsrWVA++137kFh8BPYN6EIRl7YiZ9YSaw5FVPT5VOnfqLh08UjaSGecrwNxq
0vBoW3KxqbVXzfQJxvETsQvMEtFiEZ2wuQkovr/wcDys0/FTrz4SQwg3NAod3ecW55cWjy3fAaai
01fsBLrbpRbmQdG0A/lNiRQchnSWS5fgJ9LREMVsy5PE1+DJZ+MEq2CyGNe4FT/2zZMxyXWmBiKj
Kmlaj/ka/+HXSpkD3ESLGXawSng0SiVRpk8XHa4HNJVf25GVxe4W75y/7pdkWo1uh31bMXG6/McW
p4ORx9G4mRC+uSfQIkG3SBC5rw7oP/kqMdzbCit95YtgRcqrKhMfCPPPNMQvHwrEvSsCmTrm5vwg
/oIn7Qfcv4vTjeW/Njg5YEw72h/rEab1XUf1N0no/vRCPZJlWIqobtfD3m9Sece/LnWsgUuEkulS
TJeHbChusDKQzSSpUbTVogiQQDsE2nqk/yo1tl43BRD2NTBVjpCsSuXzwSS/FOTMUDWgJseMGtKt
0LMwQDg1r4WvLFiMMPRLoraHp5gmz3utRV0g2J4HpakpuVR+O/j7Cz2mRGPwAAWb0Y4myHOPi4zN
mrwWcgQJu0YqWI4PzamKVT2O9kqP6EEGt+4Opmv1snTIaV+n+NdFvBJ4HbLNtES3enMuYc8kGUMI
vNOSUQJBh6xRc4ac3R4cQJZHIMLdwkB0roKrIgrQa0Fi6s6FBOz2PqvvpNp8ThdFYlgpK9KoAfIF
CSKiMu287LW73z5SAFfvKIbu6La3rnfHQYLQ+ozRnv+DH38eCpYZfqqtKQ7KnBBCnX52dZXmB5MN
MLmvQoqSxfGgwzCds+rsHdjX81jPjwA64BWpHbaAIit7UDTZwcxwUMQ9wd9TqKS4gOPzb9zMZYZ4
HLPRis1+SUTm6T5yjCV2v+63zmOhLmvRvpJ5HuQiRBcoiVIsPql+9FSzPvTU64LXLjfxtzx1xuWD
syiHgX1VeosTJ236UlcuIC9oPK6JFvLrPhPAnOUmFANT6NpMRXdrvy7o22do/NrJgC/qwQ65FkrL
9x896FpWjEqk/VgK3LihKUoABioLco0jyIHV2/sj+gvapwOjG7kI9oOC8KFL4/2np8Scr95eiCTT
zr1HQSeKp6UDOKc7JBXCLnrX4zDHYyfrfflaK6ksdi5zhVN8Ivb5kbP63njPqO3FFKM48IQkvKwW
WaCWHvyKX3I/0xyEGrs9PMilU5ryEeaDAefxQu9XjH20HKP+zCt0qBaeR9gDEZInZol/m3gnaZ7k
iTAfJMY4+J74k23G4FYH+QaFFsVCDuuhl4RYGm00+9U3Hp+oAPjri2el4qE8NJqpsu92RBUZv16K
xc0rXEBaF6/Aeh14/jNLZSGzPCInjWWr4MMFV3rFRLcUI30Rru+qOnw6Slj00d7bz3cWi+soidMW
wqcX3cVIHwJHpGrkQ9mscp80yYLb/H8LeyhWRBUhpH2Dnqh3BlKcw2aNepEjHunfYF3RX38C15Hh
05I071xEbHVnM14TyOJKLDzyEUWAEztwSbCvJ7MvvPqsv22RWISjvDKJdDL/kwwLf28agQW1NO3G
mngVtF2yduHN+X8HbirDCqOgpr98KyDlcEGpHCuL1AirPh/are1Eg6wqMPD7203/azBZ2NYm3B66
u9ARsZSiRVuQd2oJA0xnC5I5JhqJoQ2LmpFIiRetIGqO/yZCVsE4+AmxA6rH7zgoenUQGNU5p+lw
cCVa/WBqpB102831ss/CD3LHi865r9r2LfpHsCDvXpGN2y2To5PCxhQSayb2R4M8EHycte5R/RcG
s6t14YNWhfdk4vlDviX4/GEXswoQMGwlx7tCAfU++xdBiMwlM9lxrJKWapPYLkPungw/46pf2Yb4
Bs8xuRsleS59e4Nky3ud7muA6iualJVowBfOrhyN43Ld0tThYYIG4uCerCDKmXvsGKkdbx6+0q8l
AQXwh82xwtMKW8iJLVztKyKZcZzPmFSA3FONaWm/boCrQL2yxzwIcfu6D5djLG+SKarqdsXhj5bN
2luNVBHjG6RQKfMizxaz9ZfRsBhYfr3xsbGroXmAh0aE1GvL6mA/tTpNSUL265YStyjo7T7riXl/
/JpnVeUqhEKLT23BvPhh2r83PE+PohlfFRUWQU7e5BTN8S3PIRMXxpSQVaC06vZhluKeUSkZUC8o
EtRg3nO9yBooTyPiW8yEWWMUBHolO8mXix/wLCU8CnphHBrww77em69gWks8oyaP3LPu0axK8yCK
j+5+kpD7pwIT8+tu+C3IczTiC4VmLLIUQCB9D5Rpo+O+xvSF/k9oGoHrR5Rc2+ooXAeoB/FTRxpT
etgHPv0Wh38S97EuNk3j6hTnkKCd/2L3HpDe5CfDS3j8CD5BEHqZLMUICSCyUeBmLjgMpEqVg5FL
wiY/abN8O0QZ6482ieQM+XoWISsVNyxkn9LYP9f3pp6rrVWc+xW18/DNqGf/rdJsFDDlXqssLAuJ
bE9eUxeLFFDL3G+INgZqMUajJjCU59KLCGGb0QiQsx/IOTqXi3/x8Rm7n67vROhSmuljOfI+foLH
95QPwZCHVEFWzvuLF8CQzJbCFFPTK9i/Ahg1R0mEgKJW6RBvaXO76MT6oRL72ROYWEvVwYO7oC+0
TkHM9uJEV5dNBk9G+Z9johF3k6szFJmSBapNJa1gmAltvx1fv6cnqf7Ob52kQ6zX9FW65akeI3rQ
lkdm0T5N+6eMftILHxB2PfDLAauwYCUYTJ24BtvSZqnfh8TQFNZLiS+Ni0Tl4EHb6QnuOZVqcDDU
spjogQYAmDuLXTHwUS0BOW41jkthDxJeC4GpRuK/OHJKQiWH2SZmHH7s1vuU8drEnVpPxHMS9D6V
OU30e6lrrY7KmfpA4z5YEC2lrFmHo/57HT9z4UIqeGqRi6QgnV+5M9jwITjJ/heUUStSPzzxaJAQ
vUBPM/psY1AJCwM3inrbKvlLqP/fdqrf59MmxDmR8CCmSC4HE2b/nrgyvi4e/cscwCHMUI7xd63k
57b0/HS0nQ+9HxEqh0lHmDc7f6LKgFjoOlDQFidDz+KpnMV3XpwcZvpcXo4D9WPIZrHu/SD210F+
EeZAOkB1EV7xMidQDJ3Y+R1i2s49nDnTXthO/Wevu7EiMtiatDoOhj5r+vZYlJlqM9pVvs+n8Eat
HRgL/dyzfjlY4xojDmaVo9dydX0SvcOoKkwGasEP6nHknAe7sYCPe0yTE9YqB8WRtE0Knd3Dj/pq
mJqkJCkvuCSZ9XHQvtHd4oX0bDTbUNQ46DgCdja1T0K4hievjE5DnU0OTEdXvDGr5EELkZU6HTh3
+PxQl2Y0Rnysw3XhIq7jBSGVaiYZK0gT0yIkGlH9PwURtwabTxQwycCLMT1WivV5nF8wW1rpAlbQ
x/l5L+dRD3Ah8d2fHiEhVUmiuDh6PA12AlnVf8g8gHZupttoz4wA709qZNK9AKEEuyCfufIvQYyt
Pyk5xYLeNDDLFgZ1YZXXCrz1Esc9AOiS1wdfvABKNxiwSUzKaPFsZwbsLErBjzNue444y0J0zkq0
p6CpHNw4slrbjF08zjluhAzSrv/I2XuEtnyLNeWXeZ8pV3ZncxKgNurtaY318A+ifREAdY4k2bYX
ldHkm4WnASJkg0klJiqRAl+2m5butvLG7WIGLnFBQ8WD01P/gZTV0Pb6BMNH44UNt01Xkj6gMXnh
/ETiVo485sZ83ovBT9BcLVwzHfC9dgD0JpwUxnjcjbc+dD6uck/0Bpj68V+QF9k69nmJhB1+nQCM
/EsLhLyeNbu8h92PQqeR8vF/xyz4Px+l3Vp/dVglJe8FtneIZxZgp6U15o1t9K0Y7AHLfRJLhSej
QqQPcvycpfTG5NhnCd0/Iypn67Ms/7HwTroqbw/2mSZtiQxBxnGj9ps34gHaKpOQkynvtFmUvkx8
3mY+rEy4bVDXlc08jdFq8LHgH/XcjbX2npMtoCYfTexWSm6GjLidSb5tEa3Kr7mmZXnvjaZUu1xh
FUhlJjP0rWYnyHZts4TZxnY3FLqjgiOIWUgIj/I0LEgVApujD0hzt/E505Y+Tj6ASCDpPX+aB5y4
c2Q++H72haC30vH9yJpoQ+emIfuZfnfzZHRiqBX+zmlWu0ZSRttmuL1gsoI5Yx3/JwIT1QENjvZy
9CVKA9hHX17fW8dtnS7Y+htH5iW+lscgX3IRjQoi8fYTntPVAwKFzlE6ZdM+dlbTjqxi11M2lNPL
sw2agIETeKqJCgvbThvWrMHkkk3G3WgKOxVigLl5FiAEpzaH3L1U/jUloJBjDdLoNOO7ckJ9oTQY
q4eI+lTamBXUzb0GEL4ZXj23TK5/DtGw5KCx8GNHLKqb5/Gl1+gPIOO/M2Nh9eOV5rblF0QlbyOV
olgv56Jdu696maPEzpY4RtWA8uJ8FSZ+XhUH/F8Qj/Pu+57rR3S8mDtr5qrcfMu+sSBOzFK1Fs9Q
nurg331XBiIrcAWGqUXF7OBlpfJGcevc84erUd1G4mr/A1ZhnedbC79UssFlXaiCO8Dmzs0b038Z
AoiPbd3FRSUq2ywhSmS4BE+zbMFsQZLuaRSB2tTlsKY7Tti5f245GXmEb+/LbQCD91SFSOhpXQ5B
HwCLeCCbFHe+q6QUzsKqr7lUNZJa9+5pyHQ0yuinNH8lvi7LIh1R83La7upnlwo8ma//++Nwp9aw
/kkcbla/VjIZHrL03CE4cIG8jJMLxBtlrjzZAaGI2tZIT7f4A1kFTMrfNw5oq+FpeZqCjj8IK1FV
/gUhpP5UPBFGEE/0slaAugX1tzq2xbmkrfaayxZbas50fNGafiitcSKdZL400SXlV+23DSNRAmLz
5hI1Ce6QQCZQXeEu0b4J+2N4BE0lEQiw1PLCQddVWUgx3dy7zqo/dbzA+zW92e03hnmeP4rSZ9SF
ybYgcy0v72vmcBO3nWYTugjo4q7LV1+wx8kiHwtxVyvMfEXqTe59RLCylLp1YsuqhopEoPalAMch
iWXydhcF9WSRaYGS/A9tk2bPz9Z/ZJ9+s9p2BQZA6G4Ae4kNoWZ4eL9tM5rDiqAWz21FPEcplJrq
XZxlrzsKDZZIGrcPj8eaRBP3a8yZyaJX456JwDrHBEvCFnuAL30cYAzdC/l9cZff1OFUENggPCdY
0E7i4rPnebKoC9Z5L1PSqytsX2CnLGuaX6+Zz0VvGbq6qM5qe4IL+wCNm2nrJ0YlilUxtyLSFS/Y
7Ob+3ucs8r3ReqLnVIhSbTC1opm/K3RVmw5q+pLwdw7HJjafW580JKfvVKdwt1Bqar7W+gC3FKf9
8HCkvyUlfmE8gFyoz8QddxmnPRcdhFYDzBdja5qyIul1hJxVFbM+NdOhdksutGS4XwNHi4CHn/S3
IwsXTf+niIUw909+YslxoQhAiJR8Cjmvh0RA+lIsJXxEYpGwS4mGh/8cpTJ1VnRvkkjvwyoTksTA
z4h0MEYYcfDVsFOiMVs1jWjbfVDPRbpxR0Kn2/Z70IuvNt5lDO03dpvGBFs3gg1IC0TSy8eVM/99
PyXu62/tE5ZKfbm+YujvNKUynYbk6UkzmeXeL0T++4+qtafcQyDM6qAYDy7Dxw1Vrz9OoaDDVlxI
C7sY4qzt0HPmfY36Ha3Ui1/xoT3p+AhkvfbqRa9CztU/4+hJKr4/V9TSePeEJXo5+stwM2c0fjIp
nia/6vHz/sHoeT4say5zT34zfG0knHi4MAeNzKmKt/KaDp1nFhzpFUtA010qJMx+ydaI4HUZIo3Y
2UzQ14HZJEYOtErqzryEIKd5DBmLJrlrsYPL+O6fjJNe6bBoH7iNV5yjVQnLbHHR7648HCPI/s98
n6r2pMu0jSCTAVN+aVZMWJLVYb981fwSIOF4vYhoG9UMiDgSk8kq0Lg+sWyQgd8QuWTzQF2XdB17
1H44nL5Ayrc+Z1Yvb9NSPWhlpRJqbPMHNWKNQAOXXWJLjCEQ2aohoJRyWuSLPYK+9PwU7LMSIHK0
O23c772F1DosJw6HTtaCtIiFQelbvWaidFdZfeRTghVLQ1Z51A/6Oc6XrHgtfsjcBlDFOvOLJz5q
nMGsi2XuOTi6Yo5jdhWFrINfpHWzd42/Z2JJ1x4JLvBR9NThZM7DbUfCmSLbp0UuCJtL9u76qdEV
sYfmL8Or3mxLsg1EwffMz/0KI1JZM/Hci3suqUwc4etpCba2Rl+Fj1qzxZN++Fr1xcUcZ9JILuJI
RmWvhkHzEC52bLmjoBCKW+QOhBuUiV19qTMobtLY7fVQiw0qHVzpdaiclV+wVAXHKFURF6aFkZQj
+lRf//M6uZzeMPC9CEeQVB2F7gHakEdJGE2JYWj5AVKmNilF2leCBVz9YsyoE1l4WI8+5+tjNV2V
xJtJU61fAE38WnY+v3cN0sZ+N3eIzC7cUOrejAHOVACWWMOk2vdJ1ssVwYCZNHCB1LIKFRoRHrkX
u43AmZeNzkeLgqRwd6cO7UsTilKH5MWtMAAeB37zqEeKt+pqSpHqT1ndG5sIsvygXLNt56cUgLIB
UerlwE3g4jSDEXIfr+Rtl1ZaoSTkEuEbZqkq2aRaZ6mkBVfGdnhvDP1+K6ivw4VXk3242LNYUEx/
eOqR8QmwXYPvSchvVo/HEfJ0CIiku/p1QOoHtIvYOD0tu+ClkO24WENFioZnHLZdSLU5VRzSOMzi
v47B2KROJLA4YiNT9vnmBhiIoKgZBp7tYpU+2EuSyzS+HzSBhmB2QI0tg5wnw0DjZ7TbqmVtrLGd
hjy9BIs8QXW40OwUYIP+BhQvCR/dbSujEXjynZCffJZbaOOLG+0akGrl0qyx4nYufLP1mK0hChtL
3rWq/i/Q9+owk21DhkFnDB4mcGsCwdv4SaCAMWGQtyM4ep5Xyzr+8PGt4L4dYGKPHsBK/zTjjn4r
DzlzPnfZt0fI6H/9jp7k7XECrfKz2qBglKOa7T1seblnrYKlSxOXdy7FfylNRTzAQYK/P7pGF7Jx
fyT0ffLfNQUbvF4HBm7l1aIBPvf8xtcWOMnzs53EKFTbwXSlQuYKb/74ECqVbqEQpwyngBJhKR/O
gdd7bdIMTK9zsvWhBw7o6tJHZzsiOX0LXsohNywDEVXIOjWMtJ0qu1MTozGIQbHJ9HlMAYg/m2d1
yBjBRwfxBGnAjcwUzp9IUf058+8Y89a0iQXu0xyOgTJT1BBsAXhUGOPk48HZdlt7uKfxZx9CV+BB
R/amc8vZpzJO+qaVsmkwQ+Hy3Di7pJPhXb1FvQ9j3rY5weikyOXGoQ9clFhj6GUZjLYoFIkPh6gA
/UOahrM0yCXaiM4Knl8rlkJ16rD3wku9dS4Dxqd71DxNHutcdTIcrfhhC6iNJIfuDVL/0PjX/8Kr
8nh4lG0z3pNXGEIvrrW3rd1267ZY+oZIZ/w5nKnn73YgPMp7yGwFS7vzmc2XCLFNkPYi8wqrejTG
+y1NTZKmXqp4RifxP9z1G6QbcCzoaSVCBxFNgjm7TJLdy/lrRtT7UWP1A7T69lVIxu4BPaDKn+TS
oaGWmpGRLh6O/Gd9ydWiXL9zeRaV7NQzDjYkyXaw1d2bxZpoCyz3I6V117tZP7KH5JUzD1ly9cwH
1R7IMNaEmJ12NZS+CeVw9NOXDSiLH0BiO798ziEtatLpNu6TfeErX+/q1QPqoLlAZWKLlHrWvDB+
z77PTlDAn6C4JAdAHhZdd2qVmLRWDH9Fcv+rvkEphOP7Qqc27qqflzQRwk3rlrO9+z+6apa/n9yH
KHKT/53XucFytpsydoh+xuB6D+74FY3IlmShZ+38tkn/LP4qXQSK5SOVfZf0O13oEJXP9Ec8qS1C
8t0sP0Os4PzJCtCjHxj3osiMkGm40n88+M8lYe0ecY8HURYcJichp9TBr9JWmWS5lQvNb2Tr1kcX
O588uk8kOwgxb9LP3dohiwgJW4zg95BsikvuOp8CQ7R/oV2dXF/x7qqNsKH9DUxgfBk7s+6bp7FG
Qda33J5gHZNNG+cnosYHsksWT5jnD3I/WptL0s8btGMcueP1wQ73x/Egm767MF32Jt+bZ43K9dTc
G0svRWeEmQygtUZl+t6J2Xit7a28Xe+3ZBU3P4srEzGjY8NBsGi6uTl/ImjPdRQ/on+C1Tiv1WGg
Y9Jli7ZJKOQ+A0aGmZf7NQhLa1dXfWrgd1xMWVWAQQlZ+SvX2XBRhh2wC/R2RH7Sy79CZBiNNdG9
BZJ/77QMqMU3SsOj2G4i4exJr2uIA+xcmf+7QxQajDuLs/Ctv7/CVkHMf/Fmou3V+12aJtDT2yot
rzVBBKY4UeN32saTORCoHiRKdBNO9aT2qJBvL33bdW5aYqhokolHdfoHFEnPPU4Y1r1LmjdhlWcl
xFamAQaWID+wCGqXcSA9N6wdkA77iThBpYuzQ+faqK5F2RMTS2ATYCp4q6/1z3xKl7LlIxlqZpQ0
RedhOK6SN367bVE5xSomPWPgjfrAj68aMuFeaTt4dM/vI4cTES4jpEth5gGNYERDXI59HSY5W7TA
foOeJnrgQeN9869g14Fgkt7okxYbUUEvAyYjO2naXMqXBY3IoZuHk4JJqPzPRQkPiOgzif+GCWJu
naopkRseCGY8KLDDDXcNbQjGvtDj6tBGhLEfgjJ7xzsX8nrruTOgQHO6WL4m3iHqJU+E5pDLyOsb
uWGdYKlWDlfjblq0b/9yn48bwthiG76hrKfQO9PbKUMSHgyKF6n4urT+x6ka8LvUimVzDdbK/Rxz
MxT/GlVKqz1yd1TiYNmKtsUGyXai/kzCevhBN7bhPhAX6LPryfd02JrbeoP7uOsWKag7m68sdSLX
q/VvRCnMQstvVIU3vn+cGhih1vqA1s3ryBRTyTb2NzwzT5a8aRN+3W6reABKXKaOFk5VXHxEG0rw
O9OBkw+6bAi4X5sjezuE3xceETZUn6q2fDBkEMKV7sbqCoy18urX4ZpqCAqi1hQaMR/PBN0p+TvY
Zm6cO2wm9WukI7o9AMgAlzbo6891u0Beb7r2fpddeaJFTVoYRjSH7qk0wH69Lc19EYKNU+1LEyEo
ygnsIJNUIki5HlPiUPb+tVW7ItXtH8W34aRHIi4oyiO0NlTj2LjhiPirLeiPvJu8Xl5vwtvufFnY
Cl8WMatbKHiTQ4mbMwt67wVUkPY9Q8CdJHCwBak6YcAOFfsX2IGORHs6njTq85g3XMbpdBBJH1Ih
ikbVGGAcoFBDYOusfzi6fmCltPOUmZt4F9aM03mgnq1xp0FRcEQT8Kmms+DXUXTxBgn5JyCiucqi
QQ24wZ+RMTFfJysOIRlhmfvlzod35eC6beGDuqB4gJjOA1tyfgwEAh/qlCEQhaH0GnyGSknF4JTp
n6ZhayIRdPpkfRUKFxyaSvdpMDJ2vGcE4cBCTQtOBG+sO2w6IXzoh0oaEz8ONTUs/QI9rZHC0so/
mrKguvbqTmyauaR/3FHBGKmTgGd5fXd8fNbn7bQFbWvO5Lko+pTjzhaXieRieIgjJy3eE13+s9UJ
L9llvlwBVdN8EAyHoKIS8+70lSAViF7lZJVawCigRKRzGGhjIqrDGfGqSMKgu6VRjMuo/ihQxXnh
WOr8tVRUysan4PmISfk1rydFAabI9qMdkJ3dmqtWkDzIsF+MW3ys7pP9Y6y68VEC+KRJNu7BlnkX
2VzkJKVsLeUA4doedSfut5lOQJrKNO/Yu+JajFTQeT2VNlrqHr8MWP/nFgpIi9YzuzCBhKdx9JVq
OFTqus1PqXotgrznpPJmZ4Dt3bs8tBd7rb0auArBZhmkLshUuy4c+ULrAtpWJo/moY1H9n6ftMrE
20f5j5FhxYwY1kqkyl2kzSIRIJ0bCLqJh990mL6Mtkl8Qyn8xlrf2aGVF7Dbt5Dj6ydolJkb2izW
PWk0E1TYMo2kY8GPbESLpw1F+TGKkXUEbw6IBZI2Od20BFt231kB6Y8Ew7cWePJMhteeR9nGvoCA
77inhl7WIk2n2GFgeHSCkZ1uprVENdCQP5isc9tUceIGWWXDQRiGcZJHSDBcQaRnoATzLy2eHLOi
8cxijWWzNxHYpa1TFnOKZ4A+5hNWDcapiFy3geeDCaig9/IBe7Ew0Z0R4PEIIWeaXQzYksapnhk7
9miGnDBTVIL4GnXNvGdGLEKX+qTX8aETUu/58HqJuee5kKFUH/vKpXxHxVngCE46wpnpDykp0x4m
/NL3kzQJLK4shr+erepwuuQtx4q95bGdyXdx6BOUqgR0Hf8gFf5M7xNtr01TVU7fr4ULJ9fbb3kI
etaMy57Pcz/0Xc+mN/HPC3OB3mxoSbq4m+n2jvDUbaYP2R+hrWD/qPuAXxd+SU/izlUJw0Zypm6L
kCv9ZizMaK8J/WavReiuNoNuUofGlRXwQeGfBxPPpHWMOzj4K3L3Mr4RoPUKDSrl96+2OnBPBKm2
IPYSGlJqip7pWPJpjr49n2F6Z2wAidAz761SDF2F72J0Cqd2bLrGNkk4YLnv5nxbgBQfyCPBclA0
Uq9XBLY6Ry6OGaez9yffPhhPIUBiT8xRTED0IALpw7KByOqTHCg4WUfAibisXlRQjpoXL7yiXAoR
oen1RvL35/9HkZIa6UEGEXWMo89qX2Fc6awgCalMLL+6b+Ng5LD4qyNl+rHRtTWmlHwqpNvn7KAq
Er0Xu0zxDEb03Ee/od1QPEFR55QBLfNzWKPChWVjRJg4owI8IXJ2bkOg/3/+2I39MJ7klNkJ1kvE
rAfy1cTERUMFYAufuy6cY4vsrbYuJIqFtWq2DW4ZR49BI7QQ0yOMcz7mHaFw48W7x2F64kinBGIj
Q76PeeSajVaRqBtfrNNnLiPoS+hzu2bcCpaqZKM2uX+uA20LGZrgWcxwbL07jvepcIxCKULlRFop
1i4Pfwq6o3o75lykpVt5ZAi7B9EGdaKImjhCpEnGo0LDexKo4KlHtsFde+LyUpZ+QoTq0nVkqcj/
Bzni89YU6XUOwTGNMufbaRr+DKgw6E31sM1xmevtvuahFC+1upEgHP8y3K+/AIaSF3rHtb0FYRbW
RWIvddfdpPBLRn4YdsEJGoq+QwAvQKbdPX/GcsOevefg3+wMUf6aygaEutFLl8yQ13dS+6dFi7ou
c+5XYw71OC9KM/7RFo5NAgaLHK8a7rPJRic+9rbqgOulMo4nxpvsO/SePc7Hi2gWYMkgXaxQwPAr
Rg8bugq6G4kLgPfTxP+o+ILOHvWf/Jevh0OfFB8EX5JhnhFb4Zahgml+BRdH7bo5ubC45eTe3Dc/
YnqQd+lm8aedUl/1PNbyKuZ0gp+6Y1egrqfz7U0cuHh+5K5sZIn36ivH4F6EaH0Dnpb5jP2G0ABX
XM9aXTn/OEKWPnCwkETP0qWTw3rf6vl1LlQorfQnd8V+RYVklO8pJagHvLg960BU/wK5k8Dcny/s
GnVsi8YzwEV6E0J4K3UIqxv9jjr0jUDIZR3/mnyo7TszVNfazQmZT+Pv7ovyGwdXgg0BL/tIiTLg
ztroihqiMDF/z/Xx/oHFIJsks1hG+26ApfDbWWT96OdQKPOB0aepOgRFNYWNRtfEIyf1YxFAjDMz
56SesxR5KMnnMFNBEjSR4NZ1q2iggTZ+Aa4JK6+0R2AsBhLl4QbltzYSMFh/Mp/mKfoSNg2sKib7
JdfiOCwNjv5RKJGSqVrugwO4nvrev+3yF2Uj4rLuze4r2tWxSwvSjKIvu//0UI+cZLO4UVH5LQkb
RrJDuAgalTrPRXTqjuxoI+tvGmVpHeNE6Kqru3CFt9FQe0Db9xKncF+5W5a7eXEAFWD00PcGZ2KO
wzRuDWwBw9am1ckVT8UTTI5yGOVYKcv2a/G8yPsOkelcrT0gfbREE1J4z5Kd7SKLAskoYtXrgmhi
PCkU9LPI3WS0AglZyT88Nmww8qYSzCeRfoQfZcjVv8/RTphJMQUAJVvPs345Jm7JkVC+GSLtl27m
UTk6Tnclb6OngGV9d7Uqy3GytnvSeqLG1ZWdyD0LhQxFWOF9jrYfJaQPPfC6HkNXbckdP3zLIx7v
B7VVaPoGVL553hS7TgfSM56CwUTfSmW41GBRQBiBqSW97gSpOOA2HBQHI2oscMlz/+R7iV7myCRH
D9GnqB5n6KTzYuXluvzluQaI3lF+p1JddrT+4xEZ1AoY9wMvdcs7j/DfFlBrs9xp+zlmVp1d/0N8
j7ccQon5ljBOD9cU/X39w8Ob2/S/ohskKe8G+uzOMvuEkQkxvLz/RSFJnFMntGb0ivi+PbuwUezm
2po9LGIRGrUdA01jNYN7+LSrudxBRDTSw+nuka1NdgsCsnPpSpMQZuoMn4CXN8OB4kS+068ZKQ4V
sIqs4NMVZGLjMZqfFvp4IOtO6fMmHQ0k/6s5krptZ21Azbd8XbaaiNuaXO9KIiDHOYy57Qu96zAc
6qiQJF5GYoMhU/rgRIv9uV0d6jW1MSoOOnI9B3wEs3+KHxsAfbzqFsA6CvaX14MeyxyohfAEY+oD
7b12k98hfpDVpYxg0t0oqrAeRdXDf2EdwqRcBVIuB+iz87c7Rdgj3sNeOva4vYEMxXqZ5ty1YiRS
ww/S07y6VA45Uehb3Yu8juU7FURr92aT7J6vYQM6RcuWQnuX9xf1TxfJHJYBt5nQs3YvkV8uilei
9kfmVP1fB1C3Ruld0xWH+iIJXlkKHylgLXtaxZuOUqLwpz4VlNHuQEKOiSJJKg9eX+WJEXBFxDDj
CnpgcTn4th7yptL3pERNNhMA4cduCvDmWOsRoUXWmYrZVe7nMEbSjxpD20YDXYsH6/U1jE2TMx5m
1JEW7uV6ypLpT8Mst3y93sWJhlvD9Oc6BuC8qghsq4TGkNU2pImRjYTihW7GUg16yb1jVF2l/Sq+
XETlkCkV0/Llv6XlO1l+OLrznZmlSBAnx9bDhQvRkZ3twmM+wMLbqgplZ4hT6kbHafH5DopfVY5x
S89z8JPgaSudNJmRgJmMaA4MPrjzZSiLkOfMCHaNqC2MrCV+ZcoDjjAc4kt+d2Ogexkh9s6p+UUe
goliSmrqpSZWG8fJF5Ji4cVLDR/lldfIcHzmt1uInHF4v307/o6BrCI1qJuNJwYLaohWkUrRvn9G
0/9j6aXq4pkmnePeQNL3fRaPMNtIbEgiKAEXzJFnEVX3k9vMFvAPfNXmC0XnmNEz1Bx6+bm6cqGk
1n6e6GI5UFWeAOwIQCcG/KwMl835xc+1yLk+OgVzkBHWXLudYt3zaUqVvG3UW5fBoXiBhDnt4WM+
SFB1+kjW2khkljZJA5PH/SvZgtRYDTbj0JCfBAlZPhVbtTX2MsU09FVZZezgMl1LzFfUF6ls6d2c
ucscCxX4u9DD2DbXI/pNVM1QX/FsDY67etST+br3y5nCXRzhJTjqW7+XCW+TajVLCF4OsBYmqmWK
3BpOWELBuwPePX/65WKzNfmRi7q2GMYYQYxWXX807RBs3b8csgHDIAstNPbtvdcHOW+edz+6qxWM
ukh8jMV0qeLQbIDkFyUJgQEQO1t19QEoJSLEi/xDFs4R3XQW/jXViP0AZ627dIXmZnoVtqMYdFwO
7BupDA5pD/q/ERmp4+y6uq5MEEiO9t79Qplkbj79MkUUyCPbPbKiIFZy+PEl3rJYVMvOKD7Aa6MQ
6CR1sbe4RX5SUF2TBU47dPnPdcXyc/v7/TxmvofPOiRq9AsLTsBlasQiTCMQcsJV16Qcyj2y7dJQ
FBA+orU8G1pWSyVxfoHw7dK92tVzRqDtKVia5ycpPjp4EGzEvncy9WU1mu16X51QNcsYcrdc7Ekn
ZFe7CqXpRmUXS4Fc59wYDimM+2kuobDwZI2g36OH51FxVjtHkGumQ/5w9KMo0iR98opJpgjuYwUB
6UgBFeMB6joFQjPuZeoY+HaDJd65OLg3bq3XtK1zgjhY6Llg3DCw4CAgdng68TSJnSbO1HkNO/aH
4SasKTW4TfL6v7rt8AGaioScJwUC0ivIZvxG2p0/U+sbZaUqElHrcEB2o8srp9lXV4fE7DNP8PlW
NboBrX9UZ09kxmJhKKHNj7l7430MKDQM3xeGpn5SXIqSRk8m1zjwUgYdY8f23+9pB3DPTjxOuteg
C7VV9A6JOP4WGlzVM/h2M1gtxap4iU/xu27cB3dQ1H3CdSb6LJ9tYjjdO9dGH77W5+jSazuRUeAk
KdCvpD40Ai+OVOx98ziWLA34BOkG9+Pm2sKoIyassysv04KpEdrNerqMp61NgdjB//FPaSycGXPt
SHc8ePral2dH9zvaWHwZ9eOTPXCBn7qXtNLGxvYnQQjohSj91sQDOa+0WLkXQ17GUhzLIryZn/Ou
IfmLMHabHy+ZI9woMgC7ttFrzIyLtu57bVYZz2SJDTOBqoCVRGpNYh65NtJ2sMbbW0UX4e/7v8LJ
pqPgazYGJ9fbT0H2ijR/E72rzftVjGq/mj4RAtuOphfHGAsjrqHHvEeDJk5gz/CieDTCk0f2vMN4
nysRcDo3CXAbn2HBNzopaj0ASLe6+883Y/MFwRRMQq4KveWCOh/LJ4tZoaJzMNl1BGw8CFMT6bM9
aOgmFVyDxCfa441oCZXhXePeELU+b8C+sPze7q4JeZVW9crnLlfXazAYyRoUm75r6+r4JH74IslT
bIkY/i4UrY7hz/BhugArgMFMpPHRe5zPLnNTlrgCqc6pHZzr3MW4X83YDoP0Sdg6qqjl6qhwPyQY
kNvV9dhFRCnnOyqxmn0hWv6JRiRj8Rv04CEGoGnoHEcAb2Sa+W3iYjm9MCO9kFZZFXZg0w76Y71X
6cocs0uTfpyz7l9Wtl6wCgajWO4cXPf8Uofgj3O4XAdUEyR+bidrOJZGBoHCAhYR9qPl7FEhJCoa
kIRM/MlZVCCwdNfGIW21MQq/qK+xQZerP00Lruur8jsKxBfJ49tK2dLiCKYfLN04NJghb/O48YnK
otP/RVJDyGmP/XaO+l3mT3YVc+0HtTSN23DK5WMSlmVEpzVAh3Vv3DYpIjt0q21vPylN8hoeXZBI
sABe9qBQ8+H+Jrqrg++XKSuk5INADud8LBDclYTZetvSOfEaypRYKi1LXviNEcIo0W7ZtEQIgSwW
+tSS9QdZdoVsNOP4Lb1fy+ZttczINSSBJXvkPB2zhnBIufLYKLKTbbC5H8QAbkLWeFwnIOxFh7n9
PnxoXKzfuSm+Z2OPCysYeQs+eM7DqUI3aie5HSRJ5tj4tid3W1m4J4rwwnXnEBwvumXM5n2dHUUn
k4wect+VXPKmJHIxaUDvdjE8wOM20J8HscdANdevIlVuZKMuw7pvZnH9mebFp3l1B+FUxPiIvMRz
Dkv8Jc+2ftr++F/obdSZN19kuDnAmwDux6dLUpHVR+g+1X3zD9WJcT9NR2A1rJaM5ICc7ulkVG6L
OKiP9a3rdOgYBBqZyvWCPPCLXTUR/Rzj/8AGryz+YNdC0dM/19li/+bZ4cY/eQhyCC1pUPgj5pWt
6uFJd8YBIX7Fmm0GOfAhhQidxyCJNacVSSxwgyc6Ag6sVOcP/usa6wacIWYb+RqXgrwPPy26ewju
V67DqVNr2i9t4smfMket1XTR0wZ5k0i9khSu3O+Ugtdvzfk1VPgP/5F0NLo8yq7Npk7zMgFVP2FU
Dq26lqGOGYk8wpSYTTL6u8fCAVN0Im+5MCnVoPFinecjcgHPh22GcCD+Fsi0WZ+RieIDW/dPePH/
UjRbhP9q9ZWzjLDcebsRfLvl5fiktW/ioRgglHLF756l3mlcmG/VZ18UYuzJepwvlI7Tr2UcSQgh
ofeM1AbQLYmwf3u5SYFr1oelQErfwIPO/TE7eqjQR1okMOqbZW5mKLZRnbArlDwrAOOYHvuPPmPV
Wqopf71otsDFm+gyonfS4hPkccButUxgmaTAbJ4f7ueUOOArjXy/EYHBrU3TaFzFFQeqI9mCVTck
8Uyen1BQ5qusrd2JQnLsxK50ETZKOIbqZjPprej80DKjBmYXAD4khTxDpSFLNYDPgP7Xx4fyKh6t
bQkAf8JyLJG8L7YT9Ru14nk7exIXp6yAyFP0f9DHQHDxMi/wunp7i2qvF2rGdVPe5FE2cGO/COqF
1fwRMJbYkHbmuqLs8IOUZa6aA/hFoXiVSuYQCeyHR7TlVdSWkHlWS95Dv+lf9fP/LOoK5zhBzp8u
lFdC9gOLmhfF3PxnkonGULrHGGGzxSpaCLu4zmJCOIzRY4a9JVGjSJrph2WJnqoFdw5i8J2cwHNB
HIt0WOh+jY6TTJUf6DhNR94BiPUxlDbUWueuK2w9lFTkDjpswhEPbN+eaX6WWHSPGv8UDmLpu1R4
pmXGEeETwyWRHPBD5qpwo/7Y1PTcykRtiudRNj9kesT9LDBYV7u7aRC4rD0joSPgstRXoD/hEYNi
U/kUzRoluwr+qcpr9HgmNOsAyrEdzRuDLz81xCH/wfrXFBte0Bly102wQIU5jyOGorp5DOiqnNWd
DBWDbnsnUegZlQmHZJ7BuFIzSeEY/XI07egMa55A/9iBGLtYmCq9P6/iOm8n/HRGq1bJYGdubuAt
X4Q522z9xDp1lUnL4YU57rrDjL9x43BSsvcOChm2sAV3UEGYM/EH+59hPCwqOoMQ72NkWImMZzRu
UKe+s5q2cuaDU5ZTYK7y7M/xAwxsUzML/UamL8yz7xoyJTmno6snrSjX5pQTWQwpQcBpvS/0f/J4
4TwcOcQv+Fo1/p3qPGDJXe2tpkbOErR8+FSusJR/LFjZXl8ZBZXksE+wopzswpNdsI/a8+4UXMGM
lVAVptCwB7kwSl50qP5yAABpuZPInIQLeEz9AcFnZ2cknHivWzdoTxRFj9rFgxzS8z+IALNvav5N
O3w8Dsq/Ul+M1jnUBsI+aAB5NIun8CtI/xXKIaI0jicXvR9B4Ckss+UY7oISJTUD+hD61AZ3AYXI
X+6bO9Hh6hqEb9U4N2xXBUcXkXvcdrKhOwMgB6/8K1dXqvTA2UxnHTnO5sUeaxyOiSqzCyOOgshA
Xk56sRthBZ7DmLHyG/4MjkG427+IaMdfbGoTN9tBnMUhYo0tqKMd59Hxsbhpk9hNhf+vp7q/V4de
Tod0knLlBYrQqzmdfmcUbd98HyGJcGuaB+ybUXnWm12BBi5YgGYRY1dPXXDH942XCHcrv5UezHVo
cQOGsqfo/UbkmRupV5S2qnpx5nyn1/tGGgKNvwLx7XCrR5fjXEnSAgUdXM9MgG2+MpRZURbPdOaC
eGBgR+z/jrFJdfuoTZ/7E9q6j00V35kCj/0cjPHBCchXh0eIJj4Nmswu8frAqsV7rr6IsugdJB4E
Mks6Z5qoQOl5hqMak/1eLjVwYLrmlEcznQR41u2gnO8XNWbOtVLwd5vJKJyjEJoj7IUCn+/fBJeu
sHzTp9sGYE4abycyiQbxyK7A5MaA/ybJLch0GY0+qbTRHdyES35XzvuiwWx06LRLi/3Gh4M/92ob
Fn6+qz3WUTE2zUvTsxHhkUU+Kb/NCIbVBU2o7abLceSEZZcvUngMN4SVCkf4CPEP7firG+B4Cwa9
QJsYmo79p4oWSXdeoTMk3CPfOLh45V/YLdJPHFtY47NiKpFIVsZcvLqPnohvyNnLsAO6kOrdv3Lg
wwxkyzIlzrL+6LUJ/QLNA7aPox2Ay4w+ZBKyjXzNKl2sX0rVEwwBc+TfUjt1VDDugjnideDXmCGu
MBvAoOBv5EfKXEWFSfsuEx4Gv6W0h6Wr7OiyGJPIvR33av2MgeTT56PvMfbosSja3mAlFrERgTPB
fPisd8KTD2iZNuBXAlzghOBgvKFPgpjV2p4QUyo+jlRobp8WCfjCs1ng2amOTTB9G8JUR7vb9m6l
Jvx+H+1oI3fJJcGAADPNDWIMsi+ZEypbE+02pWRg1e2LTluntN6/xmli+9XVoB4FdqDyzASBoFxp
R0P6oFh4FFawDJXDq3cYUPQQQcGRiz4UvqrKBH13Qw73bFwhv9PdMvVrAnmOJamuNQGAeq/UtpgT
JIpy/Qy0wEnGeUfY2eeAxag2sT75bRUSPs5AO0weQMf+b1Yz7oBbMDmC2nrDAqof1jzWxsgIIEqH
RlmdOrOtghQL5tjgPUhAhmTs5ZYpSUDlpvNIuRBAXzLBcBlQCcYndVs8F972x7I1ij5PiLdFVOGl
Anj1PfTRfTBM4DpOTKlzw5oXFb02CMa3Z1LBSjnSxr40SUTSoLQQf5iZHpAyGNiqhrkjucdGikVe
K+9Ku1ANebnvmKTGckbbEAIPqQn3EsTfdm9xaAMq5o5V2BrHrAkV+XP49nnmQxkF1db7bFOxBNy7
cLpI+KVMEHI6dAoiJs9UdPVBqgsueGGVfFFumhSM+ZAz41Pi9RwG5r0D1+0oj3uqdB/alO6oqau4
SB32Mmm3EcdjyJqDezRad/LDaiDjZkcy5ARKZuFH3SLehScVn89hu4fRy9ErJDQGkwdkS3dhWhtw
uptJEuMNMNrtUwjMSRiQ0Aas/NuUFZRRQ04vZKbmhBR286Rh8iJbQnodGRge/fzLa2WzsZDmM8M4
i4SSjDk5orsOXt/S6kMpR2DwDpJOQhmUFqbBe9Wujfx7kCtb31h2+AVimNe6uTPe7/R/BUekadjF
WrdMuADWCRwg4Zo+LeKymY+isfH76Yjj2d4vYd9mL5/upwxjxnLxvmcWvRXSAj7flFflOO9OFT5A
mBlYe4mpuWDosmbRiW7/bR7rSjpuQ1Uobfes8jlLXdl69HbnxDuR2asKbDje8SGu3nt8dQtsZs51
PXnSr7xajZbYiOo7bQn+n6BmaASSaIKAHNl0SKYwI/7fOJp4y0eAZMtyTD0c4YQ9irKzRV8DoG/O
sQLHJfGyBZbKy8zNesvFidtDNZXk0bJ1MG4kdHheWvA+Orlu3hpnscw1cN8eRI8ZV2G7BdMnOr6w
lWOGo29hyRE64BHzSNyN6/dCPUYKKcnRCP+mHnMRffUzzzdQLfgsKX0s9tYFlIh2FQAUKZhVMbaS
ZDlVQDtbMKe1eyZbXWLj3kLp7VPZo9qfyRB9hBZoau+lXGgRJRzUOxwLvczUKsOK7BapsDChtQ4z
E7mnkXLBuVkZ7iT/Hk8WB+PDyV91zVnxKfNeZeWLJETbaoXl7sqShemPJOBGAo+iCY8zGnZDnvlm
XVBiu+fblgAfnzJKywwRLuU8oUHLfSFZ8Rq44jUXdTg52LgC5HsgSxc9dlNKATYA8sT5gqH9oY64
M3YozNYbmQpOeBTkMkUVLYDCtm/arGZVvF6w1OZxZ4o5Laj/0qNjUAIPijwu7X5pKw6DeMSjdVtl
ezlk5xs8utnRJ+OJVrGTCN2JWxhX76FEOyoWy0pvifIg3hzeZFIE7yRyfoD1NOcsN5PTPjfgxcds
HLnUg3kjIFkOJX1qjy/G5sF33h/ixwIZHQ24uOhEOEWDTS4OQQYJjYKe6t6DkiinqNKnHAniYnG2
FIKye7aQbLpmxOVd4uYFdK4PcnK1uTNOM5+CZylza5YfC6C6kfxSWmuV9rAO4+B3pOsdwaSQGeJC
5N+FYb4lyhRaKuS5sfjk9chPJJl+TXhQBKs+TpDOreWtmbncpPJD4xrKPaLGl9gOxlUV9VcZEenD
Tc7dIU/k+CgxUuVq8oKpyHBbzfuQ76yWgnt3wKmctke/+bYVnf6Q26hbABltzjNTszUIBOEglir9
Zdm8BqjAXLafT0bcnrrsms0aeS9HX9SP9/+pm/mKDcANZwNPdh6MttdXSpCoIJDrQkieOQkm0Qj2
7CX7kX6C9S+agND0Mp+CEWE7iFrZRa7HnRsm8kb1dOy6b34cmQk0jLiSk4KmyzkNIPGebCKI9Uy2
pVQeEAsb/FEr8rXDaO8wkVNHirbD8/2eMwslG938J9xd8chEiQtjKoRnzjXStN0hQLNj//+CufLu
631SS6tOJJdnulhl/TcQUWfLyxm5JbkI1+nlHF8mdtIpfk4H6VuAoliZAVnnt/L8e/Gu9KX7Whz8
Kwnj0TZXkj/58wvRMNy2SE781WBEelK8rhKjw1gLSrWDSUw9v2gOcNw0POXLocWigF1xRic4z6yF
Et73/C9gBzQiYfKq2pDFmDRXofpZW4zeKXRJLWgT/Nuw2w6UpBwofIhkCaG4ESkS+oDPpaPNTMg8
mUd+HD8Ogn5+f3+MbY6h6Tz4KUhacTnWgHY8QdHiZn28zVuFzK//wmlQpCWIAiozfPPPnF5n0xEv
6F8imYkC+eE4IjOm6sWMWZKg+AGjXugCipHDrao76InsH6h8s/QwaTewY+Qz3BLPqrjNr0YG/AxM
viXamfDF9u0HjSONtIZIK5/DYCJRexZsiJOh6djVmrrHUMCoLz3j6XLE8fLZSllunee1juN9PKcq
6RB2fv2MSLm2gdg4z6LJYxwjKY2Oucsyr4m8n9MUOviC9tJOUlNLKRXtuQeD7ZVx8NiImzr1s7Xw
OjtAiWpXBytfSvwp+BftHg8rUKCY4TIMBW4muEaWGjX7frXThKqeoQ+OWKKOWpPmEdtBXlq+hvD1
nU9Mif5aTL+Iygk9mEl1K15jLR8Vnlhfomg6DzdaOMvAslKhybicBvFf5QDdN7C7Tc5E1r3BfRaB
mcn/1PodiTJoojV5D78g6gR2RL+q3xvhMRdZRV97DTrW9WWjQWfHXGw2olI8Xf2hJBbIhNVWYi1d
Wa68EyLtZU+T5ACsOETGnvkVgHW7sl26agtrp/v2wB4uJqxOEpFIZaw/KS70EjV+jYrivPCB0Qg+
Ckql60NZQ/JRzUXQ7RJULSouWhoalKyqa6RuEdaRBOohKip/UxDmzCRjtNn9d+afrPIg+n+0cBkP
75DoiGWpZQtUu69JUXtRHAQhldv05H9M19yV7YCPzAW2XedOoAVo69TiKlLlaRfj1ZIPjM/SVcOy
obTiUfdyXoosMi0aRe7fUdShc2DSOd/LreFtwC/2KMhXGLjIgzNbrYMil7uwJkm+52IipP3N+EKM
yGBgzrTCCptFhoR7WHxSaLnqxYn6qkn49xba7qEtG4QEPeTkInaldaJ3Ivhm+EkYo6y5cu4hZQF9
YEvzuvR27OcZepusauqNlvMEQ4k/WH9mWjYpsRhwgsQNM3BvOG7KEAG5APEp0hOy/UXuWj8C5RGk
1p0uxhEu3+LavgmKeZaakxqm931BfubnrgNK8P2Q3HYZU3ehliVQ9+y8FMf60q1w6s6X0Y0GSYvP
mzmw0/+HDVBvZg2XdDVp2INawe8AzaHxyDRja9WO8+H2+b+9y7CE8iTMkor21lzwNQc49oiA3D8h
WO6OPja2T0FuBgbQ5xgZWB2g9bby+M4l2T4Iud2P9hdJbZuJaFnFowxNrzyNl0lSKmSZPKFD7yj5
avd0Iv4qAz8MlVxgU3Y/TFoS+LYKB4n8rQ9g/DSAuOYBbfyMnQ1kOcG5JcmyZrVSJjxC8fF10zeF
37Vwwat6xlN8s6VfqyFA/7zghCtPGLlE5HcIWgezI+L0501AqjU9gqUQ4+bMd1vjh98D404oHdZK
YnY9iVfha8m66hg4JvhulhnuQ0ClZ56rThY5+geUHDHBLxVL5H5cOHKQLayQMLgxG3ON0W2OeZHy
bFdS5wae+JPCDELwUrMSoC6XUtXm0RDLd6XQZsW6X8Bj5ITfMTkTZbYBlDjU/7aXuqdMOTRcqTAu
CUMeWHv0Yg84eoDntuj0/uLmi5KPSVsAgk9wpxD/sAHT70kxBPC5MXrDEbz2xx1qmsC3weSvDjVh
Wz3B5g+j6MhfyhGnAH2I99KvMxP+HmoFFUW3F0MUAs6VHY6VGjKSD4b2YH5XxFI+iSeg4hwyzViW
UlKVFINU18rqVzGOK2exwY08fcvpptKbT0pGcCaQyjg2XwIKpR7anGy6IDk26u5gmNVi0oDdDpea
dNmisVqhNT9yaxBvTGZZlL4Br/zwBg1ayUp1FLvQ4/R0m2ABGQ2qUbFGKSUChaF1Hl/A5mOgYys0
nWt9lwU+bf8yg1ar2nyuRboy2wroQ6nVfDTwzD3Qlnn7K2MQLyO57Mi+0huqHeecfHviP/Tztg5e
uiKM354LLRlwXLlIxCmsNpsXqcvc+3Av7uHSAG7SJG5AL3rA+NQY1zY/VjJeuJXSyfToNqQUiJIc
HhJv0eXn70mOoTOK5K9FTy+9kPBXKfhVllqD4Wst2CkaR493WLAOlohIb/ih6kl7UAv+XsYS+caS
YkU1qrC8laBE77CIDw/LeVZMJ1HGCH5EuS50v0qt7uBMUAL+J/VY9E9T/gUZkEJp93WDHgPf3RLY
wswOAXfwGcM1JIEqkjqurOAP37DwfhXZIY0/8c7E2Evc15AtIB2cARCDCupNBjxm/sOQpbdduwkU
pOjX8p5jv3sdF5+W435BsbsihcuRIbX98ljLsNhLKb/kvyXec/mbjGtbJtDsI17T4rj16xq9gABv
UPLNzam/BL6NloGIk52jhhvKfA/ciArCtfWSlgY05KcQSmQF8sm7NupjJvR6NPYOzZL8rXWrsRvg
JWyudPHpIX+4G8Av//MJGQF/NA4LXOX8hotmtDHJax8k7x8rupwePL5cTcMKJjwiEajZmJm+6OIA
bCEBPQQXe0T4ba2nU0zWme67NlUB1YAqkwE9JxZikO3o8xsL6o/02dQp3hyVlQHmCfE/urNoT97l
ocpvKD+zMbpOIbEXaA4PZbvNW13KhOrHYmeEFqHW4uPiGjyDdZ+1m2kgtRsGJA+I7NNjLm6MgX0S
/Ugr5qfC9rNOfqUTKraTITeL16yhGtkXCHdlnJmgilQgi5dbIY/tSV3n+AxxrmMyWSQQ2vRoSvTU
Iku1NNiKCPtrBkL7D2IYyaWI/N0tWyXREmXHulYJRdjA8UMb5WP0eomoj4hSZOIxqhPztCb0iUGF
gIyid+/qCPmbIem8U7ZRDVVsPmAyZ08wyQ4QbN3GpqsdcmxLj0oRSMwK7C2RrBjGWi6TrJEpZgqO
di8KOxP1MTdziuPTMj26aZaizu38TbQvrxIwy/Hna8XPGdvcuC7SKmXOFNK/clF0K1Elj+5hr921
Q1p+DhDB5DWZEk2SPSTeKKwaGP480KnbZe0+qztduQw1Uap50oUn+UH1lWhYwCOBYwsY3SaKKBAP
1QEHEPnQMzpTuomT9/EFgk8d5sW46PiNv6En7TEMXdxS9phppdFTbgjYHydXjJFaylcGjMtolXMJ
PgepPC/C96FXXaiKDan1KhDmrI9YMMyZqvhpM1b7vvLN2itjIP0pG/dI/OU5UC2XDjyMeua/IzcY
LZ8J/U0Z913wAu3KlG+pb3QgzhoOdbVChU8ivO4gAbp1mmEKy7/tYe/5H6Wo5omACRYsYipdmi0S
NurAgp+21TW/Hh7gKk7CAcWfdf9NaJcTzO2WmbTUh0aT9XCJc9ENUdo3Pok5VC4rMgbMPuFaXkKF
ka1mRKnVeYz4g1FuOSb5T3wQLZgZ5njiWQoaBt4CKWwaHEGAmmoCnNrhntIYmqCO3Iuf4WMoEmLt
jNRMdqDlG9Fj92jTEbkvzOmDPkfI34nNAQnjeXRlTxMrE8yVheyNonzBOgAnYnpGCs4JZwUnWtmQ
Y4m6H2oAdClUjByfTRSft89f9flC5IZwilUtPRA/j455uJsuIHYv5i1DoFPao19hLMAqVDDjnKoL
qKX0hKda4Smkw9fk8Ni1cLGdm2Vsf29uqFVNRTKtRdjNC9wwLGBnl1QctfgDy5PG0fg491kZBnj6
BqkzOtw6Wv0e9gwDj6XfDoTn3J23msHMlTH7E94AukSGk2rZWfYNP2RMa+HOnmIEaYyV8gNylW4I
w7qJqyfhGvmLFcm0p2yL85A8xZB7ogY2xt04wmIbaFPHLYEOUYm9UXWZ5C+rSoIUxbswphcwzH7g
mEQpGOxsqVT+Eu8bu7MKAEWPjJ7pt2VzBwEpuTD4rusMcmRvINXniz4YG987NxGFUMowyqRzxSwV
24Ni+iBZlaUbrf7JaL+m8RQLsWMMXqbZ5C+ubdVjWRCXTxbFdQYQYzD++ZjT0l0nLAZXpBWH99nH
fmhawxslNc5paL7J5nOE3t6GlJpKavsmXCr+mrmDQoqabTmb4gQkqpz/SI0VKkMyPQcQ82eymRhY
fzByGZLEX9DPrlJcY3qulCLc60IRlXIDQFhiUWQXVddH+XHXFmlJVsbZLaP7ZNQTam3I/j5WTu/S
q2O76ILhb2Kq9/dGpH86tsJYdwMYGGN2e14R/CyaB+qqvOLu+9Ha4ymyY69qNaye53kQ3nn6N33+
5YlwBr9ISvpZ9tLp/ugo6m9f/DcxXgS+S2AN+UfRKChNQEk46jsI1EvsIzf+YBnAmyGcc8NOyWcj
opkKThfDPKJe+/mnTT8Z9aOoONjZMc0iA9LWjHKAVOxHzdRFf3HXy5SO39YY3t547GulvkWaaYII
i0sr+6yOh8U72DUHCElPHvNgtb0jzKd1WtI9iiKz+Eb7NDKBv/AS9gwiJrSHoV3Gl29X9V8bHcmX
HY1oUDcZC6uCcuFKS2ZADjdY0Wl1UVzxQUNPKIkn0vI9ony8kzQkC7aHpu6lA5Uynl5EMF+Yqg7g
brRfNfoVPUJdkjClkMT6Zpl0va38wB1hxtheESn0SlV4SXMHwmEAdBE/M39GjRjk1gWXqHuVSoko
Ha12vNOyX/6xxU6h9rEvPr5JIJBI6uVdyqtKRcgmNdBP5bKrb3irmCXbcK3ACe8G224I22DC9g1k
lWD6X/JE3ShYwfymr9QpSiqjgsKtnzixDTpx5d3K2xauxXGMJQ7ULKmTfOnK29+xHTCzWq6JZf3I
1o2PLQ/WTX7H0nY11pesX1sxETIL+ykF/IU6YMpHTuExGqxOvzncNC4Cv6lqxY9KpyNv+Sg1cWn/
GvPa2m4uZyNT3BSAL9MMtymyPZf6/6xvSrR5bpalRjzE4l2nn0tAbvc2GygpARjMA007WFwZ1laE
fuL4sVLr09ASYXkETi/VPuPiHybGeScGVNLh8SF6IEMXcCkJDNpOxBh4uQr98poP8aQv5PLxDWaf
ow7R6At1kMQoriG+m5gWVXfBeyhmEONLu6gH8d72ULv1SDcewJBPNiVYLaD8gmFf/G7KRrckhW6q
/8VHkbqv7yIpOhSZGZdRnywdwqSkutX0DH1tXWLG53c5XCtrPuvx6a7Y5QTThNcjkOoRrhQciPZ9
0fEmZRn22zu+1pxkMBc73DGYEyzKF+GXiWqk28dpP3ZdhgR3NO5yri++7n6+PvzMmFs4eyv2TEH3
noJMMgbxLZBm48wmMUH1740V9h65orbWyH+RHtV4CAOi1awVumAhbnn3nqZL/wT+SbctkLJi3FpP
jLkVKn+RNGosgGMUcbH+0Kbf0fsC+xAJ/Tnsshx5c4UBjd2sm1YlDRJY/pB+iJTCIQdS7dGnF8lz
dbgY/eNoyn1YX/oLxtuQWoTgMDFF/8N3JZD2HCZw8vzO1C/fna80I/2a70igT+plSTmaFEION1S6
72hx/MNauQ2MVtiMYS0TVCRvozQMBbh3l2TZwdKZ5HkmFX58rJLdAQ3fTosEUEAqPNyOFiJJkmpF
WJcAfMKVP84o0RVadsRzS5kD2A65wPKyvAKoRXm+baNnAKIneZwzAE/Y3SbsL68WgiQ/BLj+QSVY
r0dLqy58sblU06qqSYACX9Na/yrhcA2Ydo8DQQehRTTOFH02MlCstQbmUe8nQGJtGnKo7VcqgvAC
YVWrf4P3Qt84oWJFVypqAJA93qMoyTBco9J4m6Rr6wDoPmFDbHf8NWI8yoy646DUWEzVmgjbMXSK
H5cPBJLvY1LuWByGmOe5i6pssBjnZ1IITBDrhRKFY6Q8Bas+c/zUHBd/YALFUPl/vxJ3dGxaoAcT
3QsKBn37HPovQWLe8RPOiEjItjH4RRqwzZR1yfo7EshFvw5w8I9en/JDuCbNh8VBu35c94N2VMxF
ICN1ox1RxpVjbTqSec1+tAly//iEet2XMdoDAMZyoFg6Rm6WmoqVDrYLKcDE60y8gjzqfW1fy8fo
qm77Oy3lmgwPS8PHg4sFCs6bXNP+4QNj7lJvcVLNGGU2VCkbnbQK+r/L8kWFC/gWSY41umLx/8Km
hcFFsHn3Z4n814V7CX89v/kTD5Bq4Dcz4+0b0S6qwCWqCPtrQ7dFwlBiItX/3GtYJnGk/T4L/ddt
smFLld6U/L50TRhEtvZORwLRuoNjS2G9oQR/9dpB2/5uvLkbhxRJiN0uwFEwemNHoK2sbbOeDBZM
Mby1v7dgj2qk+pxjYD5Xygzot/B9SZSt7tknUPlAIBg+zGruhGaNdtMoBsiqNqtZj9QbH+nYKS3y
ToWS2+OFJpN4IcCubneqqr/X39F0/l++SJ6wU+stwp9G1+8jEcY67cbfaeazRLnVcTJWJMD8utnY
GOyZECZ/tfYzQAwtgma6z/YoXTJAPxKmHZhpo5y3NauFOtFcgtPJvAIpXwHJfmUlJZdjG6VYUnCW
01GTaJPLr99/Rs7ulGz8zvMuHQgP6DBAQ+uxWrZBcF+wbJrizfwk3/w5C/sOzpMuhwKa4gHiqCgs
+dweaKbrZGGr0HPCPaJ9ph+vNxE9WnmcEfDIis1QARnMF0als8xOwmwiQBiHDJQcsXpGwXSH+93B
DYVJPe7MH9y4o4q15rEsfsGCatZMjUc/ucfzJC3XEnoRzM5rZEOEPLUvon5bmUPCs54S/5KqZhSN
quifAHjRm89YbwLvnwHnMKBgZocOHam8NqtWjQLt3fo9MKLz3nVPdYJq6yQrrBySp/MrVGs5jH5q
0OYIssIKxZNmWhwL2sJ60X7miZgULhqCfX12ZavKYrGsJUFvLNQivhTJiNgdhlq9G1lngtNMFM2A
DjbVfyb92J92X5J9B8kKNNJkKhv65xHV+lJAJSaf7vJQ/AErqrmJONkmsmzbwJ/DawDN2w6UNJCp
Xz72nTXAfJU/eOG2kdk4N6m6aR+i0uhms3AwFVQWkAdiLtNvRqi3PQMsc6BuzUsbo33g/LSvFWtK
Xx3TX7x9MBmgT+PmbJCzHfdXTI0c+Dua6Ul1uiXtrfQ+C6Uj2sszYeB3XPFIuy9udKKMV8c19aqD
Q7c779jy2bE0zxoTAGaY3PpyUE8Z2B0XASDVvOgtVU3/afVinMcQOrCpzAOiri8uOFkBckSWNQTw
wq6Vcaca7DcyTRROsJDD8GrJaFeDlCSoTKft+llRDyzPosJjLoxAvbzk2Yx0dUSVIz9/yLa/kIRs
mLHm1azdzpQWFUPrQ8FDS+VCFsEIc2JA/lyJo+MrWHPzeX5gU9QFq6lmEP2rmp0l0wkDUr4t1l3A
azekxfwTF0E2rCoX4IAkCrub1J/rSRA5UYq3XRwR1UYCN33O/WDzMk8FmbDkgd8umjb0MsZGgDzs
w7tLu18tKuMcLK3clDmLiel+nQSVrBQjJVmrPU/TOzWGMiIR5VE4z7Nl+RHP5bt4kcQBV5DDIlJv
asTIxM7A4cky3MjYa4OybQzcmNcKhJfnGb6gk/uCYS1yJc/8LrNqFs0U0akIpyBEzKh5K6ODNJav
/MZ3u8tv6cSUc9A19BGFJ2HaHNfQAlizkKkHgumgjwwvaEnuMaD7A6AxQEzST3R4BHQD8ICfW2cn
Sw53u20oIjxKHiF4FpUjBIkWgmZuIvIGQinBxWdjZV+VucrxXHIy32fzOBliZbac3m6xHq37RB7Q
AcVwLlP5G4zi3C+a3FgAafRmLPb6Y1amQi3C4/tkgAsD6UkgyUve5G4ACifqNUsLQYbR2xR+96an
wNoYF+PjrrP1acWWiv6jvpPg5todYqdHdta0Y3jJ0PsSZ4XUMcy5SB/VAiu5+EbD8N3s/hb3IbzB
EBxkNK7jh2ZphmPwkdKg+xsumeNjKpnR8PAjYb0XmueG0xIIFKPHFuhaiITYLOEjEjEa9C881YgP
AKJz4jikdKCK0xT12KydUwIRHLvMGJVnuHALE29DiKrSAY2cr0WwSCpCon7Jhl0BuwyqRgB1LZEM
FDl5T848GB+fm0BfhjGGlqWyWyLg9gcN7iRIfZ1aspbaYULtO4hdYR0i0tUnczUdPEhNzZRYnNS7
d3Eu0vTSmpSzsmqm06WmeWg1aZZOuFkMuPnv8vzHX0WSH4X08DYGaZtOu0d8JftoD/louwZF0sLb
05eLp8lHjhqslC/KdoGCS82PjCy9nxwCcXMB7nNiiXZFiBWWTNkJhhKxRFDXkzk2A3cU2LVb2MRp
tiliVACfZm1RN/TcrhSeNH90Wq/sg74F0BAzyX/w7WjZLHns8jotVXy9+gpVdxzAJcG4SkCs//y6
/0Cu22pOLj1DQRFddRirD8dUfJi2ihSiZ1hY/6NJjCWjamclimR4M6DCuD8cdOVBiZLAnotnEqfr
YeOKGNFveafM1IiyF2JXIiRIgVUeFgIx0Kwx148N6FDmHF+Cvkr4UDuWAC2uM4gBg/EUu7QVJDy+
Sh7bM9EDV+968fyuCC3zQtQhYjczE0RYEL6cZRfrjABBltxOiAUuCKiDOmZa0rRaktKTkuhvWAcP
RELtJAtvM6sgXrpk7LpyO4QO9rkWPWTM54x5898e7f2WzoV7ixbfN3BA/UAer3B1JmeqlTAEmp2m
01nZ4RSi15E02oC/wpJrUV4QX3kvy44jnCFXMu1EaSC3599E40dTtVqOoeF6UCu+ddvAcRnxdlr7
x7ciHtKEsHBF/wO83AG7k5ymNKAtVqNg+E3ZA+CMvz5VK3vO7SVLv8rJygVoOUTH6DjPRONNI0jh
g/U6/1la+HBAkK1QLUkh3r2MNMakxzXtMCZSMyoEWXlpmWZFge7ZSPOE4fFMLzSRf73XuJg0PfHF
c1dY3jmGbobMVmwdtMKhSGl2QmoPTFAuY1YydOUFctuqv3fFkkcnjsEsRgYEM5+fORw3fjDnO4l5
BdVExcEmeH5QDdTTxo3s/VO9RR1QhMshy47XCxlFW7y3QPiDASq5vbnc/iwMHxAkzFyjcvHX6oLt
+S/C0NdHxHbw9Xi90ry4lWaCelbqaZ0SlZ78FawnLG95h9tzdd7kYWzRq+Xbwx+QexyC6iRjwR9e
zaMgZelZv6RIPFl+RVJBwtjZPtEwFRyzo24LjMONzwilDuL80EavR3ZpDaeLe2S7jdPWEZB0cDPW
DXaTNm68Gv1TLxLzGGVSExdbF+WjS/Ug3RZto769ULu8axx1tab6b+MwVtzMiVjEQEOSYAQugCIg
4ckUuURW3J58ZGt+EMUO/EySD+VeRxQQskm7YKSvgmkmKBmcTCheKxJhz41adLeaJY1YS24X/R1j
OGAPGGGV+YvZ3WmYqONC6fAR2qaVZRYiil13m2fw9sgS3vBkdKP18s3bmsiKlo9hl+FQg38BcpCd
KI9Hkg9L+knYH5KpV16arOIpFheO3oQxmOSak4k9EgYrft7AfqBfZs0knPU8IRStSgoyUzPp6tYO
j7Qnj0ri442xu7SHyNLod+c4uiTt3eYAK9qSRMWa8u8ODexksCizXTy/ztunVcoJewBOXUcYEdfw
UoeqbDQSTb9p2cLKQ4JXns/4V31v1lgs+LAG4SorQK1g0C6u4NY80cnvBOvMFo8yQxtao0Ua8SRP
I3+kl3tolZmTH++43VL1Uc5fPLimcOeh37+9c1s8ohNtqoneX0PoP72owjA7S5dg8DhpR/kQQ4O5
rfR6pXLwXd/AvC6rHy3kFuiDncJ6xGonEinJe1dzF4X5UUkYutgNuZMunTadjE9qmTBozQdUyv39
jUdasasMj7bzVJ/ff6SzPMZq0/Fh4DGJEPISgEct0dTRSUcXLCMXpKYb52N6NbInU2gh9zEmtOFi
/y0LqZdmkRqmpjxSblnYn45YGXuYb6OcLaBrSNg1vF0Sv0l9XdWmsOda2XwGVwWEOL5Yf5yadV3l
dQE0gRPJG8xJCDHF/HLR+wSTGojV94ifI7psABQBdg82AlLTCcFaxdFXD09ssNYjVpCEfzmi+rph
yMrayul+rBNQRHsvCQfBjG2jJP3UuS6z1J0bwVGPheWNMoWbLIBb1dH3o+IZ/oGbvOzj9+c4nGTa
MhqY89+1o1YRtpUvRRn3YrTCEu4LWoGWIihVFxYom3hTYPy7w4cGRWEpKxWWZV9Xp2TZUEdN1s0E
gAogKEkkPUCtiwbPogCBl4uz0i/pnZT1a+BCDos+ZCaQPiTLvOpsx26XQEGdnIAwrE2tChuqjiTR
Bs/fQuXYMS9vemOmSwQUOhaA/B5boNx0uy9xXwpEikz6eAYYdJar/U5UxHnHBvd7YonBCIm9vaqw
+5kHC2Modq1yBhSvqf1vySuAMpBAd5mWHiz/fJf/A8gJ6C7u4+pIaDONHMiJ0yrDVZCnzaHFYgXa
UOjwpsuaqTMuXOOGs5jPl4xaI0UNSGWlbdOLKhrCAHFIMOaxUIUqnWfODA/1rcPIwTJiMAN/6Oa4
rbf5EMNQgc9RTybMsJXP6p3du+nUcB1EZN/TGqwhHCebMpyKwDCeCRf+EFVOeZyvFeqQincuCunr
yPtuUvzLU5C5yWDJxI+8ZUTjnTjvKIYRSP5FjO0+RSKG1hDLDTd2s/Nm0t15BI42ogSi6vSEiPMK
7GSaVVSuJ/l9Pkq/Nn5o1CXG0ZNJ0ABnFzvtv2LRf7YtgC6W4U7HGcgUkqgRCfLdkM25oMUiEsLH
HZBCWP6PyxMFfI8s9u7GqOHG8YH/SRA7zbZkKFKOTzomTE3Atq/oU4utec4bt+8iUi2IUDzdqwOO
UO6Uw5HW76qcPzxZ2HgdTKVEB0vA31xDEKV/dCxylnEu3sztKmN6Ou963OhQSEzjDgK4zGpDt/bi
0a25V64e/NxA3tFiTpWzFol4xvyTgtQoBFtJHKGPkI4vLe5ZuhlfQXxziY9YNAxkSVcCfxrMj+gX
auN2JKTQZ4L0qOxKSOp8oj1zVl4WvPOoUIPwgFDsXos2FsfxijRWYm8LtkJoEntPELe6kGIuzmZe
/k5H+Q7Zp6ZNN1FGG3+3CABeLI9jgi11IKl7IqIOBr6Nkza38FIIyUrd/HkZiEFWyhC9jQdKKgEn
lZqZbdP7W1kMsrljw6mYJDRhRYQC8f97/hHRMX1essD9harHeHw3aONKOFShJgHJy/PjO7Urdvo7
f0vo7vP9cs1dra30EOFzgjW7JnKDGID74UH+yHl/O5cs0ImKIjh9tpGHQx/fpJcujBeGC0MVc4KY
Ci5h8e90VhxMRiL3Ic1j0f8TJ+mKQeux3U95G3aQ4ZZkqlzUQPUqr3GBEiHMnLi2z4LnXuAR0maN
6HI9tSjKZrKx8XW8au11RL3CfmUmD+JTALJXYm3wEvCiyYhTI7ENDY2MfpuLRRxFuT/5vPz4oPk+
csn6IkMY1ZQU4/EvsV5lvdLzb7b46VqHTqDucPV57vjcvfAY6lbG3g3TN9wIGTW5Ul7Gq+0CvlU0
I4Y2x3Az4pCTT33yAk9tj0whmGqUInc0pBM2vpdOv2JWVpZlnRF+NJ6SvP7CKTFIuJYtZqV9hAx+
JTcQeoulnpeFy1x+u/unpGiEn9921gfHY4MrSQWmS6DS0lXVz0ZW7KCgQIpCbGqHtajN2dXWiNKx
mbtFNTJ3aqOYMiMSLHIH4WjJlARR0W+Ejy9Ihn6itZYFvYgcdlGCacvOTww8MhBuEOKNxVki0hqd
wdqRq9ttqbDl0oZAcvVHDf230VFbWTjZ/57XoQsI6WV/CodJbggt4mlNqIePR6+MFQnlTjDYgQEx
2svOLwIrZqkfkjmFLcDHqP4k73x2AkAKlAx3X45T88yxmhoPT9kuG8Oeiki4lIZjJyqZwmOCuur5
ttLZOTv1Y4T24D90rAYgBSp9SWIY4z3pwjfPzXfLp+ahCraC6cTIGorkpzyXiTSKho484PiM8a3O
Bo1BwRvWPweUYjnbSoTE58KDD2hhEGx0Rn3dQ1VQTwEDnkFKMp1lilgxGtlrb/mJagd/HaFpC43v
QN04pVP4AsvFcPA5OFd8/8h9QIABDzYXy4irhy++Zbxzkufxhi6edKMWnI2fWka6bf66lL6p47mC
uKK9O7c2XErwYsotR54OxGMUc+moIgUObBZgm4VeXUIU0F7Njv5XHZFwmxEC/atuLdPxRTy6YxRr
TFZy+wbq7PYj2FwvkkWgIWP/KbG5IFewX7R87yTVJBo50hh2GuQW1fikRB4JFaWgZ/c2s/wJJ6SX
b/ljSErnk/yi6+1oiDcEOt56kpxBxX79bd/RcWlB4JTaAjAC3G3efMShQGxJbdlvbszXt1+Htynk
T7PK+8qJwYu1yz4d/x1i0Tb8eocPUQXPoGFa1IRc3cB3VBshwMIbF8P9ZXNonF8gwGEX9n0aOSOQ
5RvI9SExvhHIWnQYxo8rjb0HqrpF6WgsK0dqVkWyEaZdrl598aS3o8TWKzwp2yMRdZo4VZCm56cE
bkw42MqKu/PB64CXtduIWpVAMgEhgKwGtw8xtO7k8MvGCSDt13X0etA+i7G7tocl86rD3QMnNCkF
dyEIymejxOML+gnp6Q8S0+rIRepEPK5CjW3Vvgflx8/DxDwy0v4SthKMUpBA4+B/b3YaeLL793zC
oVD1/85s2JFGGySKsVbSfnvdZUCthobIzKOExr9FayyOhI6dHSterPNkL2i3EYVokaq4Id0UQlRp
SB20fzeRK5wZCx7tfqRktdYUv6glYU3Ac3FGNWQMyjei4AZBxnBIddp7i8qds9ezl9ciS4YakjHv
cZiU+iZCmXTt8pU94NBCXynkK60CPi4QCE742XIngwC5Ivs1IvVO//PyNxbDxULuf/rm6pExrewg
72YfKCy/RQxkBnfRWSyAwnOBK1KxDuwLtZzcZDYF805cmDE6/yQZ0+hk9EVTQxw8msEqcV5WGPmb
kDd/WaZaTjtNR8HXumlIB+RNjQb9ziuWH+VOzVs5foUzHz/OVTLDAbOic2IJHvZXGZQYUHVwDRYp
V7WD0A/BiRvTL3lTJ2FsAdNmRq4eCjIvddicDGt59mWiM8AwFV7z2xdPqDKDQoletvdDM+/rb9Nz
iTI8ODUK9ISr28HTOts2FFFvXxAbbLxI2ZNtvEvGk3cC/3Xovt2j2FEFf7NanenWwMMGmJB+A7e0
Uce0y8jOrDu/oUIEXHzxyVuAK80ngJOxnWGKWPmM3RefdSO1SlM3weMG+1B5YiwRP86EBRNMeXBv
j+mw5D/D/QyVILYpfjqWIczDavLTnZ9RjX5hpLx+HGf1UpzKkcs6I9/SJ+KhH4t0iD2jmgakzos/
gSSnC6VjOOyQP8Gjb03t/uzU4E0HJ2o3vAM9NTIeF8ukh0Htjs878QTeyjXtXnxtRF9+UGXMFBzf
sRlhoi6zc7Y/XN9EvoZcO0g4BuaCQw4o/yVLeaE5a5Y/RL7H+HnUy3FAzUMmzlPE36NiLPc41Z1g
3YrFCqnjR0ZH9LZ8mwWx4Iu5JuMF8rIp7XkVjBVqC/nr/HzCwOTTtYjlxtHtUpuDljaWLwiwJnPi
Oi+zz+fiSedMRBJGAc9qSr2m+eoQYFqFM9jq5ptmt3skMa/eB3sJiqxZhFtZeqOcMqJNquhtzOmC
uTO8aBaV7hPvPYuYtvWu5fZ9yh4hHonIA+W8Jl6yjrwOXZOOSGT/Gh1H/YN5Xn4cBmclxYMThB0a
qYdGpK8DXNQp1ejQ9GqKt75RBTFWXB9IS9U5lFQm5LfO4x6ALP54cFsEBE/Z7WH6bxLpI4/Z1iE7
j9luD3YevHtHujPYmfLTxnFgBmlhsmhi6ROtHVP0uURpAR3txMtQY1zlWJcWedAQDySZMtbd12o+
BZNO+Wuct9ls8iaxYAAzQgs7cldxqNhA0iTb26y/bFqcW/5deluaerEvtO+C0Ic6dqt3xS8P7XKH
2nxbjw9AyqTMlbU2dTufhw2Anqgpdti5eybTKo4Cr3Iqzyx7mIHiU39CkNP+W3bBcGdmsqihKhF8
ZeAo1QV+Q3Me1tClYUm9qzC6iNSxDu9OiY2hfEpKThevK/aJO5G1IKoCrzpe1a4eb/Q8qqyK1UuN
fE2C+ML4OP5QVT2t+h7b3lYRUCGk5HanzfY8y65eeIwf8AjGL6RAU0nQ2VcCV74WxlfV05TkbLUX
TCoTCd1hV4jGw8ZQQTVVycy1Z5YiJrrC2yvCSFOVwKKE882Oy1NpACl563gmeERyNK0GhYu13B8J
IK8HyDib1Fj+KS1FZK7j30AJ1pkTsYfjpJu7UPmIIUIRT3fS3TiDn1ntKppCm1TdtiFwNpYSBT62
uvh2g3EFOaLmopUgi7nRm/ynd/PSiMlwZBCuUpRtuwRCFs2YTTwanTscm6Bwft9fdTYZ4RRC2+va
yXd+F/p3Qcv6S4f+440c64rq87aartcw8eWwVLoZot8sFNg8d3+F3yUjPsWXNzeVdJaNgqj/fdMq
K6hcHsZNx0BPUDIlzQVOLMse6bRZNKgr4TFvPluYQ7vxBEsRGUMEgRMZ0yvxYUR8wzecwssIhuBw
jpzWHbp1Pn6xHK4jqTbuc4TGtz50lst7CH36BDQNR4dsokdkyxKEfOF/jqLIB/XKp4lURxBy8FuV
wVz9tFfRT0jEhkWHIQqZNSYT8nnXPDcWG9w7bK64kGI+UFFSt3uWQwV8b4+1eVhdRa5diO6aswfS
lsBGmOldS94WRciJQ63OCVJo/Ym7PI+W6+vkOUoZHlr4ojr3W8RbWJ7KxgZhCjMGd1MOC806+5wD
KRulg8yVxHs2Yg0wGsfhKBAcuqhm4dnMT6p7tqzSIuzAU+SKDJ3IZXZDysBHBr3b5hK6At0pvz7D
S8/NQTrMGvmgq10ghMdGjFsQPj6vuIa43EZCN8YgHjegQC0zx7WQchSfDCkEDPvXwHb+0rKEK1ZU
P+d7Whj/BgsMAsy0wAQaKZdEcxKsQIYNRn/HUR5fKAGRkF2Avtblzy28wVWBX9unBnyM21+mkC3D
UW2dUee3CFOYygJS0aIcuJ5gRR2isW/q4Je0sfTZP1pMDJTW278hXvwtlMW6W+7OLUimKm48Nlfn
X75aWC02sUjMGnKxgXkQZiSQj0SYQpQ2WxMnmBphvVqHkw+/1QFVSP0c5B0Y5tLbD0Qtp9TIGeeR
jgNO6/6g6Zkm3ujabkfhS1e2nCxxz/SRjd1aFXh4BDy2z6p7R+brc4yYnWXVEPH2R2a1k7ShySl8
WmykEWOXwKB/pCJMZXuB/Lul+pp5+ixAM8NQ/bsvbMnZzEJdXgiNZZTmqxyQFo2Oogon7W1Clwq8
hVUZjtKgwFpuc49VY8zqIoZsiSvZABkYgPLQUqdQjySlj9mwI55yTaYIRUdOO98EFAcwNqGpYYjC
xbOZSE5dZKGfKKSPcHoB4th9n54arVWLM7i78EDMJrYYWFunal2TiGnHVIC5tBwe3FlHRxyWmryF
ump3IkYxMb/LPWKRr5vqA5sUPBcoI/3QF9HO3aVTccI3EqYTR2QYXIEksi+jDbkaz+F53Il9cPwl
BCv3PqJU9oDlbOl6rRe25kvlPVAdggmVrTlCpFBUTQHddNIOhreQQCXEEU45HY5Si8TCmB1nes5V
Ogz5VJLgXcpglaShAOQ4p/QaWK5kjbcAaNsnuxv0DiwbW8Ag6S7pLu6Naccwk2fQ5ezEUhBXnl6Y
RzQXXFfuYaDnv1bu7ZcovET71meeiYOAtKquuZsEcAIrmUZ/T1BVl0NJh81XJ8BHDF7ZmB4l4trd
e53Tm3Mlmg032KTeODyek838Rf2th9OQAaj0y86iw4miblM/Yg0ytgzxSL/ZXfDKgc3BHH9qwd4J
iA2OsoIIXMwtUYNkIfzbEHdI/HPvmlrUWCIHBDQRb88XDiJfGOrJ9nl2tqqOQBgn/TKJAtlKanSO
SAC2zm02azKlUPnNqgFUNfstmgLmmQYD/6I23FFoxkKL2+md5subdXJKpQsuzMZ9AI7gLmb1TKEj
bLL9DD9JCxf4mlGDF9SNwq6Zj3G7IWLm2F8/B4uG+Lo3JgeP5q0KVZWsUAmslVRj0sidty2CxN9+
ygAHcDiAm8jE8w92T/1F828AjH0v94vETooAj+dj0SLRo5Eb9Rwj56WJ+F87KsfnnmRAXrnoP3iz
NLIO0AlOyJjxo94iI7c7kw521Yh5R2rJHl4kOW0x7WsARV9mLCXlCP5BrT6+NZIg9RRPGeOnKb08
qNTYtO726v9Q6LIMA8kfY/VaGJsX9Ar/bvVzzO8U/K0THdfpB4NAb4POKN8c/aYCO5kuOrmNX9QQ
dv0TjzWumtOZA98aQws2eoCiQOxB20fNcyVMps8dFg+bb6t/7UeLZAnwNTIWHbdg7HEXuhYrCCeP
jVnWxxn/LL/VMj7G23EqOTol6XwrE3ZFMj9UoDKdwruqcW1yXe8UO7XRt3buVNkXsmb7JawKic9Q
fshe0UNMdmc7C7olPnsNJh4aa3K+sfyIr+R6sJBgTjRnsEYfRHZArKYulT4rzlk8fXJEGakIN3Qo
WIJKwAhJRJJz0NIuBmho/LtsyKG+n+CotS5ZXf93FOXFxmZln0Ub+n9WQ0EqDrizaWJT0o0QKxXw
e6RqMuxYnOpZ/85QSSBQ6jxnahLFcBKCCf38fsh9InARdi2DrcQaBM/LBeg+yY5emq7jW9okYQ2o
HirWWKrrR8M6BDoasS0shLw/9FHMnOfAX+1CzIBdntfC7z5Lh66FiBxb6yb0Ysqsvj2f9jKs0tM+
QkQ2EELaNAcF295G8eort7z91OKUNsfzuaUJAKwnaPbAy3t/XUNvqznIfEdxP/qwSGSPyKJfBosc
J9IMok3UWGxtv5r/WgY1yMbtvf25Lb15eV/eyxxl5xU/cO1l41UYa3vLPYw5DsRTMDDkAjk3rkoJ
kunXWm4JsAuRqT0FrHWS5Ty/sF9CVAoxDn6o9otrJcpgBvpPx6G75bo55nnqrLmfrGigN6DwA7q0
1c1BSIy+i93VK3UC4EuO6ApP9M6OVXFKv8Bfm8SfHpBm3YAyiXdLiGS5fnQGY0i7Se+MFr97S3G3
lpGde/pXMZ7IvBUEtEWeOsar1Dufs07tpct3K3LRkHWMV3W8DMjgF+C/FHsOAkFGEfgKrSlIhxrh
t6xK1Bk8Aok/tAEhJlI5r+rrw/Q4z3ozlr2uBRptfSdEFfYbq5+mM1uD3ivu6gTWKT0RRa8je2Zu
KASvm3W5A6ysot+eUisOa3iZsUzaDUv9zeuHl9894XD3Rm6p/QtQG0GT0H7q+05vyQrDxDEZCxaj
1wkB3QyMw/8/hjf9rjiPHUZAd0PlGtA9C+6AIKOaPvv8TME+t9Hs+tjnRUDVPtaTNF4EpRmUosyS
1qg+w6ouKWjhEXGG1R11Xq1ulrYa8JyqNTYy+2CHOHGTBIj2WllD+FFIcm5xFWNIftuLq3rRpDkS
ZAgFdlrrf0+3MyTe6zbqiN3rdClkQb0pEbAXnCD6qo7SW5sIHt0K2nofjl2ZQWqxoqnO0s6ekqZB
zi4OX+bbl2Af0DdKbFoFYPSQYt+yI0U8Vc6jxABhgsZZm+NWHCiefwZlqSD6tl9N1OcRosTi+3z2
NAvxXhJRqHVeSwQJlzsf66v1Ehn80TW6AHrAXuSIvyqYGCr6sVYOWi0BbDKlH5x+EKAhosWrPD9y
lq5wAFIpz3Rf4veKtW+P2jUCXZzV2QDkP/6Fn/ego3JDRXHheEm6Fu1nyH2kyvlBzzmt7raEq08g
yn/wfG0X7nIKJA5G92HyHiUHW1V/aXvxH5dcsJQIQ0JILtchvURNQytapBzLSkAplImNtLt8k1Tu
BCaMadXDwld/Y+RnLVkoixuzoFUfWf0BOfeDJQAePmRFbHqiveE4CPvTPT7Op+5Q7Qp2biqA6rE6
pqzr1prdGeJ/VBT3jNGboKoJrdm0Y4wNws+3R8Mk5hoM0wqX09XJ9kwzKiuGBPGZlSeD7cA2MFnl
cBfth+Y5mJE++w//tJ26hOxuFWO13AYLnfTFbE7GsyzAngepbbQn7xDDqdn55GdSr/WXrXsyGMks
00j8SoFTR21x1F9esmoT+WnEvTBLISgPCkH/SeYEY5kaZsAQnE6jqbLoA+8ZphK81nQMhS2RDH8H
qlUiO7AUqKrkKblyudLuMkUNo5yRlqDTyPKwRzCq4efRafXbiOSMtmt6XFAQKSAA7ePnbKIcGU47
tqRNY1ykGriocRHiU1h9XHAUCjjV678QZzH2/PGrB3n+/9fJZu/nwFD0SWfiHOb60TXtFZPzU6MO
ayxf/Ll1f4cejg6WjaioLM/8QsPtM+IxQexgMRNEbmUz/91JJcTpHQGFHVP86hOvQus67FcBRf6+
UiloZokW7qeWzjzFCtpbLoTYILASYCNY13L5JkVCffHMJ2Kzno6SaCF3RBz8GU6ma+c916+2Jcij
VfN9eD8/ZaG9TS+26NDuMr6SuEJHbi/Scia3TUyfuSnGEb97XQI0lFSD4IeNeTd83ZnAekYXmBND
sKMnopPQ2oe+lq0bJgFwr2TFKWdmeIf7zahoo4wFQjx1uYy69NzvcJcLtacMR5e+IcSbEhgZe6ad
f6PthqTcHWkBL7y2Sx6mQ2F2QnGPkrwDBFDgkKq2zM1pmZpeBRUkOOXCJ6VCTkuyZjpk9ZUGhleC
HA0Yr/r440+qhg3PUL4+Pbq292u/M/ln0c/uEwIGGqWCQCTceRgJG4LTT0KmuYn8+wXq3k90tVwF
eQFXr7+NMb4jUpEtz25ZCnQR6xuXE0zFimgTHlS5vveBPDYOWVMoiYyI/qXzlB5gMa7maQIYWbBk
wKX1/pZOvT9S2SY+Tr4WQpUrnHZyUQ7YZnOq9EvCaAJCgruoHUQnY6c8iZ6ZEulB/E3qEGZy1Z3W
4AO5py15LoI27/mP+LLDAKrkT5vEexbzkLqgCfM5VY3UIlAVM+RrEKnclsWovh7hcuX4HY2Ogdut
tYLvZ1icElvp43WP8mJlscjjabPLqc2npnx/O/P8VwjIGxpCjf14xsOf+E3vbSfaLU8Cmi7ed0aX
Dw5tgvNZTbXr+ZR5Oz8HBmwr3vnliJd5dpBql+tyHMJXNpOpOBE/ZokHizNlsYOB89lpqctmtTQN
OjNhf5Z1OEE8Rh917ttg8Q+Ec54m3+4D/4y+D/1bHS74IGn4iX491oV2RHaRrKOvCNHTlyIu/RZk
rrmXzpqojkcMKrkVRxyOUMZDWVf9JYzsTGOoxE7bawJKfUF+pjiAo1CueWXQ0U+KzXhMB63NZvEq
zxFY10OfvcNIap8jTGP2Jg94kLjzAmqI92Y6kO4+S8+FgR+vDsDTyHIbgqu/5d7bXWy3nyVtvmzy
ADlvBwFbP0/LpH2L7Rd/EMS1stLoKUMjzeyT0uKL0lWVckmf0QqP2lehBBFUazjevjKLZk2RJtub
8msqXV3Rh8hFU164mq2e1FphOzkw9XHq6/qh3ULbp39vWNSFLav4l2+DbEH94KN482gtNzlB1xpa
k36fMPUeCZMRTqwhDSqCcECZM7CCgXtzI0Q9GpN+CygqfJEm7UMaqDhaEq1U/+R8Q3mM7uaFg0++
OmB5TBrdhPvq75xNPO8NV/Be9LyvubDcxfWDJPQD1IkMrcERumXX+19mlaOdFQVrO9z0WsRmk08F
SL0eLyFUZM9q+LiLA0dG8jvMOvo+4XUB/7uulAPFva1D3YDCvg224as0jafP3vKKQGmtm8Vo4DZJ
NxfB93CN2SHfiMtdMePRGtMne605UpHrOcPn4fUwk45B+8i1gSU1KwDg3yq6bdKwJIjTTDgh58mp
8NssLw+EWL6dArbK9BQD5lYWJoIq+RyM0EOrlhjOeLK3Jjq737MAix9YoGlB/6eorkm1h4newVpp
Bkm2jVkuAP2mEnnjhZjJpjHMGMug77lHpA3ygwVc1elAaYHX7NCtyVkH5LW8ZWd15U1+41e38U8x
HdH5m8aDihp/BncOeJBbjXPsMO0pfYGYU+ZQ+xeq7Q/oYcMVVeYZFZJfUc/rMDTn9OmmIhgC7K4P
LC9QMZTEiiagurnHcgQ8SoE0JwCbmerBvXEW87W/OkLmLKunoPjIk2BIHDIR1XTV3H1xyi8w/+xP
SgP1uPoBorC5u060iziyuOFkaM10Q0IjdmXzsdKnyl+MFGRDnTRQKcGpWRljj7qGnxXZGY3BlFEt
oxRTIujAXxSe/YW9fVH+77NSWEQq+biWxIqrftwoEPQUn55/QAhKhhYQtHYC1PdgxkZzjpIqrRWJ
Jszkya6mk3+Gnl2GlcgF8fxD/MPeq5PCUaBj3le99cUrjUAJHHTBhPn4P7UmpmsuQjPYrqoggh6f
bYLQ0MuPJfwKMghRduOIpk0zbyQy9rThssiU8/N3GoDw/hKBQD8MGAqZILjKk6oMvVppKhSqAIuM
Ea5zbLAWpWscblmPfPom84VqCeH3G7BR+Me2x165v6o5ongflAtcDNqPtN4c+n0Bz0IjUO7Vu+hy
dSC0zLVvQt5YAwdQ46kxrjCcKJHzQ1vDlkZHXEF29jYRLsfW0U9JyXwaaiN39y9HILqXtDx1jfGI
V9dVgMCw/xh884EarSTs9yETlN2wBmiD860jvBAgQPsP9mQHSAq+PcUBAhKVMbqhFLu1Kd9U0H/K
ob1X7hrh4HMWMdO0vOo718XybBdKd2e0L3T6MvmCOL4OjqswZNfgM6BFWSF8HLfL0enSZFEvbNX9
23T4QYI6VXAsMfIJXgMvGvRNqozDwmXWPS5I6lKsLJ9XRdnRHKqTkcNGnZt3EDJGJ8oEI2FjAyv6
gsZse/H6GIK+CUf0yBB5VFSzk7USxlU8ny/SkumHV9yqCPmeXuhLQqdVCopeXeoB/wNnIa66O8wG
YcATwVvuS3jD3im9ihWQrxqfcf995szrmZSEWDpKifmLHZFp31I2ho8x3ntVp0nQs8VN3ntWXGf4
TFvJZ8g0Dj9qhFocaCUW+ijmq0hkczkxw0kuKlbLjMPdK5yjUUe0BPFc2zIHCcW6GUYjCTwNZKkb
HfDlyLyJhfkrMj/T/gmTwf6wsB3GOCwLfNr6HkAbDquh7LApSDMH7ZkKAfO3rxifQD3eCLUgdN5P
HNjhdHkmYX1vQW2kQYyPAsOQRbNoy0lScGyLMSb+yDoAs34bSf3VL45Amd5C2O4u5g/QKWqiZEM4
mSaSnvIfbNFTQA9SJQDwENW32Ka3h8hxE3kSYmLU3nX29KfjOgIFK+VnejD92b0S25q0tukIgZ2D
g0DGTD5pvsX7OiBS3JlGm+Gfc/FpldrGHF4WnZrs2daZigTpnj8yTVf6K3Qh54sNczzkglCxvl/Z
7gMrpho6FbykDto1fviJqpKPjlx/sQ/pAKCW/o4XPuuhjysWypETAnVx3HTT7lfe2O+r2PPO26GF
L4pwU4iNMfNyWF9aeNWrLPckxaSDXFXlEDd+pXsH7DmWHDwSDN0p9KHC2xUbSuPH8HdyqCB/WkIW
tIhsIfM5Xs8HmpvGrn++EooadqdxJmXlON39ykKIiKD744V5B9xmRZBmi2R8D/O5qidsqN/Ajy2T
IR5aY0O4g9odnrAIxR5Snb07p/XpcmbGYebt9Vo9Ic7py5o0Iko5K/KaBH5gyX1rF2R033aoieKO
RaQ2sYLUJiadfCCnyB0q7egFEsIBAav9VHqFg5ZrVmhWluTe6cc++9lvx5cJ1MPSG3TFU6KbEs3k
Nu3UQa8w6z3XXYgnZBsQV44cK5kdSz4/NlSlt+saSRvIJYteFmgsEjLhj6k66HNm1SIfUtNZvbL3
ygBmhIC65yDQ7oMW10CGQYxlW2kZB3ftoIEIEgrc0Eoy6nVmC23v9v3Z2wz/3mL87DvHSZQimPle
G12SHa6cwDy61IuxWxZ02JLu7cqkOWbFvzAf073EHvF1BrWz9/2jMvL633yqjw71f8m4kHlyU/mo
Ethaivfv96gH6e9qO7gAF2akEzqLg+Tl7EsOhPwcuK/V7F8vdAyKvuqQirufHXlghNYSQ+sfg26i
TFXPwTK+ClcXwUvs4q0Ny6OeQIXgDcOrAxc8xvUESDI02D9RgJ+BKVDK1ggeWMm3y7NRCIXk5/Pq
3kf95//EAYcakvJeRUrIy6sz6EYPnmBDssdN4fMVu3dy/k7y0lkNGAEE2dsmNIGkEL44oWG+yyqq
ySFC+FH5f4TntzSVhZYIPjP8QYqeFFFBBNuFZn+M9D5rZDawbM7IVyTO7JMJYmu6q47sbjXGSSS1
IbwK22l8b/xE0lZmKO+OpgSRBtwuWatLc6Iif0Vs+sVJsaIY8DXMpcYwUvmx6gHwGNnJPDpVUJXN
NajX9GOq7y3n9FPZW1RsXUvaCqQxaSeS6jBf13tlhh5I/tlKxQZjEuB3NgRdhVbKXNBt5Z1PoqTK
53/9o7ziwAaCRIRpO9fbtgZbdmFEejllndvvqN81Zb7lQJWfjlh646mszN/b479JemUzKxLIk2Pn
QD9XBi6fT5xnj7J0PgZVFwdMd9zj7ZTwB0GfWh86xUAq31CvlKmXMG0MpZZCkoycR7PXdglbZEAz
96IFamANMoN/Vfb1RXVNTaIXOB1Qdq4ulgtn0W05IytTQDmLgD+roMIkqRItOzOzGINMSWrXGCil
BZqEjDRagr3hLMo2LqZ2DDi5hjQgvC20vV9JXa0r0qTnISFoNKEyyaTSBCxldqVSLtnWZojBl/kW
jk1K7e/Na4U6SsQPPAaGuJQg/wf38qbs1eo6Nr0kE9yUlwJcAxBTM5iTooli6IE4x+kJSeLB4HLd
iH+l1TUycy1CD6Mln0Cz7LJMzS0HMVu/F56Aq5MNf5ON5+2VWcFFuH/3gLivmJEa2GBUblmodSau
/BZRqn+835f2ZExf7P3rp3wbr708EMVsp/k9JqkVC2lYP6Hj6ZUcWkgJ4K+ATBa27/HuPk1E8AVk
6RJVDErUm9YXpxzKBYUW9lTPKe9BEg6qY8iYNIcUro/orwSvHuR90h1jpF9T8xJ5uhskZ8gOKhdm
K1p0P6SkFsxHhWjh6sLbshRBQBuBpYgEE9c3MnA8o2HQ8Iqx89atFwF+DeEORrqR4kCR4Jtj6xle
TtL1570fq/ZXAg/temsBQ1su3eBmxQMpc4NhnjfssENnTBAmYu5gkjTD3jTHlKp4hRgAatF13xMa
iwjV4XnKSXsDI+QSwzGUoFO7PGhq7bO4L/IV8L40xUz8J5pAAEV7jfp433wAP9JUcjrRMIsienzq
hsFuL0fgXJ2E4f8FRGmgIHz4t6j50GQnZhrxXeRsZmDOiHIWeCamQh+qFElnI5fuZFfpJ4BILFix
XjZe4fqBeph90e4K+TcGrJ5FiGVHWuq/Q2h9aSmlyyqK1uVd8FxyT6w8reVZ110qFFI1UfbPXrRF
4dLQVs4yjZLRvuiigtFssjXWKgKAmuGIWQ10SZPYtAr8fgrftXM08pLwFiGaQIkv1gEElxballqk
Q+9VgW6FUlp0fKYq5stpCCC+oyjUQMXM8lG1Dz7+/62blvL6PusrJJrVM51FLgMKsErNPLa+PsfC
PqaLkpNW/FZKNuPnY3RV6FeWgwVOZQ+a/EdkrBjlAwfMxWkqTnljQCD+6ozuWBhaXhtwYRzWTYDV
9ywXaZlq0wplAPOpKn4+i1Z7rhv36xTgzNr4QzIPVA+Tx5kfSX9a7/VLC+RCpxGMeBnrVoVZsBnQ
njvB7nKD5YE5SD3mCZv+x2WKSb2oNw+EqbBthIcakM14OtjXVQzKbJX68BBEtL66rqGmlKU20tZi
GeQFHpEz9gLOu/MTUJQ6UMyZhPmXPk5YLp7CW1tmOnRpZ7X02q+enVzzAL9wrKT5yyCclC7OXjNn
EqYxEOb9tSb2iNZBmtfi3aHOhJRJndP5BIjCy9quyLXrFX0R6HRJkRFU8gfKSm0Xd2M0RnsxsXwT
swp8ja9F3PfXW/wNHOSvQFM13dVpr1liUtwoFbnBMQgao7hHkdlGjD1J/fjJwXOFICsPfpeyuCCu
bTnvqZHv1SLs32LdJbnj74Yj+Z6FnNL8AOZqmvnBpZh+IEPXDhRqhAjNVqlI2e6yCrO/OqsNPBPv
lewR1JMihhx9hU+kOy3PZMXOvipzgHXwkBvsC74Y9SKZ3HVBuCGHjKyISfupprQu/nqEPCJHSFJi
3qviCbH3yxGIiJlPtji9XE16213dUhcrLQ+y0fvxRd+wRV+xtyg7PdvoXagpcw2W2owRX3O+mUE+
YyJAjYoeuLHX23xWqvaMgk2H4VqaWvpqZi5ouaz2MlJXVAUjr/L/D23DJrgHtZAT3wNKx0NSThX+
I8zPr+PgAscDjo+ZPUlbzgJb6ZCdOOI7V2MP+YST6vmsKvs+8emXFYSOeTcUKo/I4cWJUHhby3mq
guSTKD61TYb2g78cfKzbBzAgCb2Z30in010H9x7jBMeu2x5YOeyl52Ojb2XtvkNR5SxBze11OmXX
LvvwQc7xO7ZdVogYLV9FBXd5qgaJvfrylekc/xSBewkGf0cuz8YEAyjJj76uvWAw5/vja6w7QPoZ
P29stcwXhFKSAfNLC3gIW0LREICc+VAthdqxm7n4LdjlnHGTvvw86Yb1ngll2Fm2MHOSaF7FbOyh
vNEL7uuzoS89MKR2RAPNNR3K5QDs39f1Ln4AN4nts7xCezglM4J1FtPaKfpIPK4T+w0OVVhRM9Ka
2X/LA0E8DaqOuzhaT4aWiGpGVmdK16AwI6huyQJgOFkYc3iapzk7K3CT3m/toG1uytn5GieE0Y6j
Wo0Ee2kM0x3G2tHWW9mXInyN8Cq9BqoiVyX4doda1JdsWigxzEcjM5iQf7+VyI7qyR1lsbDEEPkI
TyA/6W7aWLBiqkhOg5+Ns+duU6oUhDp0NXLWGoqfhyJcaiHfR3sqkQEJ8JO95QpFYZ4lPc84ueQ8
ny1rfwJmdfsWlFSI7dadrERzjFlrCHJ9ob6eyxazNV2CBJ6l//BT8C5q+jTB2xJlefQeW58urImy
yazfAupOqYE1mKpkGJ0TwTB6VAlQJS3wze6LN9t/I9ROwmLOXeAaXMY/i/DvmPSl1FKZpCIrMlLJ
MQjNoVsWeSlev+Tm4nf3hpnOQ+ZGDKQAbAT0V9j/KH2zQAYXNy/cKttDBSG93nnzw7BiANB4u/He
Tig+JVm2ODE542Y1IX0qCxCKpnH3rWcJh8E5ElM3WPbGzZ5LfyuAsRR1JulWn9z6Z7OvIlXI9UHL
k60LXfENDTmoXHXEDMtf7M0f9Pdc3txtGmeZkUtBJ4/f15nNfuzogJplWZXyzZGV0b3LoFllL92i
dDvMPSr1YJM9iYgvQaIY83R5WUQKrjOcd4Au8lgfPQUKfBL++ZwKl+9LOqPGzWuziXFHhFlEZ6m4
O40gb3lTpnHoJ5KTMQn03CgB+43Uee8ALVR3iXjvhMERkigP6Xgdn26CHDs4J7ZhDnMepobIMaR4
vsf7BBUiU9kB8UQNNJGKQMtQHoIui/ynElH+IywskXkpPI3e3S19239vFUAdnu6nVIsSJQxvKd10
ClewZw6Q6RrRcAqyBo6asqziQSrpn54zGSDXiWDTsuOZ77zaTASyF5tdfUfz8TPMaLfKVwdAzwkM
Lcgo4mFdS6iefY/DGbv4R9VJ9NXPXPHXTFz/VdKHzGdXRHwXfAwQVH6MrDqBiFMBH+E6FSwbBWNE
0eq4skP4NHf9NjC/YKlMDO3RwV4xprCl9j3otAhQ4+3iJTgkMiWACI6WF+nBkzJ42OO1vKHjNNH4
v8eUboIS/S2KY0pxhAZhPvkRaGEvhToafbHdT1s9yzcOU5eIQrOlm5nwBla5MZG/4wk0sVnetJE5
nMiQfCrnKlJy7x87XZ92oXTm3loOGajk5rY9BT7cGAFR3g4xzcqBs5VW4eyPI2yWoiZ6L+98GdY2
toEVoNZhtxADVYcaLWmOso4a3Y1ZkQp/Vbm4CQxnP4pxrNmnzA+NDdMrzBYjBsj061oqQZfwEOSp
GVQMVE9cqMOkLVazMXp15SJmbssb3y2fka43zh0XtfC/h+ZQYFHtQD6zi9iHIT9TkKfs8GkO1yY2
VmKKTw+yjYhO2pvL7jdpCGwuErAYJeAlP7zlcVa15BXH5eLm86W4ft5xR5/SaPuu1Xruonw1xQS6
5JJy+Cau/G8uuswVQYcxccpWabeauXGbmElVtNBbyVlJLbw0ue/sh8bwtKQduVTKY6xBJqpB3usO
9hPjnrFt6nA4/xwr6KAu/2Vxc+YAFFKTQxM4qkx8JHylFdvPkEKoAxBamDwJccVqALN3rSH47gQJ
GJsNILvY1TJtb3eUFHzg2RQlV50cxZE6d8B7dj9VgpK5AQjJJX0diWcsPSlybzB4J7YvM7jG3Mbb
hTDL/m8fwK43gL7Uh4KEstMtts+Ug27PXvGYgu1h41hX0ss+wGq5Ja7y7Le7jhYlioBUgIuZydWh
cmapl588DH2OkEKX9dXpBAMUM6WNUBDyYQZxzEOugEbX01xW2ugfYDkjWtWZjRSNyQno1e5n2Aym
ONhJKDSYULZhEstt3anAZZdth45xF4qvdFFsCwUeLaJdNJosVM3UA+A6PZS5ZU3herhbRg3qriFo
06AQJzQ9JtC8i2zmvs3uEUG1s/GLLwvbhNgL+934qb2uXzcb7txR92v+Awj6wbmtVc5XDSQeyDK3
D3377j07bDYRF6IDNDdYodbHl/SFT0JaAt2YY8zheCn1SX0GAZjTn/9bJeFTvurVVTHtNi6oQkxP
1a32Pd+pieL1jd748E+OyDcF4mhycw7dF0FSZA4pmSVSfXjrs/eIdtqSr4JxIt6kv2M5w0POm2PS
FDpjak7gwmMSxm1cafr/ELaifdZq4nip0Q2DPDRSaxBkoY1RL6KBLeKeYPbHBiaa3cxz9ztMUAS7
BjI4BMzP4PZd8fb03SqdaWjwa2lD/u+msXU7V/CEKvCwzMjqveNHQH5oh1qkjAUKW0zzzuk0TMJW
HXlpzAIQWccztmBEiuQMOoHieAsJfoowJ0Mg3pOGkVLj+DYXsS1hkxvaqXdhtJwgv5v7PhCBpgyY
7/o4QnpunrJdCu2KCOxTH4pekadQIic7nqUITfMzD9XOFsVlMeURKtnYNUYNd42Nzuf5H+GOXESz
qURMI0LddC+D9B1zYNJw+kyk9l3SGE1wh3/Bm1skPWxYNf7SBUTXHW33Gt063Q/I21OgJbUKRfYl
hpE0w7dCFPpDfyoMDViwDmvhC9DDs/W7nl/PLmT+8CgsDmRkUo1M5YjBMp7kI73QTM22OJqU51Y2
5cKW30ia5BBeqe45I7LXoNjAiy04qi06jY+bp3+uOmz9VtKqIJLtaIf5oIJX92NmTQzsO3+RukN/
N8tWjJyjEySI7FpDde9Hf7AFbcuztV7vWw4/2gvM8ax/ajI265FtHnSDjxrCMvv8yc9j/yzPXlE/
eNpgCKffIJnNuBIgGX+XJmd+jdBSqup0VMC/V8ufL0VeRiOFJ+pSQyRN39n0uvYv64pFsc/Rvh3Q
tWJ6GLHYBJsU7Z/oXkB/OQ7c2+KgFCCEnqM8DZKnTWCu7UDqWS/rrnz5VwCNp5vxWKZJpUBV5OAL
kVe4oq8PlgnQgLmbAFTjEzPdPCQDX7wGbpL8un39b4htsZU1DL9B0Sf47fUwZIocdDRlxhq1XRbD
0ujKy0fTIUd4PgSAYIprnvJePpxlSATCtJKt2cwXTqEI42TodVSZc87GgB+oQozG89t4aI9Yqp+4
1UWm2JOZ5nMw72MEMD2Rk6DluTWT6rtvMW/Kto4BK3HbH0/aYAEQ2Gq/AFAoS+aMZiGdo+6xDxdM
T6u1mrh8QJXApDSCOLXeIFwz4JapdaoIo1DQlOC1vCsg4kkCsN7HjYW6jSTrm4I5hi6mNVGC2n5/
3+P6IzgUUrB8OGUJkLy+6rZS/sCWJxNg/fFjhgM3AD1tqMb7X7DO6dR/YNO1I3llKMoWh9VHShGb
129DISBfOvWr42dZ1PkebDnIiJCS46EhCEaBD4P1gfClSGCEvt3Wgl7uaJGU30wyvhOkLCLDaqT1
y7v7l/2jPd/ouvcteXwAqKYBC+XgEMEh4EaBMO+LlttatC014xnDtHqRMtwIem27HY250EQeyJi/
aDE9tMSrxZ0xP3XaRKVLnyt7qJ67IBwwxuHTxg3/EONGmMeQBmB89qGhzKEhKgigfbWA+N5+S+Ue
1hPT8Ec1lVFDgLTnRv4JMvO1YisSKIRVXDOEiFvHel7G9fp94XNrC4Wkb6UiQWkh7HtpjgAscgB5
WO6P9yf+ThigkvNvyEMqy7Tft0ojOkBPY4OnSfePnHsaoXUHKS7hTWv/hd+pCBqj8zzmcbeDaLUa
GqJgxgqvKnUvHhbYIcqsjca/ltK8GbpRvQkfApsErTHrZt6gVQ3/2glHHTpKKyGFJ+uoOOQXnhx3
9tGyR8x7UhQeSRU851LVF5158mJhI+lvpCFd1lLxfx3H5zaZWFGnCEPxXRtYyQsERfGUeB4/hH+W
gZfoM2tsvg8I1sG4+cJ1ms27dDe+jS3Z81tBvY1kFswVCVR781BMZ7VPnOLfWAQjm/wGaHCuoLht
YECTUdV5Pp2ww85Cq8oNUKYrj6paT6U1XuBAxWVJs/hSHQtsbylgCAf33GKuPoKxJuKkd9q5Kr9W
URGeyD1QCXqMqBnmtxoznwF5Oc+D1Y0jvAvxw1sLrtIC9lON7Df+8qTBYYw1K7qGCSqu/wrq4bIt
b+LOpr1MS//yBYuB3n5+guTaKajs3LEqc56A8xH3CzXdOBvnmbnlzLCXmyx+vlFG5GQyzVfhYyG7
yGRr8VSfW1tI1vlFb/9Hh3i1inuAD1ER69VNzilHcjE6clOwUVuiIaRoCllyRAbY0q8yd/ZqG+mh
ygXcP02OGUTmZVpv9x8MCFXHabfDN1Y3DLdjbz3ReNKw7gXaWJRqrbA/lzDC1FpfEMDr4Xj9D9Qj
u+UR7i7YHHKfl5hJ26lKvcxkhxWF7Lqw6P/+BPdI1mfDqGPHp21pZEValuf20mZgHgIX4DmikShz
eFS/7c908TufpTnSp4wevyhguX/r6OXX8mgKBV0inS/idbB/XO4oGSJeBCWaN1nz7aQgFMViWI41
b3i/7V/s+c7XD5wAIXfgBYMwcQOPeIk3d1absTJl0R9vE7CXytATd8s3uj3zj3I+NFhvWUQ/xiT4
rucvHhjPD4xc/zrYkX0llD1E1kIcd7xOnobn6ZSBjEytuNFW7RUCuj6hLAqqxZKIUdR2v4PjqamR
X82AlIMnjQxzGpbOnZ/dPdkTEp59kAww6pWJMdvVDiEM8YsW8jrPcDuzknPJ4w9Xlw7ZaMX1xASR
227avmGFfqdurA2JULH/yqZ8XcXgUGFHPuv/BSnWcDuCZIe0Xxq9HJXyI3aDjERUJxft7eAsF97H
jt3FtCrNijeYCfdo39tuR8cjU++n+/eDF9w08L2xu92vXxwq4SwbTKMLrrsY1mJU3qGQ8ELmQj61
SRzCl7jvSxz6WGOZ3dLDMXwFdi/Z7Lf1r4CoJZHTjxrEfqBtNtYzfjHybXWnsMl5VWnh6i8yhgtI
deOqvf0MHKT8O1pdBfyY6HhOGxsN975ycgm8x7B26B4pBeih9yEkPfnmbpPnjOuiwWqEi3e7aW2o
mCl8nEg90IDH33agG90pOGQGaTYhMwPSBEZOKdEbqhvUJbhZ3pcQkmIyO/cdOVh+fXtw7nkg0fJt
fn74wtF6qXzDgFrakp5f2oJzV0jMLqTezjMidcYExelygJ3Siu5W0b9unxkukykBDBrHuIccJ2f5
fMD6ovAIr64JS5+ulDO53xRke+MX7EkyFTDE9WJqNQB8J3DoIbDyNA+24efsn0dQBwVnMAvHIFys
e6SCf9p/SwaIeRIuWrRgdNATQzYoyDaH/5dxidzWz7ZHcDK0++hrIHqfdInHXoaczV1hNazbPfm/
g/HMVFEOhXhADkLHXFUzzG6ZM0VUyZHVxnXntBIR5gPSoywAJjOhdC28lb5m8T7uUSDaIw4hO3ec
+3AebkrJ5KZHAsXRQ0OBM/EZQxJz4EkZWTzbmVnlovHNGvEIaehgwCyhTxF0ARsvRT/opF0owR0n
22uvSAYWgA40ZMnXLrSNyukRJyxipRD5YUTszJnK79LtJjJi9bgqj4NmzUAyWTQFrxx170Z4XoYJ
9PDI6yt5t19e6RYmf/odJolm7vtrrh/Aq4PjVfRX05Z8bm868/dNjN4Pk1Qia9U6sJcYNxpGn0Rf
9IIgfwJWRiSPDoGFAAqfzMf8sHT4BOStu+A4zbnC6069ZVxs0AzZ+Q+RMoj7xiL+sBJTmWAyD9di
UZxEJfvHI2eCzhXBKTDM2h4GTTTa9gwuIEMettVl8DncIvPIj2C8rEz31TaxdZMDLZcoCEyEHdGY
/Xkau/Flg3onB259CpmcMppjbL00SGrcG5lQ8qF+dizbt/AiZRtpGZfOn9xZQre8u9KqHm4593ws
c1TJtj8noaSwUFRGalWL660E59EfFzKv5fqkc+836o+BpnXvLg2QGAoPIQ3bLlekwOQOsO52fuVw
vwHdAasHsiYDulCIxm89ePp5/mhbrjvi4YvAUEq3slQs/uQYSqsTfF/qx6C6OtAQW6sEGK+E5v0c
xwUJYdk05yR45T7MPW9D++WLnXgfrcrzCLWTsKKz4/7ieU8ZivEoaS8A2ILbMM3jzkWEZXAcTeMy
k+e+A5C17qBrP1tTDZhUhZWvZYEZu0RC46DDgrILQjNvp1wAOZKlN5YJuWQTjNeQftra2uysDhqZ
Z4/SvgiTO0XYLGlKDUDBhS4IooXGNEBn7GtJu2j1vrogKH3dQcYCf0FZWp+JrONMvhLpCBWlbE5m
LSVGRJ/yIi0gpjFH6ncVY4/YFgiSLAVV7jT6FN0PdCn23jne8rOn6c0ExezJVircDVGgGZ6cmzO8
efCvB71Vc3DkTmO5Z6ac1HaRkSLSpSGzY/ZdBgMvmSf7Yqlx/IVZeJXHzKYq9B92+qAcWNSI0+Vd
LWX9IrbzwvbbK7YLDO0B8hXl9y5UzIIF3sqipxQSEKWQlIIP1J9ozGKk02XvRe9clNAnELAyT8EO
BCjjcD0erGDH4hZ/MOHarX26Rv4fEO+c7EyRWFpYHduGhT+++gzntUZ0MPjea3jaRsrJOE1C0Ugi
AZ9JDlYMU7Yr4nIPAb2nA2TeJEOecAl8N7WUzpxF1l4XiKG0MilaDenOGT5+r2DIU4MgafdoZajG
AGuAJdi1QJtHM2n3N+hnJzcsJO2y57R5QK89E068P/0WhGLe2H4agEbDWE4jmjHg/j+3vbKEfORm
/89VGvXJO4BZRr6nd1gw1VhM+tne3wusFEGWbRfCootsLrQ2xrPrfSlApmLfDNE7s+8YXHIRroEG
nHg0nahXwqjnBQNn/ZqbL6Qq4xb9ebSfLcotP3p0JublPPSv9kTAKqWA+2q7kqU7ErbNV9UxXIhB
gevBSdV9q6VFZfwDTLbAxlh7TgtWNsJaHaSlft5oDByA2RS5cRgJ0rSxYG8twGfdwP0vryzsKE+m
dg97ZNirpn30hql8NBGNKBMmtmKojLVrqufXO7HQDZ2VtcVBun+H9MI5R9h4Of6mNj7nX+G0cOB0
rKzo677AzNUbsmxxs7UzEPGHS0OhEA4j9nwFtist92XscHq2Ffn3i+NpDOD9TKUZEhxwCJLjmrTv
uZ7hawbY8Hg10rC/ZbW7NINyfliNPxGwzAKIWcfkD9GYlfDUoHZQw+WrPJVDsLlxPkjIaXw4BqnY
Mv8vucFlaEy1H14kVOmr41KjPUR/6y8yg016iqcS6gbo2+Vmf5jEmy4Mr/JPAaamUa8EJIEVIhsI
7JDEA1V4OfxWrYaFr+W7eHgJ8yyQuqMhVeJnmaAQEcLA1zltLjJeN6yUZaCJwNaVkFwpm+3RkzmK
xWqAAWI11f/CiAHmlV4Hp5eqzC89ijzsdUmmfndm7xDL7dyX+ihsbP/oj0IM2XAEkMAppodBvJYm
TRiIhr7kDlfBZxc5Z+6nNe7MV3e66DhgvREy60l9jw1SeBgIvtvHce2X364UH21GcuQ9rKjRTNF6
1GlQiHG9BLuGVYZFraU89IGh+PnFYW7vG7tOdT/nfieSA0T/OZ1Ua8Rr+GesV0i12SK0pPV0waVY
H39EKelN9tVanb5MOlVbPivLhIWLDC7rk33X+HguzZ7+s4YlulpnARPlCEjMjlz1UOZIVlmNLn4h
yDW0/dj5mgGIpT1rwo1BuIMu1/22qy9GUqoPuV8XLQuymZLAKt74pJF8Zm1dcq0CHUcpIsynpiBj
LNiq24zvntTfzxywaH7MMJ5LsQxB2PGPrFwK6sp8cExts+ilf3yqkeNr/48p+TRYWsT82ezfjwar
XNQXX1s3mVvwxSEUrrTkA4laEqB631z8atnPB73vks0Abb1MctjOo3Gf6y//Vcwh8OqczSzPPYaO
Xune32g/9d8lAGAvdm25/1+DBXejKcz6xwKjZuN0AHTsXlA9J06cPwfTynTA/qY+ronMbtW02hIn
7e5p+BaUf/hqMKz0YYBXdw7iANQ+d5/elAq81tAFIHEUleTKsXmE6WPwsnybckWaDC+ZCQMRFhT0
gZV1jLa2gczXgnv/vexM15Y7xqvvxRcCVnyIQBpjazklvJJlJ6PDHd55MWkleAo+EnJSoYd3lU56
p/8Lymw5hgdBypTjMRpHiAFBa7hQvJyVdzQu/RCQyC40SHes0LjDs49O1XK4oajJfYbO3A8OyJAv
vl7BVtehGFuBy43P2X/gTufmxUUTOJjDutQQdM9PVx+5m70eYBa6NpaXe/UqLIFd/qKfjJm64JHu
ZhWzAfjEwqQm3D3WQCLodkp1Hm5tpScxUgtTmK8GtV2/0Kyxqh25yF3Gn230wnM2cQ2k+pt2EL3P
ts9VsmAQeg7bpVY0nm1XmNJYniUkHJS/XPisKj4gSxLApScyByOA/61dM6XmkWD95JCguW0/7YNC
//IavafKfB17q1xPneqU/4wSYfsc2YCkHQnPa56NEddrx7abQDddH+/hTG013UzPwe+QbfL8V/18
1Jdua9F/la1+QI3Dy4pUqQOWERbpXy7kIn/ts6LkJFteNQoPGRVMCJxlnp6XO1mG17QMtw2RL7y9
fTGzJuF0/0u3v3FCQX6ga8/HyBYgzVbAIHM6+d5NKj/9zkKE2iMkWN0R/Xpz4OmyX3NpNKZl2FKM
6Ed4u4PxjMwCvLk20YV54MOcANvlnl/QUjKjq+4Q31xPtzm+n1agCaofvz60pd1qPDDmnXY2PjtF
opjOOuRxfNXoeIzFJyBq3I/dfsc7SxBWEUarZ4S33+FAGd+FQW5ka8THfxm1IHLOmtfiOzcbeR45
bAdFvaMNZFaEboL+a9xiam15zkD4B9qKtWURp1ja+NiVamlQTKHAZ10hm+yc58N15ucISn+420Xe
KGfkNqzgG7nqEJtpW4tdSiYf9eIX+WzKOOLFnuhp6mKZ0iAqyUb4GVRz+77NSqNvVDdBai5dGM6O
E53jFUcV/GNgHlu/sbuLSJF8gvnyEk3pVo3WbH8gqUbc/o6HSnt7v3Av/LJ5tBfy24oun69sR+lF
sSVBpfQqGedMfekL7v4DJd0Ec8WIxfUPKgdvEGVhCHrmWZQC4vIqTnTKoakIKKL9YJ72IBfxoorY
uLLgHOCbvgLRmPgDoM44nXJaC7LvExljUXFTjxEPZd7Tg2665YPepENQmpG/MI8Ck5pqVQfzrZgZ
bHpUTRMATkrGs6sYatWLFrv+0FL8B46MI33BFh16qzyBUb2S7Asq2m27d+Ga1nLNVKxEfH7ebzU4
wi98bfUID7ftQjSwUrRNh4pLY7m2fU3gvI8izPEVT/w7Jn2/YPBgYFEJHO8jgNDQJ/4sTuTggBHx
gr+WnyspoLbA1d+qQnu29skT/JZDg0PwE1AwWv2biYDChxky4S7BEsNnqcn6p9rldgKu6NDJ5TiC
ij9tTE9MzS/ZalSPxkvq9gPOILe4NfMh/fu/JU5m1aSY8kYA/B2k/HEBN6QmesHb1ZYduok6Nqwh
owtJmOMwdaDIkDcO5jx6ZLAgvwX76sHQCcYi+2P29RRpjn79CohO13Bu5rcLqZSqptbIvdYo7S6/
DmPvwz0BYMM9l29BaESfle2mxy5Am3Si/Q0jMilZy+h4WfxApJrVxOF4pS1xrPGYtT8l16RtmYzO
oujcVEShBzylNN9eAGQKt3Eayv7yORlIN/KgmxBdrV54N3PuBSK4G5fikKzGklZGcjkiFAF7yJwV
XEc3DzpCpYU2GO5XIZTFwGaTu5X/zMGshva6+UN+QtV2xkD8iDIBBJRfzLZa9ni7WBd+tBHqiE97
BIGD3NPp5G+NJG0fY/H5D+V1TjmGyAqtwryTA1R8yEJRRa09Wtea2TRwrEPbrDM5yAbgugEdz+xd
+hvMVa4pwGkhvyRAymesoKHcvBM06prC02HGARLw8H3Hnsj/MYzIqXT5GYloJO1OUn1H12PhUkNr
7ASOXoUUrbqfQS1Tg8oRYngMpIHdI0e6HAjS9OqQbhI4N2SBfBkVxymH1sFB8kfMfUp+PH6v+iq5
pfZ84WXUG3MuEUAvb0npDoCqS0Q9yXNSOSqcxYMDFhfTj7rZimGBYUKjKvwRRZ/q/hISThs/OVMm
XzlJrRa26AuMScuacQXa7ezOSiasGSvLubZbvKL8+LzAYVNYMWPaWGT1zFRrDAUhFTsotK9kbqsy
jDgZOktnR+xNxR3eRyhlygPs1CJCrQmqpd+kpr7KTgdKTYHqzsNfTgir8LpOkaVV2PUavqeVaHwZ
LrHyIvw9H+T/uqfY65FYJs8p1x6cgev4OPIaqnyjQBzk8oym1+bLhgiJKEGGoNpEASWLkJ0WeqpQ
b0oZkZZL7ojKP9R3q5glZ5EbF7xcFdmy85r9bySEMMF1xZFAYwvf6i1cK7nR9PNPubF5wp5w1aP+
KKI3EgfBUMbN7PGSkbCGoZdVoS5J0b6gDa9TDZOM9Cir+sV/z3hXdzNOWyr2sM0/h2/XENpYm8a4
qUnw6hKJMZEnF84j4bIPAbJ8/Lqvn4h2oIH2HGmpsesFLwV6bh3QtIx8ZiFOlSuLbFa6UqZc1fBn
+4P/tdaOuRlIayok/vHShfvFT9DT12AKZ/9Ry43q/yGxJDvyYXNZhd1epKZllBFHouB0dfTC0+LE
IWFMfLO9s1nbqaPAttQoDX1gz0nDpffi+O17PaysHpPYhyauO1Gb+1QivWgIsWKanNUTnZaNKzWw
JPEcOj/kdG157xoz0tK4/qbB1V2yw1VbyI1mnCa0cRQCiHQTsu/vcZ/f24wnsRY6/hbkiCBAXBsa
9s59EcL5XIMI2+Kp6Leqnbs2fmwoYpFvb2h0sBFCNzQvNwg6LpbcAsTWVpLPWEp3TISBmF3ckaDw
6JtDeTfvt0NipirYvIsCj3C9ez587NJEOPOq/dBq8MXWtjKFin3I4S++oC3h7/et0zIjal/Pbh1m
OLF8xRLQ+Byj+MTyGzwY+x//31T+NX5m/Xj5nCW1Yk/dF46TLAgk7lIH7V0KD3+vy0pT7eddEr4J
5Tvw11183HQeDUHtzmv5pkmDI5dKZtBe7eXWdWtGScKLeEzfw0TgFHXdVv6LockvqCW5ZqSa4ljL
mD39wBikAjWiWSHfBkrA96Bo17aeXO4fIR/+kjJZ+OHwD7G61QzgxrkND0nbNlrumIMGHCE/n9Ih
T1rgxvGyQKrxYNoBqS3Ey/2x8TEZSQFoVjscGa9jtHsUMPfoZ62WBEU8l+SGWK9mVngwbbNdVh5j
rAgEkJJYkETducGg9NYSnVWZdE6kGv0fCd0XHATfP5XAjCTqGJvtCizv9q8/FT+w0zW0lfk+ahBS
tzKBVEzXwmLTYyzd/dBqxi5t0kJWppBk4/X8jWPJQ/Juhs4VpWUHQ310Y3GQjl+ZlNKgmHKG0+y+
4hmppArGjtkBySOcCrTfDAwNWykamyzqfu/+DuVSHbhOXlJ2u4F+47l0tDsXGTpywEsRSgdaznbl
XX5nt3L3UsWvPE/Gb+zW1GMuuTd4IX1avfMTMCDyO2YAmkzEfcBmsOig70T6Sj0NEg0rPiZuTG/V
e5xSCDusCwJczFkB/NvLi9YbS7nv9qPu1fzUVh2d0TROfywWK9n/xiMH0zuElVjphwFupf4xJJvM
fNWFsDoiI6A/iG3jIC49Bp+NGoxyO+5lpdH76vR0bdx2LcNdNiB7Dvxrvt1CcTJs/98RNty7FMrG
yjdhrVPZx8MCh2W5j57McSe7rDVJ9Xs01mXrscYAGNCsmTXCTsJfAw2Er/jKd8NpqGFjJ9Xghdsn
kk5KOR82kVes7TTtrAJ1QYJXDPXuwaAlMCaTtcQTdnNNHR6/4s8TrI4NFhsEUHExWw33NXloRp7M
diGjtem+gQexIGPzCaPwPiUVxQfkNluH3lbknBPZYB0P4oI+XjOWsdPyu+zgxDPJQ2qSlQwui/x9
k0kt/Fp7XJsNa/C0mC/ArRRjlPLOvu2im8h0GWCMPx1bTJZH/4GggeTS34CF6idyL8cEp9LK8yiR
f2sjRSV00ElsTIk8yabruRjPP6sRS+jg5JUUpRqqL1JyngRG69YDehGuwSbiLgd18qgYbz5rllV+
DaoHd2Cqok9JGdw/4QhDX5Q7JXDidIg4IYY89rxV6NyZVqexTFyBP86Qgr0sP6Dea4XFgf6Pw/K/
YI/TuSbyPdQ+YQSvevYF236b8ziq1a0RdgEykIE6V2RMMxb9zehTZ8jg/i6yxsoZ9tRv4IVbFfN9
xYWg8qZCxAmsoJ3hHUbmWlx++MGnwQ8IxQU6Eq1eiJalHvUuAT41QgFsEtNjfQPMxrczRl4et6ew
QJ6NYYTGCBSVR+ufeMF3YQD0ZXDI3ndO5RknnkzMnnd5hUO9gDBLsXysvOmaFH7m8ij4UWuc9fq1
zqfYXicmvq69EoowWY1LD+ZR+5m8Fgzoajy9rQoiuuVW2DCVoILxk29D0rZXr9hyQ+cSK4J7aoDt
X511F1oPXIfx3NNuq2l2lL/eCvGwrWqgrCufV4CCIv4CFJyqCNQuVdoI9V4MA+dXms86rTpx+bqB
Tb/xtMTSIAxBAwSVlY5rpWQLzinK50Zm4KxBvL3zcks2+N4WQmb6KHiu1QoR/E3VMFtJ1PXKz1ti
Cx+RiPphEHp16VHN1sihHFmI+wu8CAr8HdIU5JbdRSPrK7hlDs/BNkUlkGlhYsRnjw9EcSnjwq2x
O7kbigaib0q/4+VBzZcx4sZrO6vGFDT3AbQZMa4h6C/e0KLwpRrhkXaUP2IjeFuc7qpNuyMYSJsV
VXW1jYsrieexsoqtIsv2fpNcCgkdZhYnCOl6IbdGha5RnejEkuIScVe0lbVnAg1RAeYZW7ATZJh8
LhocA4sQKZcYlgZNdVebOd9g/x+dcZveNgN/ewSWNzm7WiWVqQoHlbxCSDkiqvNThZst0oindgDo
vSCFB/acquIjh56N8bDwE8CBtQG82uJjrdM1f5NNYI2U0iTjeRG1aVxT2PfS8k3/B3m7Q+9HST42
QFOSKcnvub9zuh4Y4pOzdTjsGUheyPz/LogCJIkLB772krdN7S4Yzuoj9sFrR7jagWELvJF3MOrg
oqLL1lSr4/O5SHTgKFyXMs+zpJ7ovNDdfq9NYxW6fS8u/datCvf4x9ztU13wBpH82h4JX2PmIPnR
6xb7GJnxKfq/d7UpqNtXgYS+XlwNjh+wY/q5cF1pXel62krruY/2XagCJ0E1StiUa70+cXHp/Xl2
xGFkmJQ5B6EEH0i6FJbVVyQur7WJO+aRlQADGLWS8pLWIgLGrSsBtQ1rbqE8+vCfZ/hOY5xsZuQX
zxNd6jXKN9InVxq+umY3vr3XIhUhQoewu4OCnhfJun+8JT32kDRqBDgRLtsxMkdBYhEG8zc2tstR
Sd3G4VbyJE7c4XrSx+oKK2pBEpzmTwKT7o2UAbScG6es50CET0gin1lDy2oPqnc7co4AyjQ3I6tn
VXQLwVWcHJ3YGjpamCAs+FggiDphqhW8UaNPq40DQ7AGy+YasY2Ho2l5zwCGUUDMwVGVcNrNp0Zc
LOSmyxMYLxKswnAsraLv65GTn2S0jCqNdgwyQI0Og8ok0OzO1mTJu1TAAfmPfIDIh7F7SAswjynZ
kDyl6pJfn1Yaqe+D8GC6znS4u55A7aOhI5VFKu7B98EVA8hkpVGOk4YRmjfY2N6vzChEfpBhsKSE
SvQ2sDszu6r0F3qsmtGFJ0W34C92/I9NoDGDM0EMVhEzsh7YDyM9TA7SSrjmAmbKu+OwpX0mRGfe
sPTaH9y/XrYLDe8alBw9g7ghEf7lq1N0qcfCcWDwM6oPpRqP6yPi+UKGx9q4hz54x1VKJS8N5MnO
YibJ21WYyQW/RfN2SzozjO6CeP90gc4EHG8VOAEE+/bF2OGaIBbk14Gx4t3IvXeWIRaoTlmbEbsU
jyaS9upomRut92UQkv5uPr+kUYsvjAOdGUMD1AGd+cVjnoZdjQZm6LxmbEXhrVl13JS5Ykassvmv
MvYXghMQOufp+5YRI3kUtDGlZWXObiELyWvNzbKMkWfoDebM60fVQzRbwaR5gs7NL18wiWWhtVNd
ApR+hYelM91Lrj+ySCCHxSZ+AsmGHmGNmGrZgSpx26hcwJeKbGXMuyENm0MEHE3VO+8iU5xGP7ec
oPiY2Sdd9Ja4qeQjS2paHm7wXdFHXzKzKJF/QsUg+W8x9iMn5t2L4Fhcdl0uyP97QiGSfQgE+j+Y
Rt0h1clqdrjSgbsrZBg9YXFDR+YaB6HggMmyLrhDNM6WTo2CAhHFaqXTomvVppQgZoUUZCL2JbSs
Grp9BMrtCw+ZvMcswsYhzVibA3wse2qdNhtaHie0lmjHkzBxTV9gEnjHjezZqLkpJQvv1iKOrKeA
Xr0rFIl1waz5OGdmijw/WwWmH6PW+LxXsXa8iB5QBsix9XHKbBqM+DGKvyKth6w21ZktKHKa4bHX
BB5+t8fHBxobCKuLIphYzUfKDDo/Y9UR+tuoLBCoLXrZD1qYOf8ID4nJQUNMHzrdB2n445c9w4ym
j1Uvn8cqxHrCB46NXA4kS4kSOmnyqRJGJAuinTEF5K2Q+VnDO5c9u5WEr5HTY/V/dY/vnoAkrXTy
HesY6a2xBRjel5FFAnRpMrOxhT9chqYRs4AquVZTRl3hay/ezSTqregA4QHhbNUWyVI6JNzGfsUL
45JflLnf4pNKRxIE1TQqaDFfJDp+5PO2KIM5lZYiVTqownwRzaEouiJvuHtsJDFUXVivdfqtMAGV
u8QYk1yHZTm0xq1KR4z2rZFaSl03ADo4j++AVTlf2E7Ag7M3K/PjgNd8wLqe8KFAZAkalZ42bnhG
GuZy8tsokRjf1wN001HER46RSr/aRuss41Ii1V68e8h/Alt3yQo39iS8TQoaoH110F0O7UhrNeCa
Wp1f4XU6Njj1sixF/PKJ3DSVOHglWZTT4eMQcMJ82qVByj+0ID5Qir7VuCnXHJneqiqOtz7ypoGL
yotK9rGThIDQ/J3p1FQ9QufbQIGYCbY+1E4tHKnYZlFwVuSekjTgalwGewJpR96tfUIADAnYF3sN
HR8UCZlOnZdTQfU3WL7MXr4HHKXrBnVibW07SD0Gt2YSVYxkbyacHl1MdaT2kt92jYBdDTdD5sxa
PPn4a4R5ocqcpqn5ARP8ld/NSQwZ3uHfJNWh7BSSyirJ05XfI8O+ifRsC3C1vhJ5MxJqnduk3lOT
tLrV8/LSlowekynEFe9z5h2DFmJ5ZFSecVP/QIPRji0A6InXK/65gvfdta7NnKg0MMIfCTDjDkzi
lxYqXmJ4TTTLXSafSw0tb86Ww16o61SANUZTKdxN0wj5jRKXYvxe2oCx1aqvjeja2TK8tb/Z/URA
u4a1miIx1xWp/QJMgbDhlzhq1M9lLFk+hYm9mnxXz8QAAa7ApvHPNeHZpYtZcazBNsTpD14KVbwa
kyp5Tab4stGg3htyKVLThdXIVSE1p1lBSDGXNUtjR3JNKdr+61EU8Zht76i17GjVXY4NRaCctGJ6
qfSXVSVuprhaebjKWFF0TcXzS/Nn84cKf5kQ4vUplR3OpVOe9IaQv73YDub5zo6xzVF+6uIxSYKs
Cz6v36szeDs0MpD7t5LEgA9ooe5OymmZsA1Ng4UfF/xydi6IqFHuZhJVEodZmZyDbOZ8dK1phqVd
Axk6XLaQeEk+YBLJWkrRg2jtHlmYfHq/EnH5GxprtUGMR9IwaAkEQEoQsxo8xXiEWrtwBTXqjcgX
lgzNdNZmBOVX3wh9GDPgFP8IqfjPq7OePImNJjIqiy3+PLjRCvKWEMXaVIed1fNSb4Mz8HmcALMo
Yg1o/itS0D3qpUd9bC62EqJxs5ziu0BVnv8W+bZXJhdT/YlDykJm9LvSLdZxf7Z1wDFw/57ORMbb
VAaodxxrX85Krwn8WOLfCLKDdlS3y3hp/7gHLczf681KwMfpcGWcsv9HRCy4JG3Tyzu9ipJXzBup
ST+uaKDYZnS82+8RjqquewL3xoexDw09xtgLOOdj3jTniUqs4m2T7uT8K7BfzPoszjE+SUFi6RVo
K/EpIMSyKa70ELoJnXIcINDRyqtM33HX+zbeAA5SXBAkheaNX2LFPDsOiueaHA+JcIO9Y9tm3fbG
+gLqmAv4zbXPPD8BT5SihwtFU9Xd0+b2Dl5A8hYlde8TJ0TmoLR9YQRlTOJ42t01/GMU4GexXrZP
blGt9taQ5YTWv72kUPmm/4K1TihJTkTm0mj1xf7UmeNjRDFvSyIdHPyVmcc6j32Q+PFENjQB/z9+
RpzAziKDCo/rmO5aeUhk1RoMdOt24MyF52rsAvy05EWDTO2ILEu+Bg69R2TXqRd24/FJGOEoUwuW
Qda0kJyPINLVtjTHKE5hySCg57N8Z5Feg/KEcAbA4/ITkiUN99p/+X2adP6a9FbLDh2bxj+LsG3g
q2gcrF+4+7PporzhhDJLTueLwqIApS2fvAZZ2QaXiVocHKlJVCBcPWBNL8DfuCLV6+1UZvAb+R/K
mv93qAuJgjbtQ4ONlKtFrMMtdYqezIlT7cjTiD0wG3VXiJpDb2A6Vdeq+nfw1QDaE11Y3Ydd2+hk
3JeCQ4G70pMNx+q4NXDkaKFW+WaQ2rBfCaa/HzxoPtNcn7HF8w/Ki5rY65D6TLItTbqCcbUFIPfz
0GjJlXYdBTUXIiwUL2NpmQZCPACaQeV2ke3azaNeYY9bGEfuCgcjH787dX44/pTCSeZfAvcBSyZ+
oEmrMNzKtAVAL1z0xs7/nMblPmZ3q2E6eNDUo3iOc0sn811LTM2Jjz/CMIaJkJNYC+HSvEpkeHVI
b7WFbzfJR1ifW35gyJ1wkgTrUnXIYWxDBmSNy6NXLD3gwSezBuPpIrulM47Xl0Yc84nLTgpVD810
EP2uN4Dw3RLkwet2CGXxcl9e3oKk2sui9/GOBbPL1tvaaadg/z9pImGkskDyFZBmiuki81D0Ccnb
mYkQFYkM6LnVy/bn4kqSE3k6VMjr5kKyKnHHKS3rBgRlhBvZq7eqBqFLoZ70U6ekrUSetjWB/Z4d
xJFO1gy4dd0JbXWGwDyrvactfOLwWNZBaEiyeI1T402TT96vfNCubtbOclv0s99qAboRDXtz8kC3
73yrrS+fHymsXtRWcudsjpW/RKrvczD/FzRz/hN1SFKHWstKBDkmO3q8k0lrDxDKkyGnGO3zPpCk
rIT6kuUNNWRQIX7/JC8T0NlHSB//GrPIwoKEiH5TdqInF1CSB3pl+ZKhbTjmyFHssMyCsNfNar0I
jOvXnVLMudyCtTDuICTrWJkNWapGUqYMDeDaIba9qiac6srUUfW5swXQeJkiR7hmw2w8IhE1xsl2
hVn5yNOZ6cbML30q7WvZq6dqv4FPRM+3LcFglrR2Mxku/ugteebhjmG0PWhawFGCilFDzTzK8W5Y
YswiXTG9Jk51t3RcYAQwEPCQ3xSkmuL3Bcen/b+RRduem0VHzh+iZCdPnSTi4gGHklncAhTCWYtf
o5g7qs7Ogllw8CXeMC7DNQx1KKhB2P507EaPrRkeZcjJDHQKT2TiMMJqUdi6taPOQGp/V410EDUt
LH9j0JWPSKZsknqxOvUT6TO7hoiauqOyR/GhU0SFB0Ox/Bo/A8AQWwtnmaxglFvuRlNi0YrbG0df
lbnoEy6oM7EoIPjiv4N3qFmamY/1QPNtbYiOqkGAwBa+ZVYZ0wqqWELczhS6Je2AhIw6c0mNXsHK
mMIVULDjFQmEF5HrvNJ5ogCMaICy75hKomDY6lTKwFGg9FximYTEZGvx7QRq05RZqQT+aLM8A2fC
z+v606k0uqtsba2kPeCnDw8Rq6Fl8Tod27X4DPigI1gy/p8bnATgniUM8PTp0bXkLimomB6JFIOm
YjXa5u2XSTYDYAv2DotTh7z5kchtL6EGnL2mNe5h2dZf88QYND0+1qVeTQOQkoTIRk9BWQ6SQ4W0
3DoZURGWiYkMWH+lyj4Z9II/nfwRkwBPZs2wSzRWEe93hhY5xFzHMVqWZ1W1IbOzDZcpGd2Ui3NB
hhF1WjK+8c6EnR6sw8CXwLgnkxy+Eg0rxOLoCBrS2HINg792C5647ZBdyYgk/Z1I9IDCowtGBv1r
K6auPHKCMzp7ZJnuDMuVt2DJJM6lYLHknw2L8kB2h7scJLsO0R+SgbKpW9Jgox9S2X8fbFe+vNFN
eUfSh9xllop3HXvMxPp8KrlKiU7rjA6c7cBex9EpVVw9adMqnrshwP+ig/lvMDQCM3fimohdHLyK
r5IuNKBOs4sEwTAnv8ZqvhAl385gTo6yPGAt1GDe0aJiWY61Q44uszeIJlFAFOtfg0cNAK9ooaCJ
vckVD6BfOhAQDx0hy5eWDeN8ZKwWYk1jWPD1b8dmrciOSwg8s6Flpj8m7GY4w1mYoQDZtF0GSmiu
ndzSFzTM5Obr69iF0ujqdfzSB2EK5Yu5o4mDot24R061i+DGYqHrD3oaIydIu52XUi4vpcIBhSvn
0nqDutyp4fQ39IBwX+AubWcwjBlSIJA9sMjn4/w8cIcD+MMc0Rn/NL5KKwaffG7ydPduUk9wPZG0
Oqy3edi+zxshI/cEqRXd/6IZlGMNKaic5qyLIJlilUi9xwLrmvgDKwKtR/1Ne3J0Z23HGkEdC3xQ
quhq+WciaZVq4vWFZ5H5Vc8cZkthRXVNyQwdC7hRH06rtrojRzVHLreFSqQi/wWeR4aLQ5lKjE91
LhSP8fK7yf4OutaP5tCRN7crx4Ai8nA9lbWBbBQAY3HqP+ReJB0zwvM++CdwQe/JPIyCVRe3b13Y
+waZDRO2oNi7NAdy7osa5iqp4ZEoTf761Xq9/YKElWhmFpiBaKEH1slwbjApMB6BpMxNkJZoyD9g
o5eqYCKrfOcyRJ8ZbZAcsZWkc6RS1jMsKOcD9YWzZ71A8D4JCF/KEezT1jVJIz41O3Pyz/QMuWSK
aUaHak3eNUuzjUiBRyrLoMnNWgleBJa9/b6Mipt0wMNfaWG3IUEC0sPZQoV8nsQfk5lUebEfpT7c
73jQyXK/AgTtZr4f7Zizz2NHS7Tgs2s8MOd0pXDrs6EAQJsJULKhMMFgaawc5wRWQnfdS1Kq9vgS
dNzW6spzpmCTMoo2gSMNUfPhPIPHSKSK5mz9kA/Nn2BIYKX8mycxJpocmeK3c5Jn0T8mjUkIXgKi
0iGjfA3ZoplwUUaGipfpDPwd9EauUE/VZI/BEGPZApP3jj/F75jJy3CQeeFC6q6oL+8gjXfsnrAU
NYVADvA0xYEzKSOdVE/fqk8r/vlj3tjJgVvwBL567vzmmhQ1EsCBZlsI8o1MFc5e1P1j8qmdAw3S
iwvTLqRKRp8ayVMBBBAbW4SkkFQnbTc0zXcbOu0AihHHDCg8AqoODCH1JR6HpwEnoQ5tgJePfVJd
X2hAKKwIrf2mNNuF+Pf4hMX6FFiZfosUAVhjKdL3D9YclVbsNZVYGWMiplr4mPOt3FCrv098UPz+
7vMMgjEzEUVkvtTTKzt+O7Cwp+RFbub5pGdHAamYcCvSKUvGObICUjrOHqLunY951VAimfk+oun2
8JYWIbqtldd8/Wibdd5XPIDtKNtbpaul0DIdx7v3mm7b9BpMm9q7+u3Tb0q4fvdWj/I89E3iLg30
BuSw+rnthSaAs+mE1olSTi3ONrWo6RsoDrYFDSmlyc64u0kySSwsleMqSt86jHIKjDmqhowIBKJ5
qMuGleBUtW7BLf5VStX/5Lk40m7bFS3n0Z1fTqlbosDqJ/9l6S5CBwPN4BNotSWukihjQI13FtMG
FdveRnM/hjeUiUbJi2RXLfjl3gAPgCfL9Si8+oSRST80dz8/lX42kdlJIOeoBOvbCq5EQp3NHbnW
7jPc6RkdbPVGThLauwk/AU72XpmyflokhJHHE6VixXwoo1JOCI+VV1VTAH/gkKirtmAwe0yX40AZ
sQ16MNa/uxwF5RiIdnjR7VbCNe62/137xwhzqTsDo5JzCloWu1WLfhY4vdlSAlAAANTR8PrMo/Yj
6NYJ09yFFB7wxNWL74cGHBRRukSyGmpoD6D5zRlQ0xor/2T7LTYFsAKjhFdxaR0od1FQ2hvNiC/H
LPRHBki1uVIj2fwu9gfSrEce1AbRroZiyGYCBCkBkhZUEtMMI25LXlGonEvrAH5XeClPcVcEPZWe
RMwzKGlCDzvAuX6g+32E16S+ezHnbHNeiW5uQe2Hw1BGPjUjEBPW+JdYmSSNK0/Lc2FnX0puAWZC
VT6IicMhwbAzGRa/alq/UKPulK+QqagN9VSGkX7jjh8FOdEpozxXI4urJGiGqUlvHSYcvwSDgYQn
gVt0EDOSkXSUz8+xacUye/dnjwn0ZDGgpXpvTnbFsptbavtaMCwwMv1tVsjLdyTiFfO3L6gPCfI1
jDRt7cJh9p2UM/Ge3NemaLZ8IRVpnBYN9tnUOTQwfTSdlpy8m3OQN65flX29kG4opPzzcX80Q0tN
xw9y2/u49C2L+WDRT883gNfNPOzKzufdRTcVg5iaQ74acRhoRG6PB3Ec+uuI7k2Q+ermxlKYGBaA
eSI/TrzlhwHrFtMx2EoWXpMWSV7AHSDF4FwCPz32SVHB2OZhEZAH3eetjOGMs5FFyG0j0y0PrCfb
UpsPF2tSXsMJoVmKrrh/ZSv4sHwwb1nku0NPELs1RMluEf09FJ5MtpiP6dBlvqah/jFwLTZeisOC
bsdU4sBRfX6UZupwp0O3wNBBZodEPNAI+v/D/pNC7fU+4Zm1n/WIRSJ6RF7oxE8V/V+ianDollQB
wEdPQSj256AbVsYfN3mZ9zwViJyjTXVq9DvrUel1nT8mBRcqEIBkLOffVS7zsWE7G5bJg1Innj5+
EUUDX7ot9E/mAIfgcoD+nH5VHish3ljGhLP+RBZkO9rJtOSRGZpg2uI3QSU8cxB9k/cdF9umtcZd
9YOo6GQvbukMtf095ZVx2K3X9o+GZG5sn/UvNiu2KgCAcCTWGpSfZgsoJZH3uXbasrUS+hxUFElD
D2i/dysPVhTOdbkTEwn2olMwXM6gLTp5ovVrATBi0/EVPTHvtGjHj6LvZEXjwxJNdM3UBtAtwDWG
ZlvSmYYoalGoXGVXuZKMSa3Q05bsWa9u+IbzMjaUfY61znLj8ydZIhOTWHjskP8YVLJfkbfWvGrG
7BOLvuq7ZQcvVibPF+D//2HXPIDMKWFlnAft/1jBBKC1SrC4tcyBytcPPKqPsbWxplW6aIm9gLbr
oYxM74jDlD6dhAL7sw8SSnCYQNpvZ+pbAFI8ATHZAmBl+w3pQ3kyXb98NqYUzVkbGsLKo7EKtVX4
eua8jVY876favrW3TuSm0ET36DMvVpTa8SuEYrsLeQMoUcBBGgqHNwQZKA+9/Tj63dXv/dc+KiJ+
RdeYj3nZ9jAzD3Q7c6El9ZvofKfIUMPmM5EnPcd4s3JPp0rltfPghzfBovlBYaTHkjKN5O7lSG8l
C0mf1XnokBZa/Sk0OlQz35b+AWfoy/UuHyEmu+WVLar2Ub8NuoLYMyS0VAEyJncYCleP2JVs4INB
8mktVgxU1cSGuOTC9qfOPhlSrKlNBnaTS+EJ0JiLB1nhZicvafwxOaYEyiYaea+4FjrAYUY9E9c6
LXxbiiPoBhIvHVsKMWL6PkSO6Lv/1vo86djaBdMOclZAD/5xDttecw7EmkDNr3yzNKE85RfXNB98
sqA+lBJHqSlGk1I09s+6q94tVrSjoQmRzVmATIJmeXbroZY5H7dMSIf2jTLv+/fvIgtPf4632jGv
LqTHCmrdz6h0EenNoIsPt7TRznt/zmivtG567lVT0atOwXWHnja4uf/PgFHp0l+tuL4kkhG4BXNT
WH5AExb7IjhCLTdKmmq5gVtCXU9FEtPA9BFjOCCQQzcwNirSSxqzq2hyAq7VZS6EgHEMEe7/ukdn
iW6yDtHA58M700BGBL1dFsLaETep9ew1ojhSgevdJcuq26lHlwfpaP2rndt6t1jhEJ49QJf9dsG+
qkU4qflARmBJ3GG9+lq1jfqceJHRQ1iawspmLe16XxG07AdefHD9T9KbE81EFEBOAZCFnNWEYM8S
jJTDUNpSg3xdTa9wrjwpwbWC07uy8qYjAiHEfY889PpefQbrkNMGpjHVOVehFqQslGu867SbW9nU
guQIyxxoNcvsI4yF4s/q87qY4TpSUXyb3ippwSN/TZS13p8/Tb50SNDDiVrXc6DyYpeIsvUqYB9J
2FL0m3gtxj3/Bh9yRdUPgqM6ETd4tChwX7UWRZNp0QW/NHxXYBgdmz6FCKhe36mXL/2tiA93cxV7
VMrQMyKF1HPrNxbi7Gj4cUbD4xYa7Fz93vyF/cMDBfpBD/IrpdqzJjDeBoEEA+UnJyoiTgVxxvoN
V6K6fQInAN5pcjJkQ7lWIxciPHrCZFpFpDvKahVjmEViDrrO+Ph8t/BPA7QF5XNM/mbMXKtb9H39
mtOzrxPVc6aDLVxERAd5zVeSWnWUvcv0X+xHKkzCjeM9Z+lJ9M9oomHjQCXiVi3suLbOCO79Hidb
j/BiByYBnWVYFnB5onJU9Zd0ishTldakk3cCQ2s5hGa3FUsyQ717ROdEnEvRqZxF+dRNyYIkSE6I
cNGN90cp3cSht4BKF7Bs9Wxk0iaHM5QH5B7pHaM+ktnhWTDCcjb0hhvL8Gjgqqs0AgBo+tZckfnb
DFeQiiW65WccC6WcXhIrykMDdjsRFtIF00I3spjA/1EmbuZYZIvhmOvaJ1JJdAuD+7x2v+SHgWXQ
r7B5t38Hgp/AtL/8LC06UAt+Zkr3ZG621Uy+fPeTMSJ1pqN5s5jpc/c4psjfVQy5xlc2svfg0ah3
XN9FcN6uR1vFMKuT9sa4g0tdrPAyZgmQDX9H3ViCS/xRMs+NYTZF5uOzqsCaeYQ47Zxl2TWJn+/Y
JWiY0axarQIZQT9R+KemdCqrOjXnADCgpj2aDMLVn6h/96Xoow4d8BdptRxMzsekRYatmZpKVjG9
QQAFEkqryIRrOLmm38nloW3vwLCOfxstxD05M548Ayd4y3ZfDC6FI7BN6RJGHrSQ6w4ij/74je1d
mNWMiA3/Au455ClOJGmakVLmjLfYc4Ir2MrbIWkGJ9zAHHsqmcC0BOb462gisznyLdxu5kbZEOJw
HNOt7292/LsHenZhXHSs5b6REsroPjLlH242UROe3OOx8BNa23tAhQxGhd85h9di8Mz6v377iU01
T7oioX/GFwe4rkUsN05nB/UrMKV6zSDCxqDF8JVip3XTS2+2/pHNLU75guoue5jjhcAcTrUnmCXr
9xydqML5HI7ZIO/7CJIGZd76h0lPhbGugmPqowopps2E+gxLXqmP9TF0gKsKDzygpjvL4UzN2wL7
SbWV4h3Bks/pOmHQWuvNGiOFINoXOlxJBuuySKZoX5AKFXti8O4Bfb02+uvGA12H4ELnZ0noWesi
i9LGjPxWrZOtbNmDfv7K07p0x1fDvs7PbEAj5aNhp3+vaNDNPZMt4v8I7wYr/q0D3AocKRP3E29N
0DVihJF5pRhcNCxT5iId2KgSyCS3JdllFIzkp7OXJerwEynNPFylQ8ydVW9rsT6/mKugVY2+dIvS
A59qOqrVx3oly2AvZz0wcAzspXirhigYtQ0xjBX9WUOHN0xDCHH+lNvx1epnOSRDKVfPaLwlfw2A
Rl56Pcj5jkpCDcG8N+jD6Ucw2Ce7szlyYSFXrYehrDjLJCN+odXIjF+LMvBxt8a+++B3BKOyQVey
XfAdbPNy
`protect end_protected
