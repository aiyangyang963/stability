-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rdTKiSC9m1h06+yzUBThQ58VAED3cU+IZlM0wbIVcwkfuulrrl2vU87bDjhaMRImaoMaF2rj974d
E2HQAF+C62Z7yaPucSglOB0QdVd0dvZZ+Q70Fn7Vp6lyCNdPFCv38airTqfgx3SZU9LKnttfVWk6
COsVsVqHxtYG6qy42XwuFe7GtFFLDuA8RFzehiMoS/7HTT4YVr4l3b1JCsYJTEBnz572/7kZDt/7
bp4BtLGHJR4WoLOEGPAtCAGG6WbRvynBkwg29M4AopjR/ARy1x/AYWnH8WvEd7VU22ktZO0RurDN
Ir4DvjeOCMMraNfc0Op5BLCnCDCmhBtTls7KOA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
f643E4OLv/3Q5sZR6RTTsA6z5LTMjZjHDGPkmVvHRmhYzGe1kYewM7kQ94WgCEHJbf2vKOtoDisA
WPvz5GJiBbjYCnKkoofct0dj1XJyC5W7n3OkzbjMybKSnBe5Fcoa2zXmGwX51UIqrbbNp0KKUVRq
Av0ucXXSRLlRuN4K1evQP/rflKSwgLIazAeCYIMH6xuJ14lgQY6yFQa52skhgmevtNNeIWPROE6I
P24/o+BwQhfMDBcaedku9jbELD7/NO/LbVTKFmieih3UJw7LJaXDk76ruBrMPzjOIiMR7XlyHryw
cKfeyxzC1/m9yfO4J5ionqudrRvfyZYps4xjWbuh/tSlweIAwA2hrcE2tXJxhRHtYnRS5VLCAny7
ClIJv9WA25Y5Go5d++5nx0VAASqq1YnTT+jgI2mV6d/YorqDqElPzRG9DhDhPBU17vsZYGZaWxNl
XLAHRh3iAZYw33pB7DxXTLJuU/jFjLTDxBpLGKUeiGY+WkwyjApYaE9tGQwbszzGiFdRvABTgp29
9TQGSS7dKv2p39Cdtz97n5J6fljATaAXofqu+MR/1SAockqEj2hBGivBzIpxa9astbyInde7jcq0
StY4pt+qp0vrf/MNYeGtMLwyE/O3cYXN6O/HmL2T4kBCIFzfBIMX4cwQNwJ1bJRfbdbakTimBeuL
DLcxqXlJhyNq/D6/v4A0Tx/OjKRg2f995EP5i/r4v8ww+ZqAUbcOkb7bYe9FT/wvoq1gxahND4g1
UShXORBiQyUTB4epNEaKtw70eUDLvC75c04cil1IkYTkFlKTeeQ4SjE9ozpOM6eUD6B9cAV2kyym
G30g9HCTm3Le6aFZrlPE6ac6Ovn5ZJfQyFbD3X2TcdjLvI4B6zlHdT4ggEEk/aKZ6RnndWZZQCZ6
bjwXMCzEikpb8mURgsd3az0u9YuEbjx3Xyqoya8L/dkQeNHsFQM7LxXznQ7WjN/Y+pvWennfPm/O
ovsEinkjH0XcReTrSNbpT3Kk1iTnmbkOswKWu9BZwuLAgktqhrFmFHMO00zuQzZiqjXz5Sj3NEAG
06yMX9x8Bzrn5WcLmRX7Btf944men7kCQL8Gwpm37jcN7GGWCjsOwOq/ZFIQHvwrdfV1HxU7Y227
JaVrbroVKvEYvIi/Pf/xmKmGoNQsm/doF7QA7gqAbZBJqjsiLxMFdbXPcbtISBLdf4yCbEmtZqGo
+OgvUnroV4oMbykkFYP6m2N9O4d8ORsraVCKhux+Q901HHzmQoFaCN1euo811Hjg/09w9RfryieG
7+YMIY88vGFWJOA8iv/p5AbksnPqr+Dd2HZ8gY3/e9YOvbmwzheJdMXc61Tmth8uaDMeOLd+x5wb
cU/9CWrnP0ISRWd2kIlbYpUvUSn7CAGkS0bJ3lVZCo2C+AUPsaIQHvIpzp5BQPVFavX/XxqO6PcD
yRyw4KFRIb7qWHu43bgcd2BkqDA9xOf9JLm6RAZ2cG9WiSpHLPu1cKXBlDx2sweotqrLN0UlXmvB
Fc6L9JXQY9PL1zX1b89YNGuVRVcDRXwQSdKpJjSQr+DrG+q2j5olL8t7XArFSV0rCTy0Q0Ncq3yk
f/SHRAWk5T+2I74hqV6GQFDXpRQb6iiowuV87BTZLOty1ZpyOQdRMP1X/pikw0Z/yO6iiTME1U2D
SlZc3r34fqdkpV11JB6Ws8gqsFYPNv0oUsFFA3TI5ss9oqOegMgZhimnKtxk9+o0LAdJBZQRa3tQ
kUUhrV9P0l06UTA9C5TxKYbKUYIwHKVR/IBR4CmW5t7ZPv1v8+4Pw5T+rO8drKHg0/C0aQZ5hqXT
SJgB1tRd1G2XfeSla3Rm0SBFIFrpCGOX67XOUMRc0OV0Y0yWTpHDV70WhQkiCvYdo2fGdbdlFxUI
wacqqWb7arYPl8wAWVu83V+yeQ5AJOuMbuXfoEnbNnmDujhLxw4IFimXnUOOci++9ix7+hmynv0U
q+JJJOka0VYKzyZgBwM0nj5exhZscFodywDGD8XGrLR+XJgc+Dtvwvi+O544SJb9iIV/h/RGa5fj
h8lgXSCQ4KYRNaUnqPfjeK+/cH23InesNHGqtwLsj6ld3b780/nDAGkM9XhWP0d5sj+3E4ybTDtw
zKzF0pbIh948bHyeEcYIaO+OJSy4cXxI3eF1EHogo4/jtnRJlfMniaecC8QZoNMRV/4OcKfsSXVl
tuxPYI79EL3DbLqABsUCPmmLUr0zdOIjnfiIhilRHH4xz0TpnnyVSfVRRNhRyPuImrmwHtTLyLpH
kplRPKcvHpD6BGrq7bd1UPlh5jLIQ23Ze91wpzTCoO/NDAoEOKK6kV5qJEZQRdqr5ibiMzPv3W60
6OBtUccuOUhLnWAxHMaxjvHHUTy6nkRDddqYn+P+mtLAfS/OuTIf7SINllsVLZ1AoKLHLloMYt0v
2LwsnG4u2AF/74ELg0CDsbCDLKjRqEm+aZ6LdNW3ZYj9dY5T0i1nUZ/KqkLzV9TJdidhHd6amCIF
Uek7DXm8BgKXbCrFZQdlYK76h0V8XodmoodJLZLBAb28mYuIU5F5CaLPY7TRLQksCpL6nQ6HpgzQ
vA/F92zvRDw8jFS3fig0X/VpAcYG0Gn2HfJsCtWWkiWTO9h9K0wTB1JF9vF5bhqzC4x4O1lA/6L7
hBd7JQ8bVpkWeenPQN7uUGm8tkZTQ13rYwSpYW2+x9tJ2aLpfwH6JZ2+B3jodRVQ8fNuig25t/v3
3jExxHZ2KagS9cDfyqov/TElCdCJ3ekVKySLA7aWaNQNr1VD3JGiMQpzhXxXDDJ32c6ari1J4bbd
se4oiAx2mTqXn9s+H3o+X8kNzk4tKVrmxtP6KOnWKL5zkOMttm6HRArDTNg+2QrawyorSQ1C5C2w
A1OtmNtpU9oZI3VSV4iAOJODztZ+HgnS3+iIiGiVuGxhApRmBBewDyQlX2zcYAhxn+3AZeKHq8h0
CmZ0k4C/yLp6ZUniNgFchs6wqUhTCSETjkgX3iFfGY8z2DV4NQfceD19LbPr7zCsvEDhpcaF3yl7
4/idB66cy8mqo511Fe9HuFwJYBLYwtVW3IKSyZOpdcdvuDgL66AlLplNvltnEAhKxf6eloKTrQoz
ncvg8W9XdUL+44btKkmw0jj1BDGUCD7mKxqpm9WzWI8NcLlIk7VP/+QuOZu8t7pwZ0JJk0kYCAGj
e/y34cjijgJ9TpQgwQt2iMzVxEWPgHeQTHdgyGL3UbtJw7nDiD2WBRajdl1CnNpXYi9xx1siv4kg
xz50YqvgEPbzv2mB5CTgkVIxLYmHTGTUg6mGT8DA9G8syPyM94G8QWQbhZLmeMCx8c/U/10OGefK
Ws0caeKy5TSDTKYzW4uZUb1OMXkwaz08/+oGEGu4P9LaCxU0CmFfN0eKub/pV8OmDpeFdfWxIBGc
pDSYekJHK0JJFOGciFrp+GBnBwW/RKwp5eLQ/nA5PPUm8yZvggE/tPng8q/uhv5oR1IR7ptFGiFJ
Jad4j5pv1S1BqKWop66IXBB4YDME+BpQ50vasc87P9TQDrkMfGZdDubvJpZ0sf7BhNG2dEOIRDQW
M6SKieeZoqhKOsFdJQo9bfmxevU+XcmabhzT4AKTVBLdGwtgjXZUPYPIgzG4hRI5MA29adXaOBTW
8Yanti1ySBdKnYxJ7lnu4N2k4deNa/gomyoDf6ZQf3agrH+B/G1bZpi1R891mCxSLUgf9I56z5RR
ZDIhGolI5RtCFH6rvQGwe4ZEOEKsJyNOunz9xOZqx4VtB64cDPBAEmcdWuJopExJei9teBGlGKdf
7mNlg42ZgnUclp656yXMNl1DE4Zoaj7h32qIwh5doALyigIncojTgEPt0fZP7uZGxKWOILqiB5R5
JxlSAm/+UfbpHDFz7oJVEgJRfrDuYK1a88EVZwkNEW0FqcCJ2jGZ/fReiOb2AWag/JPa2KiQaokU
T5AfYoL3yBwHUuaXGYBXeCgXk4AgPxTpbbYqoOiXoiYSKaWBn+p1FqJVxuCSjYfqJP/M5eHOspXW
m4NAz56+tA4sr0SvGDtkUjx+gqJfREVMomwWngfrUig5Nfil/Bknz7d1WwhhtMzBfLpzdPcFZdkP
uWEk/Yv+zBtYTvMdF/WyXmR4IX3Hh8i+3bWNcsMpoMnPJVINg3HRQYtBdszK6XPd0Re7iY71cUSE
+qyoYhKhDxGfCzUwgkM/3n3OWyIPM+FP4THORvNPTEmvTSUv9nys5DMkOaFGV10HFfjDu7pjBTTP
TGnNN2evpnFSNahQVXgNz/oxy6ld96hS71SxIoYrwsKVDg7y5P2YSD0HRx4GbR1zJTedkKfmn2N+
05DUjFUhwiNpKf1NFa+ON3nT1oBSunKH/D8NMuM2kmKW3IHUKCu13QQ8/AiodB9tcI/yYD8AF/d1
RHDyYwNJegujJ6s62yqT66kzrYfpzDRIy25VlXBzQDZt02bQGERUnBX24/QRt0BS5WFdwgNuLnJl
ybCOrJYP4J1TQIjQcU6jrWNIVROpA9NlOrUdRfuuz05L4lgkYj3v/q6pd8ESUdg5KMRU0hQx5si3
VSuxIgjdu+83oARCRYmS7ZTWLGMBD2jgXXA3uBYC/WlMeEdUKRO+YX+btKryPRgb/D6pjRuXiLLb
VTexc5JJHY2TX1RpUr58iK4aYvB8ffzAjRlkQxBCmLQdoMQfM+kGx0glOzE6gGt9VUZFM1uMEmbJ
kD3eZ8z4VAqbZLXZ+1ZZHzp7w8CioKGh+d2kghlCCjsCfY04NdKqadrPgJS266o52ZkaY2Vfc9Vd
NTO1mla7G0bJbzUAsnFu6GxFWazQ1pY9vMC9g6869v2PQEnE74mApp9+ZrGk1wK4TRcn8y+O1zuh
q+9F1hTcIwVbUx/U3XCMxz8pIYofQoIumtQKaelc1f+8wHYJKE/kUkgF4El+HdCl17fQLvmZWYO1
AezgEKdygpqaIseQkQdn3YcWtjv52BHrE399tf+3U41mjlddRa/vcVMfEu4ERBCWu2mzPQ0e4JVh
xoG2FWNty2k5YFAJUqAUoS1jMEzwl3j8x5mmfWsW3VBC+4/8bMnJ4lj/f/IjlYGUDh0+uN8riefJ
kssOqQuuDx4kJ4J5zGB05Rx3fchrq+8B/BH+FB4F8ZIkK4aygKFcntv3CGYldIKpgbylWjoaBRj7
ufWLwG6jJ3jENMvJ2WpjptMNt6E/1oguDfk1aMBKBpWP9C8hvSa0SahxCOUDKCSMQoxrVvVhjU8s
BdMUytgJ9Ywy6h5MPosD74XUUKj8SYjstljsuZgaR44uJ0jq4lvIG3qIAHIvWLb0E1vBt8V67mjS
4e4XWRY/QeVmECcV1MkuqS50FXpFXTezBK1rufBPyf/M4r34wQM7qygfyZhsvzPsQWobwHU6yeut
GLlyrRXt4eCYVRmQ3kYW23FoVh3aNadK4RGJTBjR5NiFqxji3O+F6zEJ/gz9Q44kLvppygCurpa+
zVcn/L2x9OJLmbRWpgayw/+VDQKgK2sTQo45z/PL1VNGzpcvbChHQfcaC4svMPmV9lo8wwFFengL
wHlSOxB5xGsDGSvtMJ5Qi13csTnyxZzzdKYcOx4R3q0C6rgjY0ui1p416W/2HR2c4/wX2QPbgCcF
Gp439Kn+ZfyMt5RLTCfQ+H08Y/057kJeiZTmi1w3nR45WyhTjr/J3lSujGfSj9OrrIGbCX7FLgiq
Gq72+KAy1RdnY9fPkvfN9Vgra0PZHwRa1kLc/zEx7CgrJD+JDIsX57JdblRVcnfFkWN6XVLC3UiE
RCGQEdiDQWa2ko1L1PhL4hrE/+X+Pk2bK0mz/pHSL4hrnFmj8G04Pm+Fvm12efcEITv6ANqRBew1
fNeU3d6LPNEb2e+5JG/kjPUn/7JxDrSj02ABQB5S2K1ua+g9D8tqsJ65uW5j72evN1QlECcezYZh
QG8whI64/5zMOdxKaoAweUShlTUvacDbQfe5V1mU9qENHkIgLnV6yfHGhJfEjpM9iWazL526vp1P
HzC9HvETV0OoL9kBLROFFnY3fEZTSBnEy78uqm+8ZFUr89dqBxJafqD1hH6nC9POFr+1TisvQa9r
uJyO1FlMyL+Z7k0jvLKASrcYw4G3wHjCXlt8moWkSkvG5w6DXNqNpI21ebuLKXqeqkPfc4D7UUnD
Q27yEG613kIex15nsjlG3skqGbtcXEmLkDFwLcdqp0g7g+K8SXEluW+1HoZgVDXYXWEZ7r0dcs7T
O8RwDamNX513KDxem+0Qs+ML3DhnvTMKY2U/BPtXinds9ZxhOAe+Y3+WNZU7B7xOkar/CPcamz5Q
BqLriBoEPNE/LKhdhGKtsohhJjW/eG+qphhYqygff9g5wR6PglfOG4a6j2G+r6AdBYldccAErx6n
qp4J/g4OxT27S0R4tsqVIA1MnU/5EGHquUIXC+hMyY/LRqMnWE3eK5jg08v+oRNukqHkaNKAhWx4
1dutZZHYl9gjmWqbrXyW4dg4Xs0zAB4aDxC1MqJ0iMiN5dpc738owIwrIrSVq3H7Hw8mPwICubp+
lhRvIaMiiL+SQszUro4dj0KFA1gA2tIRznQWuVFM1GJKaez098WwK5/kwL+PpNcuernia2lYeOVE
4Ew1HFae9+DQGKUmvOkfAkg3yft8KQpaJxzFBy5bWd973MORKtU7IbVIXrCvNdfpwYJtw1RgA2x2
zXRPc8xIeQG+RRCyckTWyAcgyBGhkbKhW5RKS6XBYb2dkr6NEdIQxiUekrMRbroAsAWRtWqu/yMF
izXy67tnIT0cUvN5EoYxGyWBDauxBwgprrQjbioqDdXoVMuyCZ4anYocSPajSrOc5UpswTaxhVBE
l92XYWhyGampV019bGJ10KXCC7EYh/lKtbT7vTu3F3CgC/j61ZKxHCLPalxQNDsW4qfDnWSC6kAC
PvQ8QYqtTgVcXCDJMfj/bX7laSqJukPlbeQN66blcqk9O8c5bdSv7b9MoEbFx9mesve+1wox0oLd
H34iykxVqLHcrTLOqtKYDsLJ9OY8D0WPzFY9V1jOZVxbFE4Fupd/PAO7Xq/aSLlluRkxJNaVUqvT
ycaNMuOfkN2tPUFAMxR1XlOG4LitzD2Wq9uTpJPmbtIty3pA8EsfsWI0Rp2rx8CI4QLzG9vp003w
L08D7ocG2JyisVDmtoVoJNkpeUxzTdeG9kO5A79DsUe9j8D6IvJzh7+SiEIBmtWR6bQllBg6Fdss
godqrZ7Q+/ncPP1LEcWxTMiJFOR8rWu2YADo89p+CRnHu1Ex+iNe675kj8QLOP11Fr6dIshH0yQc
R1BpYntmbGMg81EfQ6SUrVQcxZOJyhCzcMJ72RKhuvZL0slBqfuMSjjYVX1czuMKKoXrhCvcdCMp
8JdGX2fdw/7QzD9w5z4aWL8a9mzBycp8LLxIaQsSTbpG7x3MhaGVGE/s1mThQV0zLbac5drEATcl
9HxfGk4jlkcWevhsvXLv1ZkfvQU6Tgr0B7enq+yfo7k+AHQD2ccy5WydxJvOx4L2QvebS1YRf7QN
fHiW26Ot/EY++zJRGCDIolVub3CQTTL+8cSz9DOKO+VGHGtTpgU387x9jHyJrCXcEyR0AzyHlDf7
stn1yh+kXOmZv7Y/bhALGEnS8zQuS7i1PjFf4ouIP78wDmpBzBZ+Uar1/h5579Xz2T+FJlGU+KWM
0xiP7LoqFxo+QfOtLx8HF//nV1u0zBApcpfu0lrPOsP8hmH8yKHWMPBK4t8do3RIuaTP3ytxLtEP
awfAKo0JOw5B9yHnCZXwoZwoR2GpIJ/6rk7Kb/DT1Vf4/allffrfzuyP336Q1GrQym7rCIuqRttz
F1Gm4fRXjUZGp0qJfZVTiw/fg1Ja6NRocOywDzURYVPBlE7Efn26eEFt/CNtfEEEs11P/Uz/xLxx
OKRxHRZMj0fxIEaylb+kOmTJSBuQcscKBSBsxierClgLYH12VIUiatC6p9NDP9yu18IlbwVcaiVk
mlKjdm5LnpKALxMZO4HjeY27pgmpePPqzsglSt/cbuV02iExmOn42q4g8AFHBr7KHWwjzU2/sSak
4nX7SklqtXsYR6rBiOW9Iy4REFSK0hfeXKS/TMk/KRSepgF2HZMfwg5U2QrkdAxAkD0VTeWtTUx+
88X9RUlIk2xsFVuFCRKgZ2M4Mw7eTzL8jodIvqqOUq9byFBPPhfMpbov+2tHsGTRIjCbJYKJks5u
XJUutv2VB/qD18tRuGwDxwlvwa96ttMlCVpfMYtP604R2xgr3Ic5Tv5k3pTL51yybZjZc/Xk9W93
eEFVF8ibE+nnIVzF30ea0cKkYauCIDdJ/PkghmdlD5puk7BuBHrYct4B67xj1GgjCsyZjEzgpxiK
Qy7HIOkqLoKCW6bbxw1U6ViLeeOlDOo4+elPZKTcZ2VWoPs6NmcrSiDOwUMhlUja+BedH4miCXxH
ucjI2jXXmn8lslsBnOPsBP34QSA3J9p5zXr0SyWozmEesXaPjcj6QyIigOTCkZnxVdHRNBccnCqZ
gHFt9AzWirjGW6KUq+5Fc96CiHCxg+fBwdSTbcoBmZNCBklBY6AwsC0LRp+fHnHv+QxmFu3VVE2J
+g6PoOFjnjkdozHrj8K0FKDQjuc2pQ381FBoriXfdKkpnE5sA+SypspBWpIGL60nsh8xeSunaTTm
HxaecLlNuhIAff/nKT8B9JhSKfxNUdrGlTql863Ik0Anfyd+79Ws2W9Zw/RIASY9UDAx/si3hkaI
wYP0REsRiuwxsrz7r09coIoHHWapRdnHiHh2c3+dQlLmUoRCLrq6tLksJD8BYwycugefTT1j3ZW+
cxIL6do8vBH+d6+Zn9PdIv9MQlC3pOLGt1Ybh5X9wq6qhh5hZYB8b5z0odxrT1IdWqEeI9WjpTtu
dl7t53Tzr4DThTceAw6xACES7jJyJVVqkPR1iZZGlxTcqi7n/ti6Y6tx42BTwg8GfepW9aShhbM9
ptaBedWsKeh7YJJnr/sZ6Wg+XHzluPdc8lyEwXWA4zGe2HPl9fgk1ec0MKuKF3/JNkSQFpe+7jCO
4Yc5Uc5CyyZGWcX2UudqwIxoA/4DVbXDETSFzS0WJgPXCEeFKPlVB9oLPYcZbbaFGNermZ6d5BnO
5dG/LJaL5QGxMoKfmJH0vpC/bnCjYkWnhjJX+5D5BnSCxGo090hKrZnxpDqJPbp8nR5ooHzs4d5e
p8ZUEHdaV9iJLuVtHuPMuX/iyQNsez7tK+tgCL/93Prm55FwCBPfVG39nraMgVF6imn2rktPX3S8
vCfcgpwLjeew9R/kb6dBrw2UFME3BGF+BuZG6UVSno7OrhbXGj/MU67tqcsdNd1fUuPNw/AbF5ho
U8q/MIlEA5OgmhZjhqoiHYfbD5yyYSzul99699Gm1TLTer/eulsaLn78WJkaYdMcNS8XheQoTGg1
etNswxnoLh+2nKxVEnWd7M/gjT8EZemSaPS2ZdAhv5pxDI1G+ApqUbM3q/PUOXUtn5SLg4HhtCbn
GVMmfJudxrZbBitfSyKvOxJZy15/GaT8G004kxKF41BZ6SnUUwvD8fPcFes29w/uvo3e8Yr5yE6S
FY1aw28bvWmnKPUgxRh3u2EN93rEouInqjqh4blYFWXbjeov/Gx93iOtH8RMAbQaY+NxArzl/q5s
pf58VDreQ+4cuOcBhDgYxmO3IM/xK22VXclh306/Pizw0Ud2MhPyClebmGKPvMKKfDcrpleQmNbv
Yb9kgHZh2/bMKCDEhY3e9bztPF98AspEoHzMYO/vphMuoN65UbhW+cXYVL8oI5kjlv+7wJnCVfmI
JnP2G5U5mjk7mspJb4buQeF5VW4b8NEmmg3esi7KB4s7qyBk/ob78Tj6vhL7eXKTAkn7Zgmxpy15
snNRgCs4Qw0KWSr87NmdXOhoBLh8/orc4pA++6hxu7H6DF6QHmmKTSkV8wvNEKkfxoONNQzA4Yd9
HOcZIYXTDiKc1oNDl4XkDNDOPlEqAq1oxRNPoY1uVlrouQ+39ol4QCP493DomoGf8xnaSebErmHr
YWcPYNTGf3txcyNejVkPIhW5zvZhfG5lA8uqQiS+/r5SDx8R1E24lOoFnn84RgaP7L1VMMPb32eB
mMCgC9Bld06GDuIsFcsgpZ//XzqwMJqJP+4pM10FTAtZEyaJg+bZPo8oViitdE4NZobPLBt0/jPe
bXGje3rgZyc+aABXm14T0q0W0WLPIlip0DqMoHF/olQyd+bU0XGBwfvArw4EjedFylqqvs/yW6Xo
ZQF6dUiSR6lk3mIbqEaRduwZ8MeXjIirVU5FHB7B+7sYrP1eiPChiFzptP+FFLy4yWxDY6BGQgCx
lhobcqpNEw1TnAAeBN4j6YBJmrCytzFD3GwI5amBh3O9en+i2zaqHcq7lnJYvJIPSL3phhSCzhjx
ifEU084wIJOtNRa2okBjkCJH/fa/r1I+1u5wHpDi3+kKVa31mM4kPmhqvO524pr3cvhDze7VghGb
18V9INrFshdk14R260cSrBtjEXkqlvMsRqCBCSejNGedjEFyOhx8pOt+BS9QmYZMCfU+PAuinJph
ZzC+JEPWMG6JSsxNG9L2H6wh1nb5hLAmH1Ae5UPR4MUcsSbS37/BX6k6FOmQtEG03rE4UjpSBefY
7WidqOUPYvQVJLaJx5CJ/APu4r9NGZ0ySXgtYQH9JqZoTdxgPS2B7MerEPHip5mWQvSYsHUW35fb
eYPWzdktjyzhbpMqDijZuIRSlxDo8rz00280Us6N6a8MG1303+8qXAO5rxVwBuF7NdUaSRse2Qcx
rMwDphsM4toxLfRQQfOaV30WtWPJmOOsF5QwTJHY2VpiGfcY0iloGiPAiGZLL8nwDGs6l64+aj3+
i3MvxxeZNKLeVm88g/pmPbbonCDRkBRGlPh+LjhPKCimBjV7wrI5v284e24DSn71CofJ0c/dbkaW
CjZAWiHe8LOA1vm8Xn9oUYGOZkKZWhFjXlcOQFUUhf7K08hKVu6bvcwdznG56OO7P1dIFEevuiGg
+eUCnBegkEPmFw8/0Qw2+zZRaHSnBXLz3Askvzcrk/l7kAYyEaYckTN7P8btPXCc/2fyzSsfuRR8
MWO+mZcyqGN6rfhGo3bdAKZ9gbMLRRFy4gei9zSLtB+qPWOKr2jAKrC9s/mTtL0CgP+ecFBCDSlI
lD5/q9vFZitN5GJjxs4m8Cb38+IXpdg3VM/1IgpFv3EJMqioN7B/Vur+jQ1rTi5QcdzCeAGh23K2
Tw9+wIzYJGyH8u+f277vGtuLEgHMyiH6Caglsd2eSxqz2MhmoYJdE7Kz22X8sEMfvYI1eS1UYPS+
frBMrB33bCB+o5HcK5RiwcVptXuqb/ORzFFwKERaxtSeg9yt4WjePVwzl/Cas6f/dE4D8ks+2a7c
72XzcuJQp8j5NkFP28+CojEArG0DtaNva1bnnOWcP0PPRfc03Qx5GytvUMBwAgrWPf65Fi1ae9e0
I/NdTlXzKjLaGerq1CYV2RA6rFnCPXNJat8HuPQvoWYdBvawqMljzjuY/FJyoOOWzGG/MZ59l/HR
o9cI9gUm8XycIBuDUESX/lgcOhUsByXtlZH0Hmhqz2VJo2JcBJGqMKzXC/zBVcSOB92mo37okRoe
u8kAeX4l5ZCPhOx4xys+4Id3/PnwM40G8Rdi1Dlww3QHpZTsZcbY17sOJqQNTEzdnherN1ISCron
IEghcb3UQSbIadsccRFPS91pr5O6tMwZhkEcAc+7KMJAJUABouzZalAQ1KooxWHS2AETfEV2aTx8
+56JB/PNssN3Mhf7QLkLntu20ihCVnYew1FDusW43VgejCoJWKIA/AXI/l7D8GfH9DBk4vRMt2E4
zuNq0gR1VvOoDYxicuFEElNkRx3bXjXxmVPAdLRNbENXKofoSe8QZh/6+eb1a8XpCVvtR2dRWQ3I
sYdvQuivZtYfe+gELyg3MXTa7lkkMIMpI1ZKzjboDzX23ABQPdQ46mgish+S3cipEBPrTYnoTyZT
0SD+D5vpOvvOI2iXq4eh6FtrIe4mIw5LblULzdk2Y5KHGjpNMXCR+W+KczOgT0PuO73GWJw/0ylM
r/UvfsVvhf0GPGyQ1bWeC0O+G/Yi9+tY9s1cb1yga7g2HxgftmrPIzdshwxiyKDbaEKmgqRXRQz8
5IGChy1V/ZWGZXtmrv1W+dlXeN468RGLDx4iOtv5OoFrRy5kMuWs39nAO46pVcD0RtSD3MXEOKsN
kiUAbw/G7SuDQT3aGwh0y3ps5uNzXHEexuq7CymslNDnM+6LtcaVr3HSTw1rNLgV/qNpYatFGrXP
2xYE2HkeNBDlv68uau0wye9BVgpT80Ga5wDnhudAzYk/bNxgo0aqwrimUGCcqOgGSaVMiuPbvbgW
bTBjgudOfRGi1Jya24MieyMQWF6/3Sc1vAbSMB5Uk+/MD7vFzVyy0KArlei3eqZ+Uib6Qlg0VLG3
DrgFcIoYIvaYHHvo+FhPpbclHBlyJOQYWQS/T+0Vmk3UAPQho4/yywCYEsndIHKeC9NM/3fClWgU
3NfjL4n2uwV1xfAbeen0eiuqgK+s+1vHONGtlI5MLW0Az5An5G+CQm+QHGyayaVg/oS5J+mUCNbk
z1hzDR8DDcjAzD4K2fG6Ohkh9kpwusGLKZJvmeEPyxFEuIc4kbCN8+NjatoGyRoO+Z2lfui1HTtF
N+31uEuIlQ6RBMpjAf/Tvz2KGcZb8yFZku4BjAgXStuMUIs93EQIWOQgdhywprNFlhPENT8WyhiV
Fs5J758e1AZkRS877kRgh+vJ9KQPrFfp0l/JhipooYhtzPlZeKvGwlRBvZd7qLoOwjqSA45C92yq
Hx0Ic/5rN1mfsjNyKn4qHhMa3f/6njmevnVQkJZ8YiAcRaUrp4VNOtj8wh6QHI6mn8D3apGRMYp4
f+WyZZcqqvkUpoOtKWZ4LGeOpu1fxRvwt85bAVby9lPTPITAVwjxjnv7NixSJg6ZvgbO5QlTiX3L
DZyHquVy7QV/uC/CwmOqfex39oxDNWOvB6L501/Cqj8bCe9fIrneQtoo4HgyJ5zCcGaLi8xJXdgW
LImk//TmpxHFkFi9wzCyv1MZNiGV698Pfo5N2GcwmG1T/sAdOAmirhWoF4992FUtjCZ8zvhbpcTx
Df/dVeDsBcRW0uilfLHZN8yeeVBJx+KG+vzXLFzGqG2Te8fuUi4g+A/mVJOFnlb8QIejLfLXX2OZ
Nf0i1i+Pbkfrj4xZiUCH1rT0ktg+g+W+APdwXHtq+t8B46j41azUT7HFurtk/Su5ZlfTWdhfpRIa
jiDNJxBm9bEwEPZT1p3QfGsQC63gPYFxomW+jin7mLb9oKp9XLcICOcii0rp7Wficv21MEeMWmbF
5IwgA+uiNDpSD8rrkIX7qmiUVkC/qJh+SZYxExEvX4yeytJF5+0bFvAqpKQ2TjuU67zSeene7ciK
jjqze6EmvmPfF6yfcBgtpF2Q8iEOtDmjS4dMYkuegMIXjnxB6SYzTPD+3FopiKqiOFgLJG05cTC7
VxXNKvdDx/GENNF6Klf5AnFtzYCA7j/hCaTPZlr7jCYJBBmHEwyasuYTLvx6fUKgjo9rNvE8L66W
iOLv4qBWWxURAHZ+S6oMGZXxCeE6n6GUKYIK0zNZEhztFunKwGhZ/EBTtbQA5S6w2NrTInAAL4lE
slI5zHeSS2PP0qyrHL3DWkZ15zTuTaCw+DoObr+7ZVdEfQqxfu9rtJG1I1lnY8kvvZYM43BXhBnc
igHT4mUVYLLrvlER6vWI48tZgO5cx3FAStr0tofeupo60r92EQzb90SQbQSha6Pqgq23V9jTDWJf
xHLS1K9fZsRKx6CuuKzr9cGBw6q8axISSwjuOztjd+Pr+mVBxw+K+m/xqoRarGhBUjJuDsh5qa2+
UqkT5/W/p49QvXw2mtIr154kcFqYeh8Li+P9p0k7AqYEZZLEc20MiRbV6gNbpYehycLame+i7fT3
GJNeA2vk0pKxA+BumkEvc+I8iTnLg9W09nOt/GHIA50P2P+fsgbXqn6gEp+32ATdzhNc+5Kz7unK
JyKdhp+DMtiPqR7bOPZpBw0MXCeVpDZBxH25zeHEWMaTD/YXQkgg4lZ2ibfXJJw4jDGFFqrYq6Zm
vNYDi15XpHYN2u86L6IC1+nXLfa0o8rpRm8/FJnWog0aMtbt6oMQQdK+kbfn+nFG6jE3oFrHlBRn
0JoTmGPKLNQMLJH7wyeafVeeYLyb3vaqcUFreTYnSnztwyGx/u6gX6aSl2bqV8dUj6qI2kVJqIfX
SpJGPoeD6KpMk304TN0t+ZxqBiXxGz4Pf2B5GUvqwRMOFw13g0qPXp+bgrqSpHLt0clCLCbXZXK+
+PoF0S0AqiwlSxzgeI6BtmpLZ+PTYCiPJNgYCL9Y6zOWevC3RbY+OGMTbI6XCGk+ASSLJP3jpJZJ
jZJ+Hj8LYSl0ynl/a7SN6ttMsro6GLsbiJ6XrYfCgejC3c/IWIUIiD0rTikILlURBBKoorJ39J1f
tJ+n5VDlMblPtuUMlIYWJ3eGWm6fcy8UwUm3JkAFcx3y+/ws5vJyF0TLbibaG9yIqtvCYzbQhi/y
3f7KHpO+tohzZdtmqdYwZ1ZOr0+hFKOGjTf27JhZ/XOC+w1TctQs64nMEBmQnovApaOTDr689Lji
Ww7PDvghcFhxQTizljx/TRWDwXFGcSO0bNHUx5yj2FK8XJfXwNB+reaEGyRCn8cSQxciCuRWjlvM
FIoOcTBdz9klPhKecWSHKwCuWTrw/kEpfaK22oO1Dv3UfHpjvYUFHgmyT5+3CH9HOAA6SMIWlG9/
pKtV0QrdX+PfiymR+jt4fVTyaxsQp2oQd6lapbN294AbtjmQ+4bLFY3+4AZsqz9l7B2Sv7irFCCV
ICgsdUKBKAKudSysKCUUHvKDJwUyStmQMJk/DqTfuO58G57aX/jGYDeyv/d5j1YfBgr6VuZEK7a2
Nlw2gKn+TrZmr4NwdheLc21jmBTLAuwR7k4LJRQtrY1EcTT38+sF1CS/OnB34V19mkM1V6jbQDUG
FGjrJa7kWlbqtRCK82uao/wmOIaAdpoZk1v0LX8I1REqGvpcRch+x30ygveRJb2spW+mTwPg6HaY
Q9p6+L6PK5+78aEFLacVfi+Ch4uHUjgLtTJsLFgc78909e8B2UhC9dL2GKwjU38WQEJ7shTsCfoo
vQcKw6JrvJ8nel2a0RsMUHxdPlULqTLIb2jkiyqVBcsejp+kb3sP6t8sBpByCw4r3DQr3Mu4p0uG
VltrxPcLPLwcl9OjywaSK6VnJSTMcDCPCb5MhmHnnNjY9ccdewItHlu/+gx7Y+V/91cqukHZ9Qy2
SVzko2IWQg5WyfAEVVrnuK+hb4VJVkVkILJa6q9UYJZpNjxUsZFunrz/lkPBwETSqKPmkL3ljFTi
Bo95cZTzkaDS11a2USN/oVX7Bn4GWCCRqf61tixkSvaX7GQNhdgQHj4U2CqFNW80xL+/tz3RSXRd
4BtoCgfzinlCe7/l89AlWAyvFE8QGEezDnqmr8CSaD5H1X2dryz9YSfHxS7ytXqN3cy6+6ufzaFL
zMzx6DlbpQvzGUd1cNSERER29ItxOXB3KuPL6z0LBYggI+bUVPmtJlUElpqxHtrfy3uTlrBH9uf/
5UQ0l64bcgU4XsO90GcvjjJzkz4+958O28BY1Wdp7+0SrIMhoFnQ2sXa1wdJnRWA2Fx0EgW9FqfP
vlR5ZJz4dA9khzCfxsYz6NhdnSmc7rUsOM0m5Lz+dBwHPlg9O0C2Uu9SiaWzYZy/iYOpOQg97g0q
MOmafPf5NcunalDUg8S4meqjSUGeUoK29Cdxq8bJENdpWubQ/pjYsXrnBHnBAOeyogSlS4OC14ER
9mZDT/dBJbSG3rhE4UPJ9VvnbRFTAFxg1KBsuB0iLhl6ZPY3Hevucf/a2soKwM7ut1SFnfajwXju
W4rIORVbk0PTVpbOfqo8z6t/dcgjzCKLBxvTlWSdPMQluTJI8q/B34TsZoFrzou2xsw1DGrIz47f
wDEUgs2kv80O5bbf8GgLhZtGJoEXPV1bLIPctX2yfEMHMkV7CTBYOifr7o7Ph/jOrDYnFCIY5ZsF
xkwCd5OeBLPC7WiVaM9ZhUXKxjyF8bL5JF0krRl5yA2mG+tP2rYgbFSuqxTvmcX2LHOODUL5a0qv
+lfCkmTd9WKcehO/DNHzcmXm3d1Ra0lx3r5o2QqmjAq+ua4tsvMzRtgrtUuMQJis6t/y3R5r9ebb
NAmFBbLbALaKRGszKRvhMy7qp5kPYtwF9s3dRM0OA19YHAgilMm/y3kvduUoB+aAjmHRjDNOmVUG
RE2Y+sO0jpvttgXar9No6NpTQERwY82Bm8OKVsTr3OdetXxI0Mg9ugHTWBFSHhCdMXJzMV/mT4di
iHQue3wiKSGXMMT8cdqo2P4BDz1FbKiSz5OfuRX1SarBRuuZ3TAaLFtkFC5lgrsEJAwd0ljS/riK
1NtE398VAa5tp5tOyKGDGSZdmuSEXTL6MYjsRW+AMbesJYkfKkZICvSo41clvaO7oLuBjuXmAO5e
bdP5XhlYcJN3HZkLn8eNbrIjMzlTSZ0nIJTGC5wtREpvJp+CQAwQ34ebqhYCEj21I+tNWb7Ujtoc
acpbwsiE88zPaa4i6QybUmJYQAwtvFs/43sTaUZWNqK32KQICzEG781jCVxeOGuu1un4xig4hMwo
/26ikLK9pn2+AB9ca6gycH+Gx9QNzNRJlT6EnqbHoPaaZojP29CGYRgLVVTVXFNPNSX3j0rZGkyc
2iTAtjKEGh0H2+Zss9rkRcn47QogzpJqhBqYoE/Rv6suWREogonXZSAmAg3u1gKZjJt2rAtUdSVs
+wvJTgTXEAfL9H5ATyRBzgLLjopQT72qHt5LuT0jO5k+XJ4LvIQp8x9Jvr5JlIYi+I0vi+m3SAS3
zxRhTGlgIsFpVQKNWcDb0FMDmOO1/kspYkZg8J+v0sBB5/Bm6y6vpoRfVchByefub7Nbyk3+s+PC
oNtSdYDrqxrpTdEOuBs1mnNPNyaIZKzt/NbxgSyRApBJHwwolJnciYjtBqKZiXqdRcLMjrGpNL8s
hYMUC46FBHk67M13q0O0syC71seywfHXrUBM93ZrDTYEkb4+lSjX7m5tXDUTvXY6f2Qh4ck5q7cK
iNkjCisIIpgbS8yeJ9K8TFiMJsNci5LWoxhqFuaT31b37B9kYLTyXC/9v4SkayxfiVLg0JwSn/72
69mpZtM0peUND5DPUujMIrdaMboCZNaVXQbZfYAIdLcxhk5ZGzlM5XWiZXseaB9QnQceRn5ppja4
BhiSM4clRGXMSJro2iV96GqAJ6nRy5ZBlpczbc1nIX60uioinUloxeF6EmEigSB1N+j8RAG7EwF1
+2SJnz8xfrlOQZPGZyTYNB3OJ4WvNX5IHVadYcXk+uUqklZDj7lrBJlxA8tpimA/2/4e+ff2+9Uo
DZzQtIiG1/HAy2r0u/E/WXupIqNb5hjPL6QJoBtjsSO2sES0njSeOep6cs0lplTYbBFVdTStn8YR
ZfRxfGTAI4WJ2YlsXe88usvR1Ama9UQi0GGuu/aNy2O3QJJpAFgqncFaBATDZup0AJ3JWFQqwTmR
06W0p4tXrtq7cw+yuEcXW7oV+0r9zoWZ2Ii7EOiXJzn5WrMLTGDyjF8i+gYKaP/bgvYUsXReaPDa
oXc75jzC1PtpKGTd2AqxGCPyhK9c4z2mmnRxHNb+LP6nkDc+pB0lTlR0Mc8wsIxK7c1OW4+zSIxR
owrQnSUGbhYlXjVlcArjsYs0E15zurJBmf38P/Yh+mmRk6+9iJpPSt1eW/v0modIdtrVQHboy+yf
3VCxeV8nFp0lLkPP6i92s7qSXzLPsIJpxxfDY4amXfNllngB63rsT+8Rik/KVdJcDkoTBV2nov4A
cgzBjS631++YJo7eBUqLdfnGfl2dtJ9lqhcJ5bmjFm8eBROh3cUP1+QgsHutvpW+jn4KoSAICemo
Uf427bxpSU+7gPxZ35xvIxUrKEkQWkl9ZzG2UvE1jys/WdRyA7ec5i5GgFxZg28pFzR+KQJcbcGh
50Xb7Yy6Efrto5mkquU5+RWAI85/jlw6sOHdr5aBPJVazN6EMnsuxqB98lFaxNO9dzo6S3SGiYOB
BWZOa3Ysy9U20wEqxf5jw1jo1q8DNsmO31Q+KZR5BleChZryjdVmXNHoye0HZHc3FdpAMu0qAMqT
PSOrcXGjO//w41khCmBx98dDuQY4MxAexn/czRk3Xiwept4ECHtZByr4emLGcNnqEsNhOCO+PCgy
bBC2el5KeyQCgbWIHOmW0DXPsQH2LHwEcq76crg50nz88Oozde8sRHt8bsTLp0gzNbA9WVX2W8r+
mKz3ptM5VptFC1iAXinczpeeVqZAQ7FJwtPFO6XCnk91LIdXn9PCXY5Ln30/DECbmQKGm2do962l
ji14D5V1rYZJMaeSjKuEzEeuiZG72GuDPZghCUhOoce24fGtN5FSUR7w5falcqdeoovWnEX+tvLt
3yuBhry69UkA77FdOoVK/28eMjADD4yp/IWEKd4AiA/srcRlf0cyrjxr6RDmI6CYlaXfw4u+GVqX
Whp/nF7NHrD5+6gCpTPv6bnOd6jHThe/AsYDX3Un1oSRXYf6N5Iu85Nh3BB9DNblWuWV69qDAIro
9Sng9eHqc1yno4AHUc9qOg4nGGovpNlQWloVy+ZTMAfKzsItDF5neCSPoSQ0MlR973u/Ltdg6qqF
orEAhIMdREsYIZrK3zfbXe3NnY66bdnrXzziH1/QJaEnMYwc4BpI3WYFchfyMDrMOt5klBHcVfhj
RUgqcZhvE56+HdzSFGolQI0Gh7DVueGDRRdIqhsY5SY5DbWeF3o/HkV6E+s1lxVEdVNxw2Jl0DIZ
ddM+KMij14nm3IRFhnVF2R/ZeD8tkLl+ZS/Evk6zgTO+N1idRHzz4AUFZpGLG9O5LQ9qSIN+Jy3j
/dcnrrFwJs5xFUogMpilvtfehOmMz/dp2hkNydkqHQm1h6gXrgFH6t5z6U4NcksyNHUvgPgmbBCr
zhtjnXeN/jMzUAC6wxyDQvMZXSVJ4vGpL4gFKDLPUBH1QmT0fZIfD1dT5YboJmlnfDLHPNJxUTZ7
RSip0QiUtsIMCljamSS73qn+IV1H2rhekS0qR5Gmw1fGCaGE1hycRjLie5TDaqx2oRo7HaAa5mun
B9+WRciezFXtXpUkJWUagOzCUe+JWgRgHZFmkpHA6+I4hV2IaJjqwjAAMKEidcgVwCBsRd6uwQh2
fNe8v6MyeCdnZWi9qgfdIRgZLiQux5rwrrXwW5MkTkbAOwDPhnrXAsSGobG5kWNzUkX4sNoJqnHb
lIQ1jB4UOpGnFYZ4Td8Mv8GfxnpYtO3fi2IgO14gfSB/1f084EUzG2ptvLUL9DaUNk513uVbAtNH
jZTP8DfvUIFa9xirzOHf2wzSsofsJDnd2EJXSuyRnNwif8fRBUMcFFLTbEdswM3wYB5D/6N1v6YL
I+0B0astCa5dToWrF1MeSoNycJQp3FTrvdVIzDYjs73PoiwqXZCW5loBlxhN7vfmV77nY2Ioip01
VuZim/3G81MBY8OLJf1Bdsl3ut2V6AqLkzLmeskJn+unkY80zVGSBbpAkYElg4i1sHsnfMb9W6Jb
PjrdTzd5lrV0+ftyK3OhoLw++JDIhgWBTYCKMa8FIQrTDe51OKXspiT+1sRgwW0b4bphA+wuEpr3
FPnv/+LUVBrJxNcZ9/t0x89Tcpi1317jdZs83iLjmrxqJmFji2zBeSgaeiD5C7JfFeZoilfs6JN5
rmLQWmISZrcl9pJtrmWqQ+KHMACq2YKc6LPPk09/o5g9iicG9GmgEmBlG7dUbvfMS6N8fn8tVo9f
KAQ+q4dXEUkbuPr38U/2n3Qpns31Ka1uzGYKC6WFgSUa06+bnxN4hiwW9i0DktQBI23OgDgblqh0
rTJ12Yv8HhGXqwJooonfJgK4JBDx71KluR25+LOyecdxIOam3zJ5j4wZmeEcpXNr9neQxvcZ/IDH
I8lsFEzeDRA+DXuVJbrCTMuIVSwGN/0KirWWmFVLIfrVQfwjGBH3WfK6i49BXFSOhIVpvycvxTvX
aV4FmIcD+TD8XR0sKjSL23W9vl2al4UmlJqgmC2iPYHU+/yn3UF/L5MSkG9QRc28TytZ/FAfz61x
MRqHQIW2MYQFp+JB2ItleRuhIC9caD36iIGq4dxB6L4KToL6PaI4R+n2z/ZWVaG9NZ74ofkRNBy4
CFx3nxo1iNTgz232GmDX/gyasSjEdlQP9MyaEJGZZUqN8RHvrJdAO5lE8Nt2Fp83qXWBKP1jPiAf
jly62ZtJxnUx8EElrtvcr+TkvSts5PgPH+YWEqfA91tI8Cs7F+mtL786lLCpC2XaarrVE85KS3AK
cw9LsM1eojqYDPIwbXCkYaGuAZWydCQa6nDGnDeBysIJZPF89/vTiDtk4VKD13+WN9RwaVhpfA3T
oS/Arf3B7xAkG494JPurfWWq7pDxYDRfz9U+UJkUv0klq55LgBGAnDFZUvRb1UTAIN8RCp92HIdx
k4K/Gc0LIOWO8ICcWTTDbkMwTSAOHanshAdB4R9hOFhAjNLFx0EnFFxApzMyCYa0M9xEHdPLAZXL
OQU5fRYMOgS65FjKE3sI9cZUYjenFpSNhR+OdSgukIjJjnSp5YDCbcMKq9536HBE3UdtAa5a4WDo
CkejFWTFL0F3bAsSo/s8fznfLs2lxph34LxlMNq5LxcoXDVVCm9wwtu4dFnZjzkTeh9NQX7SXHiN
+BBUaVRIWvUGZ5pDdhczzSjhG8RIXH8szFsTGRJHchCeH9sXVEdJXWz+PODHN0L8dFK7JSPF6ulh
FPFizqpeN+zU7KHjCuDnKeihFPK1q/r2LJfQx04kZqXcy9doo3tBDBevgnKUpQehnobnN0auE/jj
O4XMuMd4nSFVp3RAGN5855d/UBD4tBzSRHzh8j/pwEmduyenEnzPXBsjQTM6RIkPUVCAEXVygro3
L4JjoRRNgj3gbpxqrVN3NZyifshMZ399ENb3YAcoHqrT/aNeuJlG6LyRguANcTrqfFrZjxrJP/9G
fwBxJj5ZAYXEAd2XrzWWZhmGL1vkQ3UpGzNrX73LK9XcJcdVGhus8Fh0xJ+u7vGMeebMok/1zrOY
l10sYFImMFk3PjPcntx8NyQxEX37aXt126NDjgzHLJGLzqGGCFgXNl9oFpOxOwhgyfUkSjrC+ws8
b53w+pSO/tTOUpFJCY3OdKuoSLAGKhvtUv84Eo+qX6kYAn4m2W36XyGHxdn2WdFQQ20rlxgkBKM0
o+oTihbIfGS/gcm0rrtQwMS4GWMobRP/vRRS5n97PBzPG7eOQ5Asfp9JkdhbDwl5FFt+y9zI75ML
VogbX8NPUuimtVChouES0tkjWeqBaTS6FMj6AuXOJqRsQ0RA8ryTwFgMdDg52pPQujgVKGYHVCeO
IX/MVuIbkVsbX8pzwVFpzdJs5Mli9l6irQQIjHhLHskRwU7BD0zetcUQzikCodz1mb1x3sNXD1yE
WiFnFXDPzMpr5KL/CwD/rLpWGy4ZdM/4Mr5QSHI8aZXxD+sAbEEONbtwPSISxeMiFhYHCV8DGHCi
sSYYF0yynZn0ZlAT6y+z9ok0rQfr5Nrpi8JXZ4PSct59XrKk1Fc0UCp0Erglmozx0+dABpEbY5x6
pD/kfLVlDtpcEy+NbsCceKVIp8TenqqFzIC1AJ+SctYXg7pKJpZMuukXMYUoHqNLgbr7GIrvi+Sp
aw60QkPO2i07ks5Z4BBcbGIheLgT0H7kPoKtGbwCNLkSrevfoJscfdjBB8S8Js9qNTAJ7UPQnSS5
am7XsJVAAe6CSpherjST+IXUS+NGGO7TlITVbcPTMMwwQTFiGWoIeV9bWNends0Q3hskQcazBFGw
yHzcCT7lEBGCPRPV3mqpmQJVADGU5Eb+Agl4grQiKkjWfLN5alKOpryT8mUgQ73xNAgp0vQ5Ppzc
h+LqYfJluBaqsY25oB4r/Idz0RZ9vPKTRMGvb3/vLo8w9jG5GVLqa/DDdLseHGguIH8pYiannuiD
aGKWxjLfwxgdNQ4SGD6oy3ELimpCDQH7wBCukHmfFUL/mKWBB0jQe+jb0KsxpuN3h41mq8bKE62g
5Wg6TkwGMMp/GJEARX5lBTiMNOXoABFi2JCR9rtA5A97s/g0ex3aeKv1+oTHI1LMG8QzJmp+9SbC
PH1DmPtEaPNkfwSmxLB0ESd8ywBkDI9sRzKI6Gu47ZhR2aIGaPe4uzZ5zPKf10eoal8D4/h8F+h/
TyQ9mIbzeLmlfJh5EsNAWG6kwzEUStQ1y5h8WQLd4qQ4tdyoKqhwf/xs3lQJs1zAC4zbYNMYp6LI
x9yurdG64kH+INYYysSp3QGeVsVcr01bVU017GFRMCqMsLN89U8ElOIt1y32ohkktR26fBBBGwVP
NauWktEdmIi3phIViSCesPJUJO7/5dDIRGmZcHuAfrRScfSyXI5YMeS3owXmrIp8DwSfJIqfjkMk
qpNrfADmDRiOwritG7Uv5tInGis4rxLVL2kwF+SMJK+q5Naf2IpwmD6x3+FdI/Sf8DRZBGMZoYHp
3I4ORlu4Q9flqDvMV7ZstgpTbzx1PX6Uk/qypai6sksjyirzK5BdOhQW0hnsnq5mV7XqGJEDGORp
0m3skSqsX1s21BPhK3mCoOxDRS0Vg3ePK/jJlxqn25KhI9FkWtArHRPjSTOPzMh+JdSDl/Nf1zlG
2Q831k076juUXMV3b+sH2GoI8BxfD7ECf/MDNaKg5JNItgF1Es54bFkrbvRsDY/fGZMR/cR8etT5
+g5/4vlOa2JdQIz3V5WeqSVE7B5eooghOKsapK79RKLXxyV6VXD+WFCyWgDmY9fVL4v9cWUykZ7h
GLvS/5IXOa7xPLzNQVAmRZIrJpEGlmZlzoimC3UjL5SD037r42WK2zqWCTO2flerAIiGEA5HywQr
ZCe47Rimz9TtZMb1K1CAYAGCBhqEC0R5V08gyMVPWez9/GzxOZRMYVihLpOKpEayt8IyQz+gVCLu
zADjfcoXlkR8ktjID29butClXoLmjYW+OnbInMomrmv6J1YZXtXEzBW7gdoS94GkGWcn+W4kKdUY
N8tndANl1dt5zT/dX+gko4obnqmlLZduCKU4FZju+zUYbg70WaPMDSbylEpG83fkdb9JmupDeeR/
KL1wT0hSjUREOfvVMb4nCpuAxuYZKw1bS2i9YEWg5tgF6rMl9XEFPB6V7l9oYoeJ+yhpTJbStYDu
UJ6UVG5dxL7INFa5Txtdro3PwyJ0/acR1n0/894D9XPhXB5nNzCWDahhxA61ChWgUdmq9XP6WH4D
T2rCPa8HcmCKcQQDN3NgFYcUVnXW0991pQ6rNEN3mndTLFo9+jJTSNLbNbWgMpZ7TnxZbHqMXdQ9
aoaEdhzLD0n0Xn3rh8XdLAK/AZYnchxK/WyuG1owVZgd/+syubgqxBuN0tvOkQv9OVM/QdNiAPqN
6Q6Y0R393WXyFDUdXZT2ilQ0hcHSx2wN2EnxrQQPS4K7ccDTQBswNtZYVh17k8sjKaQ2jsGNMOo0
KQPvusxY37DmbK6SoSLK78OhLIWozBIDLNihjSOsFIXhyBGoBNsfL/l6h7Dp4PnhqkC8xo0O5xka
Uk4UNa7EuEBZBTqFjC1oIBKOTkl8j+aYYxLVEDjOqQ1W9fWKCU8c6atGpQdivi16sSyMBI7GJDjs
yo/Ghi6dVRX25YF3PdL+cPNGoPpzs+I8EgSyKPWlPNWY/5tYh1mNowkhmz0JosS8DqxOhFwZTpH7
NfGMQ8FJPgAnTZUY75EyZbj6eBjYfSpxbU0RUN3fG0G4Aj7pwOLjfunAQ/g4/52Kv+CKyZ1If4iS
HKzmHfqYDRR7vs2O40Z/QaqgxKJEjcmQyHls7NYs6O5Z7eVo7f+W81W+nh+DsBTmzzlcjHohivCI
TWItI4W7L4/tsr8WI7qUI1+3saupTR7vTcc3S/AXoPg08FK1tt2LZ7SoCX1JCH1MXwnIvR2aMNIn
fTJCao+oBOQVv1vC1uMr4y3zd6t9edznEiEl4eB5UQbmEfFn4IU1JXkOumQWCGOX0GQy57xTcqHE
n17335VJdcXdsqncy7IjblT7Yf7cEINaAMtq3oUDi8LUt1OnH8B6F0cw+u/VBG8ZOoU2kxM6LL0H
pMetgLpNi/SMGL6jiM7/ThYnXAmbbDWIE95NlXD8AAdeO2p+8iITlrIk1I6Kx+/xPmYaxP9fiXm1
lMDv3okOD5evF7LzKQkRnZUiALl9vLXyhoVICb+5hYPn0Sk0XNT6JtfpSYVFbFwLFvxwHS/7Vgd+
2EuKp7L6brPSg0QZptK2rcF/hl06ypaPkS+nBxC1gjk4yLrH0WwTOH3skcuLUa/Ict4ypqyFxCEg
aip8lFAZnbz29j+dxTp9e1RQrLj9bub39Q4tv0xqikSnzNCRIP3B1/JuW2D5eVrYRNQkGHSjj+ms
G9f5X9MN7k7g/6q8pF6KPD00ImP+vHEpVPYl8bWI48I2JH6PIhsNNnrhzZOZYt82SXF6Y6BBugW/
lV0j3oOkkTrUoZidh/wj3Pv1BGRw7mlA9WhPEzxuHEQv8e2/465H/I63cC9te4kZnHqot1HvHh3j
cAqwcnC+g6SIQt1LVFQqOlQrx27mibfLA8N+m/JxC/HMKVuV0VD+I6Kkn/5kSsH44auX8KsHgqMg
E8JFco2I4hQ/qenztiLC/9iwEDvj+zVAguBRXCL2sFaWpLeJvbng3wnIQVsSXvRjHYB9gxyP9KOP
wti25suY4Ox28QGuuLqH4Z4KHXhg2nQYl6m7ZyDS1narIJ6eEWGZgcZSolGkXuqTJcOsKBD4Trfa
amMBq5q0SnkCtwzzhTB/1T1Ea12IKDG7tLwcTs48OHVC+/yl3kPn72O4YgS3BgRL1fNdoMpkZ+Bh
PxiLoBL9guCcXjxmO/WkRiww4kLwkS1dRrBiCEkIcmkhinFnijQLN/cofsaUAbYr9ZcS/BtQZiC6
XDNBXSN0SQBxI8IyCgbnQBrFS/LSqAo/dVmS9UqWYJ/7ADr5WOsXO5heETOkMkzloxnQeeNSJz1c
4yMCmxpNT0O434Vx0MRQ3bjV28Kma3Pw2s8RHKTtou6jKUBnVYf/WiCnn81DtimIeiD3kKv/QTRw
PvFxDwMGTrnzmUe9zBdALYudMPQx9ug2z1wcU/R98BcVmVxocFZZFySSFQF/dObDaZp29nS3SiTY
ehRgkuSRXPJfELLZ67iWf9a2Hl4FgO/MkpEGn3A9KOYbLafTD2Rw6luBzq/BSVHyYhJYs6bB5LNM
4yIln8ysq0WMK39lSs5nox7J4uG1gjM//neUuzjGggbfonG9NJvsrabOx1E5Y9TIIIGL+ji52axI
oNzORYMG0ga4bVCxacNN+/qJ6pJMEJV/iRhGF4JnJGWNy+afxIubVzkZ9stAfgifZ3DM3c9vz77M
RV55GmF6yuclC7/3AjxgX5nlboXkJJAGej+gXPISXqGbc5xSDTs0R++b/H5kr8ISyAS0zF9tw8Pm
yMg9NC7Ii9ZCoHBEOsJct3oICzxfP8DSL314LA+LG8E80K6HSBdxDt6GXVAhE4dWobe3kQd/w7Ah
5aUQImkqZLYVElJTTiJzeTR8gxtGi+muQ3hJbwddjNcoqb/wSQ7cL7H4Yixei90fFjGXpLwNAsd0
RTXjn5+/AL4rt1uM1Ol11j+994x/GJad0tA78JsDWUw+hIf86WsV8exjscXrT8zOPOjYH/Ew5AL1
Ua3SAKCakj8ZlNZvU2E1jmSyybx7fjZkKtOtmQySrQM/4g0BWCkKZ9S9tXzRMidrIls8BN61F8oK
wWHfF4LYFyOto2a9HofvESeIELKPYgkiKT6WPXDPAkXzlAmkmC0UEXZpX3vRI3JDEfE13wBkeO5+
6/o1Eg3sg9QZi/aZ0QUyw7+CEZqOwlAstC8TGxCboPzKSS7SYOvUzasHq4XLmDssab9E1N+YrTCE
XEHCH6QhHed/WNSoyO4PehtO5M7WcijzQBv8pr6KF2opJPHMtQpjX3ffTD+/cam/b6wfRi3o6siY
jIdY0GUDylSUVNr4bCfVfvV2ZMWZZPbWrNPOy5yQqYIKAfDN+oe/j8w0is1CGjKqrPEsgeRdCYai
sjSVuwLe6IsFgaYogl18qCY0yLyHIgK3jKimGjxORe88Fv3fyXxTKqj1mAU/UoSnDkm9g31lOeBU
AzG5c6B/Pv7O2ZxuXw51fOr753OfxZTDuOrtSDca0O21WcEPcbqCUp9chmEZrdGxMh1eRb7HuWS2
bJ04duJHW4jbPzrEPOfplYPD2DPx5lCa5IrzwEiLAo43bsq6v0txtm3RLUyxyoXIcQDPYzNpnaqo
TB3hVEQ+xmG2xnnhjDBKhKyqEmbCzE4eInox8ygA3WmF8Cd5u2rhnQ/wEZEjo1e45J+l5iQ30csj
z8e6eUYKyHzDLFfEOAg1O1Vk4x8wPqe73oD1gRBDlWhrjW92/KDsGpwmWIbVV8Ua1QXxQzZZpBzN
xPn+HUE1KMcmkEG5wwNbPo+xJScTjYA0aDip8741Fk9pozx9r5vYIn3BcW2cLFHugpj7Kd4lel1P
I8WIvrsNJj/7YhF0V9QNBna8eU2n+W4wWNLYEIYDKGf4/xea/f2sj+3oE7ehrwWC8Va0/fWwf28c
Brpz1JTQtMZy5Xl4aivPZM3iQbk+FCK2bGnsVUI6qz4prZL/TGoq1cnAj+7Pc9RxAm8fgt2O/8KI
nQ6UdqZ1PzpE/sFm4EYFusdxZTMlQvc7FcPDSe690htlxXr3R89VD9YBr73blAnseVp3jQnCO69Q
z+APgz6acU+ww9cppQhH3JiK2HnRBoGhnmLQ1xdIFRqrVM6MxdaXDYL2PXqumEVB1uTJVLMQNW50
JK9sfML4HBHGzl05QlUKAfprsrc7aOlTmJV2DUWuSRfi0EooumaK5VKmVaRlerWpPv+Bgi0tsieL
ZyBdHoAFfs8xMp3+9fl9A/juygeii0u2ovLtTnuSW7pfqj0t+MLn25FzL9WoTCwYcQ4gxx9GAWR6
6NbREtdbQIGKkPYCFP6pHh1+vtzbCQAaVGqTSbGmcnNoF5SMo2n9GIWI+UJqtoHqbEJZo/cybEXw
QnQvF/hJsFcUTXm3ri1ssmqbtMrSCR4fIzWOgaqnb+pbktoZ8GOetJcH/gzZSHhMuwzqg6ez2Jzz
wy2oP6ypFW/NV1pg8k6DJZ0TM5GxC2SSeYBY1C4Uz4K4Bjd8OJCJET7MOaEITsUr2hsAiE0BjBfo
P/US/VAD5ut6nX2grEYKg1yAjkWCaw+HkdfwzsAvNLCGFNFoH2hN+OTeyNduWwsrOQmncVcOzGRD
U93w53lFQUQuVx3ZErdmLxYjiX1nfmu2XZyPNde+AJMyaV6t9WMGUyq1pTX+zTVvJobrxq/tfmIV
a9WKOxbsslWXP3OnF1quc1YzzNPK2+uvLanCYslbYsqLpE3U8p8f0JR9fufVqoHGRtLGXh16dBub
zk8JCf7pMewSpIGtHAP1Q/YvmiqFZsPnPxYJ11RPTy7NiTj6gNJGLs0s+LkgB3Sn4tmPG0+fipoh
n3SrTFRj/nN7AWsm3qrojYj5RozoWeOSV7fz2IyNIu0PygZoB95dUOxYTSjCKPapKRK45X2UgwJr
VfijxE6OWBjZI5vi/RO5O2wX58s513xlOWBEEjtNp9tiTBsFbG/fhFoXu41OJjKsg+DscwrAEUB+
9FTkl/6sQVMuEKSOuaBwrwqaiER7xrwG3KBMZJZ1rutE8mOM5Fn8JJjs8xah1+hsoMK1BCC8HLvs
Z1D4KdE10R3RvWVRs4VuaMIMcB01rdCgnV+immquRPvh/5pL0V6B1iS04+I/yGNS9KN3QouZbVJ1
KW0C95CJxGc0mhqIyH840bp2t8ebQmeMF52OLT8hFOJe8EXexgz+52JVVmi8Vw4TqvyGkMxTi9r0
G9yupgDHLwf+Zheq7hPGSErAhgVpTfGstEH6Nq3CCP07in5iopOKA/Ce9jzByzSdQnWYvATTWMEM
rud3VMfo3sk8fupzHtpY+R/vHyZOEG3mfyrzWQkUiAafksMyFX7964NGSvD2mj9X0gRFNnhqk8lS
JnFYk5bASgum9K6RiAEoHywpgJ89Tgy5Cv3b9rjOZbkNXdB4Y3LEoU05liTIir2Zaoy4NRFsoatn
l/pXsHXv+83oN4RdjB2vgfOzTDmQ82u6A7csOXU8nM+aw1tdKTSRUgGtnD8ga376Z5e9NSLgWdM4
HGC2jjumnHWZkUdv5bLedo8bobPVoWRcG/f05NbpMYK66g9L9fEA3NeSmo7oSvr0dwt1fS7kn/zc
/gLkFGliFqCkyISqkB37mUWG9B0OyX7oesainOC9JsknHBI39VzmLyfRVvNvzRWhLx5uwtt2wBMF
YDMf2pUu5MC6iyYItW9F2RQbJlYCcSdDXcWgK7mcsqep1BEm8oIWW2YR2g2q6MWRiFP2/8ckXJvj
O6XrF/78V5OrFO1D6G2bpu1xOS/74PJYmfNAIr3KDm59BadKJGh574U2Lw2ijAD4Zk7zH8isx8xs
0/cSUXupCJQQv7QRvKsJ2re0Xd9WOdw/CxFpJGvtcIFXRjoSXsuPAibjGwLLeOOzV8fWKUiioUuU
K//iAzloFsqxwD/dPtq9eDzE43TzDTL0RWYDLVWJyBoWKbcDq1HF9NyO/HjhLXMrLzRjh/+rvKap
Uybb/pXK+U6Ghl3iR0/Ohc+jWVSi3nqrUec6FPBnoBX7WI64csLHHfiVuXasvZtlP/qyI44Bi4dg
pJrszn9Am3GnzAzT2ETkph2nX2/ybzU4KR2+oZpgbCxortkJRZKO4ROTsJJybcqSNhAoshJynTpw
5809sdm+WzkL89R0/0aogf6rPNPfS80MN1vvPrVgQMH3xBgOWSF9D+LVcA9ix8BBL0XGZSjmatCd
9pQY/bhfmg4CMsJ1qoCpO7IIE5VCqXN8kj8VaW1aSakRy5eV/h43ds5hBeAHkfeyAIxTONlvaxOu
Lel3OmHe7qwAHV54yqUOoYSwuscZyedVPwAzEBPOxD2Qilx94cWvRB+3ODtaqmn6Gpmsj9Oz8seg
FpUfyp6rOc5HPRCsSbT7piNyAdhIZOYOveZ4unApz1B6LUk6Pq1LrRHyfUbOG7nm6FhTsRywSHwy
GkSMONHYeLoQ1xeL7xZs6/IEw+yGeoJMxPc0ti+yOWCQaeHLxKs2PX60qq0a/wfiTWODmyio2d8Q
UmnpNwYXVCTfhm0dM3DWiRuLtZ/z7q4+KPnhDehh72rVbrDwyVJVPvv/EZz+TRjdmgBaRHLsfSno
H9P0kbZ3SVmuHmti9LpnkdoD14kwjO9b09ZmxrSM/nYQ+KtmpYoUIWDl7Kb3BMMRgI+FLwUXVUMg
ozriu0Mxb/11kFlSTYtV9oEliOwusJwKkfiOGiHwJGGV4aOuYNl+GztKCxkPJaTDWw/JpSFlCw4/
XCgkU3KZEDocPO9ZmQtfx7F0ZYpCaMCpiCU3PT1uYsIuXO0U78muzjVi9tzG0RmRJ3sXOErO8JZJ
TR7NYwoSO07WwkGky+10tcBfFF5yJ4a8QXe2H8qv9dDie4h1UtIb/M4SEDH5LwZ6c5VOHjXW8wSQ
qlH8luHZbCFA48wlKize2/znZTC0RCxv0iqTvwt+oSNlmboZ+r96+CkWsku8DccasmCxJnVOpPMg
7wQGJ24P6n1U+xw9BoTwkvOhknzV/hiOAIWACWgB5FBlLtN5oBV+94jKpYXKqCrsvuJ9uWDLyWTl
eE+MLN8CDJJu5l6dsuwFLdnoWQ1pNEn1uYdgMbTLK5TtifCnNtQxVqDp/YYOYETJPC2NTFxGRS++
NSB3xghJTQWvj5dQnwyNmHLul6Zzt/2Fn5N/Cpsr0RFan3WsN7stL4dIiJ7h4L79ZZqrPlCQH9YR
IYNBiv10XfLzMpxQlHcedyaUVH6hfmJE23u21+t9rfjjV2uYH0zsy63zbDBjRUkBlFy7ZYRAyEVW
LUxLJQvGAbiWKxuea/AeAcepq+M4ESc7Imq9fOBMYFo9+3KSEHuqQOi2aGiISajxDu36VfnpyRho
CX2zKTJo0IgfNNK9r/pDpO8xfxJHsv8W75D5XvntQkl67poM07tu1CBpX0Dcy8HqqusSiIUGUhyh
C1fmQGQEyf3qvMLqgFKgQxQF8JhWNqFOo0WTjDuI1fxBhWXCcePa8WqeT/6P0C3QG4Djir7zGAv+
C+iMinxaJcEYQ69wHO+5P8pppOQOnZY8aOZe17J65o7lsLLrwBSok2sLHTTHt+9QOAq5/oN+oOC6
dGCvQunhgUdyI91TdMJQ+lUOaSID0hY2schla4S8UkP1G7yog+hXlc1k471hwAYbk7uOCgwo9W+s
1JhnbsDANrYFgzV4iKSARiX236zBmYcLLMK5dXN8Shqwi9Qk2nZhcbWmhmsu+evxHSC+E6cayCZ7
6wWTqd/nhSgQO6Y2RHeXiyfxXurljBVMl0lzSowJ52Z0KEXi3y/GKVuye5fzKn2JjSUXYDFL5R3k
w/uJ1Rlbj1+saus2Ri6QuYVo0ovwT4CQ1fmkFo7pa/lub/k6IiEaqRPZvIczDM9kPSE9F+WdAmqb
XPjB1MUaG3w5Pi63f9fhiQ/Cp30ocQO7veaeDu78VIcDXEcCvwAHALRkQnaOtcsPMMpJ7eqDPu5Q
mHR3IhxbwOcu7pqsIurIIblMAVk81jkNg0qMbNtq8+NC6z6NZiTYsLx8ivBFEzzg9+3IQqRrPwbS
sjovckG0JuU1d86mQeHk5m4RCkswQMVR5UwIYtivY68eo5njlpEjMeMlV8PT/Wu2b4/bhu5HJ+Q6
3fIYupna4SRnive9a/knDaHFeZjMIVsPqFhuwIx9MVPgrnJSbZ5V/3fWB8bgIfHmEOn/eJHuT90q
b1G5igXbhovBhFy2xGZcJ7PGUK33ER0eI1NaqL9pgIUyKTbPXlqMu8ctze0CuUZyTl/l2iGUQ/e8
bryMVQBq6ySkWbXiQ87k0NFuet0YAE7CEGcUEY25lOWkiaDkeCzH5iIl5LADFN8J9GPYBgIJDn/b
Lx/zXBAXVNVQ28ey1FZyxtMS92IolHuOb+/3YSTcVlsL7YW2La/NmTEM9L5iBtv+uvGUSlAbf4ze
8KinMmbVjtxwq3TIEtwYpr9TCBbw1g5f1A8ViaphxUSF3D4rOizyNVtPQIBHfhHzv68yuWbDME6P
e51QtJ4IH1AMeKf8GA4sMVBnM56ZFuopsCQpcaWTtlcB4/mgrdELbyodRfkDMd8imAl9v5NRSZGA
YhEQBMvkMD9HpIPv1DramL3K4vwdgDho9Os5w548sDps0IkjYN1IJWm0dUKLZoZjaP6UM2dtKLHd
SPg9vlX/d4rjRsBGel19f/LWhWr1axSr031CPxfH955IGog+hvnRa8xRnmfcHLZm/8u4tSN07yfr
RC5P4gMYc+RiYcpl/gBaMmtVaLaCdys99Ae2OPoh9a4RgOiqcwhEI1Ato4K4JslxjGow92pMgu11
84JbQKZs/u+yO7ZscUohT6cVAwyE/7WmYPlXe69RgApbxCaA+OK5ZBj4jAhGXIjIZL7QEE7MNCcL
wKmBMnRigsrbOC56fxYfjDFT1+Tcl04Ssr01G+VxqNAwPMqb3r3LoA2t7IY8tK9G1DAClGDKPUVm
PZTKA974icEDUOksih39PH/mMCUj5GlpQ1x5+MCRjy5FqvnMfeUYSKpellLyW4Y1Zx1C2a6VKwoU
s9flD158dc6hf5Zvqy3AYPn3fN6xjpE7XWcDLbWq3TbGRwchq7AhJESbEt4hEzNdwsXy5Dzq/FPH
5ZhSmwvdfnDTNDc8d1zoxC9zAjZJTyuUHFfihlGl8wFup5hfqDVgJwW0ckaOEV8sLMteK9rW+17n
0OXQ4e2nnoW8rRphkF163Ydh5ZpSjPU7VHgQ6vEwf5B1cQGrsUJ/bfT2uyX6mV9Bdx9GR6gAYNoc
uOW1HUZtvZuTrqpffG6+5tIrWhk2qmng3W8bOAHcE1ojMuXG71pCUzFZ3rp9Ey0W6tqasT3WwoFZ
D3CS2wiDwIjHwWonn9/2HqfBEkMu7HC7XgUiCExzFwXp2D+uc31aYV1KhlwvaGeISLk+zh6UT+CX
EVUmlzIVCtxbfj+6jNGzUyBxuW7Jw16ma9EpgoF6BNIcz9fMyn4njLZEXOQSqcLMeMN21btmGR2I
RhnlQkW4KZ7cwur9JDRT7GEA5c70Te3ZZW27vA6MmbjcykV9OS+F32UGz0AoMV0m9Xw+kfjsqA+5
G1B9GtesoCtJMwtJ0X+qOHsMp74YJRqiiy8OT54tFdEA3x0vRcuuxG6e+F4TCvMqoaFn6GB53s1j
wFLNtZCHGEolqsjJU955uBUda0AiSPvz2K8MDBOoggiS2W9hkc6uYtN2nHUldfnew+mH2QRpBgia
Xi9ujv2oyP677cyYZtv08kF+MjFsDo/EBwu5zeGgZCcPAdsvNCG1UgfIkO7uX0PYTe5K8Dlg2oQR
wga8ekMc7sXbAml2usGUlC7FKecgli5RW06Tb3rkCY3Bu0UEXEp3XWF/FvOM+BD529ShyxDvOima
X390/MxNwBDVdbrTYkGrx+x5SO+WsqE58wBSBRhCrzCo78TzX7aScDRjapkSkt4DoBYKRekMGhgv
9Erm9t5ySP9ud9ebcKYuygoDtzSzjov1WKPBKMiy12r8SuPR/2r8Ii2oKIwTtjXDxwepiZpO55sU
9mTv7fpGX7cZR81nHzYotZQdbsPE/095YqI3fg6v30i38CglbFFIaTtojRUZZ3PYpc3iEX2pW8HV
m7eCXMQlvo8EkmYAg4GIDfv01ExoQf5yzHhdQTPm65UBJ5nD2ZW/obsGJMCIqwt4zu5rqpGYErKJ
lrXfVtYJ76iJDxb5TqdN0AVogXqV3GkWbkYIIiWcNuHCbWL9uH9AKY459U+/O7ZtBs9chQONIj5y
Vxr/R3YQlYDnluY/5WHMfhfkSwJVObK5177Y2DPKuya1l6QEXQTev1QkD+ZRPiCTShGZIZ1zyXo7
8m3NlSS9O9SLGYimcMSYBvSObgcmSRhJPOoDaxv7b+7GKDWsbPp5SroCWdZyxsANWcIoaBqQkVhj
MxXPln8TiDOUGgKR9dX1nO/r/bVI8swP/7LK+mPztAP+7e8z4FZEXCgo4h7g3t9dn1aYq/eiP+fS
d9/0CTn6YQMI5br4FgB7y7Rdx1jGlGkGWQk/73usutheYAp704e0ciDi+Mzk3CKcnzrAKMajuTz9
yFaUMfvsAlgVJpc4MmSgibs4EM+LJ/uO1pMTreV6RZxBX1/jyNmlXjfyDCK5rgo+ePb3lB3fOeMw
uA8TLle50eYCzFtj8JvWWans/t37/APcdmMjoIk/H6vidwuxJq15knaCiTJlT8bD5Yj81sNwSa2J
Fjl6YMINx/oD2K3++LcN78p9om9WW34EHNGDgLv+x7VUxsmZaPWjzaLDHB7Q3btEs2AybOz9UDY2
UbQMiILRvn14OwXPvc0nBx7JDRw36bF2OqDQwPKCTbvGDsb02pLEwc8sXl7/SuqbsjxrWE6Fv3Jd
XK0BUsDgXBpzrOT4/z7vGCd4/tkfD6dWXep3GUBMPXtBpy6LRyUga+kjVBvkhcTYA81+BFb3vckr
azMKDVeePHkfeCIkLGA3x+z+05yGW5WkUuBdG70un+n0lWkeI1DeXru5GCbUp6MVl4Fmv5r19LjZ
el+ZPw1l2qcKh7HzOrEnL3vlMJSgeT1iFfmd4pDsAgoccUza3DCryVY7KEc4E0PfL49AUToZeFx8
detM2Sz9rI/541PvqKgP2PQt+EwK+kIAU+SaGsgcK16Rtf3BRdc3+7EUaisQKNEIgirohhXiLDd5
P2REJ/NNeecNe98WW+OSVqaqRlg5HQX2/bpxK1QvwBsVAl2N4DeI0Gf5o4bFo0+IuezTCgDrlbu9
T1Xs5v56MnRP/IyBWWccSnC2MQwb98Z98fjkWLatlDmMRVZNDgCm59dte1/z7ncGDWU7GBwNwHb7
tzLxXSrMLLVuDTHRSwS6c7mxcmaH9vpxpGPy1RGZR5rACm9f1xWfd9xg1JnBFehN2c4pzLKgweaN
DZ+4urNzsmsoNJTMEHdD2gnZdSScxExw4GiHrcu1OnJ4TtfctbDeWo9SX3oSIEDkKrC6IaEBmyr0
sV2xd59ibVuDhbzkSfYudsYPPf+aPgB6pWHrlhZLvM1yMq1jnd9H7+lIUraUQ9bXEXh0LSgyZO4E
vA/sg8AuAVTtJiJgYTQQvy8y+Uz5nnpVzeayO2t2JMpj5ce+KU1Q3+z+84ouUAmxDLzFDTU4vdw7
xd6dbbAypdDI8k74ps0O2c+0VTOQjp/CbJjuIYIgSMTjaklhOs3x5GOvaxK90C30QC7+6X5+Ipnn
lci0AW6C4YevY9fk6efftv4cMRtQipEbcTp/fEqZuEQU41sWpgsL5wvc2iGoumU5loxdZJaOhIuz
olDFEQl3gevF0++tP08bKZXBT3UvqQFqctcekNNi8cSpv8OgBusxv5DF0Twjs/JKcZ+V01qnRNCL
81T2/jVsZsNOoUGwOGkEL1OM/KLsVVdQqk0LZ7TSeW/tn1SY6vP8FkG2ADvM71hhfxHcSLiKiSPY
sAuph3hbcpkKc/PpcBSahuTbk3exRv8iuSkLAec1kU9MVgB1gcem5WNFOMkDCwiCmJti3xCJJAQb
gK8HSKre1eTGDQUXsR/WqlX08bn1xaaPzfh+GBpLx7s9lLRi3pA0ywmjcqOeoSsRaswzWcrjeR9m
v4AnLF3G7v49BNZnN1bCny7XwZklyXef742YRbMwoeusEx34R2c9CxxpF1EwlHq2X790naubD5X/
4FP74funeJUf79bDls5oD4UJeEhfxkBhjmkhZrnQ85mq1tmSJS10qoYHxyTUfjqiYDiWhZTkf8FO
5Boy5lr9UBTe132G+i15tPWKVd36fDf597ZOapsBQSnqFpxeZ818EM6Jedsp5tGHXOWgZ5DI5My7
HaiydGlDTpDpxnlZ30zT7lTLvVo1zGcGkl+qkYjpUCphr/ga6e5kAe3VFZ8U5TPR4EuTw4HzuQ8R
wfbnYs95FttC40uHNAEAj0T4w2vMIyKeAFCrIO/Q9FHjDsyHfutt5fHOvTQz32X++NXrz/+CAeHw
Bj7drmaKjb6aZOb5VdvJDQDZGx9Apn0JLY6MbjzRyxxPX1fMT0tys8Apt0Hi4UXVDw3r2j3GmGNE
IEe3G7Xl5zvDz8UiQ9xrsEvvs9G14c2F0Mn3c1j2y2KWFaDIY61KdSIqccGymBNBCru5WxABBnCR
gXF27S5iqACzUQI4SY0x5JIVX4CAN7g2EFAr+qJjAlD78f6S1YkjX22nLF4yh3I7V/3IsbvE40qD
h4uXP5Ukip2tDawn8qwEld0X2VGiXx5/h0zpOFgy/rw0FbhIhuvHPas02ePojVLdWR4vhfO6OgNz
t0+T5Spu5tot88l8y2PBszb0aXsk57wD70b6uuh0hoqcYUgacJXmvU/sbC6yrK+yft9q9LjXjolk
l2DGP/H51pyMw9/Wt8hARy/zY+nKhsoN04tUrU9PrxJMqYMBz21cvw8v4XnbZQsGtITO4Oj98AvA
XpDME/7Ysmfyd0t6R07K3rESdVlI0FHnheHDuYEJImM8oPutjzTlDunKhMJkuvFZJJpcUvbQQxfk
mcvvEd9CmJa2WLsnVX8rSKZMyaP+omD1d7PCGEfrs5Yg7u7skWYlR+jRpcvJpW+3yfkI78Bvk6Wr
CKxmW5CpGPD6RKIEYsmrMmVAW9J1VLd3ahPcXA8bb+tyKR8ja/qwLe0xBi5E1ktc6iPuqjfJ5XBo
MAjLCM4jB9AByoUsOOcZeNQCHIk2hvXzSUTQWUeSrSRqT6LaQ8b750HYz2HQYUN6iXEzTeAONArC
7b95vXSL3hI0Lag/0PrdwUcm7mVia3iYtD/WjQBr7saaHg4eSfGkItPHYCuLvfEFsyjd+ZuH1uH+
7YDMt5Reg8I/LEWB3NnCyllHRbdFrCK/kQHyzEvhlTcQJxao2eewz4DTWNVZzmP8azLiqtHtOhO5
JjVnUkNG4tOOS0dt27NhWbxIYtgvnSjYPvAT9CsqgIKCBCz8KXQ7HXuvbzwfzBozA0JT9TpL0YgF
azwkTSom135u99iwwWMg5xwvBcO9CgIrQnykL/Qk4kYVvUShdftzaT/MvTZmVy/LN0SY+TZR66He
lxGwFcWZebx3B3yOoA1GscaulzVYIRIGyx/Z6p2M0+DyB9lUwJae+EWx2Zxho9NekNg2qEhKJAaq
d77Q5iz9fF/wCRhkeMvQBLiVaydavZqY5BUlneYynWgih97VQvBsDIdTSexsaKu1oDzwNIh58v7E
5vPBf81alOVscUn6yw4N1mgUtzIg3E4mc6er9Il72a+AlHvZeu2yliYp+RPoAO8GDe4S5Ag6UTQL
UNILWcXd8zMjfhBfWqG6KHJsTLv4O4+ZfTnpBF6YWVKNNvmueUeFS7ZuoXBFHwri6tMfNjdpKF+B
sgL84LgAkoxDlsZ8nTZ4gbTTyoiplGI4lOi0+6mp1ZV3LCFxgbffKbUSSP754kXwCy3O1gt3fqcd
J1JOUBmSJ7aOkzSAKCZK0CBLHBosBFwcHlM6EmjHXgSdmqL2EVIyJENiCtAHbt/Js2xsKKMbhHMk
FErZjZdAtofs9WiL7JEQjpDasU5Q2Cg2iF5CTVonFnm0h4DKoODhXT4oGPoEmBoagKl6TqW+nW1y
ifOHklpGp3mwR4AeSEqumfTQkCMykskuDhwAH77dqarFW3sCMVL3ilaGzTjnlOT0L6wdW2ZAiL6d
WEStJofA2DQgGa7GaBc5EoiJFIMc4D2LpufrGMrwkAP/SQN1Pp3XTKdq+axPmn3tdzAAKU1dO3RG
xr7QNDJ3ByrcsOxJWrt5yJquX/2roBACBZKUTKa/XMSXwJmQrrs4V2/orWepWGOqgE/pozEG3Nln
F6as1HuXyi46w4mF4uKndqyylwsT4BTTuZYXaAQtQWqDIFMTK/1Ofgio3xO41+0b6PDyJZjfDsqE
KHj026JTEIwpy718c7J2xxQmjpYSQR8U8/P/36QAB5AvN+BdrEekdsIleiobN/MAoBikja4lTV2Z
+/BTKtt4UiEFPtyDBCr/OpvKHyHsGFYWYlLyVFYHFgkPyHOK/LbzRZGKaGuhUkUfuZrr80vqeqA+
yO382qjYeq2UsycmGjmB/xTSW5vStZYnvikiqeubnlrHswGpGqaFpVmJ2F7zWaGrDdgSlHfnz04c
WbfZXGMhFDs6nwLogvXLf66EeJHR/cb5YcS65B2MNzTOkB9nnPysgllV8ucK/NXJHSji8+ILHZUX
iz4cTk6mTXJwZj044PNFAAWLBqfL0hxQegJhkeLRbUZFzYoyiL0kRXcf7vPSZUIfzy+JPNVKfcHX
QgV9vkxWjMaUIXXFjbKVgyOQjP21xxyG4ORMLjefNwIMyltLpF1kzS8PhtzqSJJwMqpOGG17AV4Z
NRmnZJh3QwOUNxq5GYZREXM9Au6fwqZ3lQlpuBMRNfBuc5OdkTXo6bitnOr/AaBRwZ+JZ8SrLaox
92AdyebIC0Lfkmb2NGDms48VdwdqwKbF+j5Wbyp4Q4Mhat/7Bj1PNOS9P8Q8IksMM2rRzhjXDc4N
pMvd6CyDNgeLfmCliVC4yTkWB7H0ht+ypMxYFi+bYOHxeYjDKRNix8Kr2ofX5qiQVjsjjpXdNklO
/LP3CQPp8tCFgNclbx521mQfUcpgtSLyihKPYlT/PaJmx6JGui5OdC877Gba+l8/2z0mI9XoyYUi
+aUtUbIR9rRqnLdjRfKXjluyAaTTqp4UjrLP4HwzolDHRAiMZI2n4um1Gtozaj/cKdhJGzJ4b0zC
jjhD36gLakqVnIrZwzkQ2t6eawbQhUJgRaLc3Inu8sr5MLJjV8uDw4FFHVuvDc3ffqjmLBcojYUX
cS3pwHEMUhb9FtIdexgoc3Fz4pCbuE+v1oCuFD1CuwLfnzakcog6Cy3aUkFgaDsepf+fejV2LakD
+3u+CVbyLCVq2WsN5bL9t2uHyEQ66A4Jcc0hcRhEdkLMmy8pMWqtubppHHeQvxGKnDKNV7xxEYPc
I4ZfhBnSo9Phk45JLJGOtJULt5oAW99Yl3ESUOcs0OC6JwJ8/17oS0eeBfsq5bgtCw+DQw0qLYM1
QOTy1n4n1e8F+t9TA3rwv8u3ZvBZr/bF3k5InPBanxULG1BXfZvDtQ3N9SmxgYgTTuPUcEoEST7C
IKcwPfe3lmpu5s3qeg9d45uA6KoslimbzSUBc761LZ+2L/SJsv4bin22MJwerKezQCxU2B6N/bBF
hoiqSsVjSaYgHhckMbeMgjnqaSHpjAmFvghibwdk+JbiSJBqBfxBvXspngTuMIcvoZSVZ/vmKO53
TtAqxu87DVpdoMcOMtc3JCfVqHRYUemG6n9/pZTW4ocaAt3klyCoUEaBqox3691szIac9qSb09Gf
YpdvOPUC6HHof6DCR0fHfTy1pUEfcKQM06uviqpby/28M8EIa+oJhVYh479eYiwerIqOq1ik7yVJ
IWtU8Rl9B3yawPRkWhpXmpebjcXOPgU3EapfuT1idxEuuIncYf7XS40yXrXiXVxgCX6JP1tDYcmv
RtSeH6RtoYySp18TiHYQz5h8kg10b+rrN3w7qroNb2Wh+BFEcBU34cc2/h+4TqOgsyCaJIJ0NBsN
VkwUxoB+xNeWJTMwmhxcMqQTe+eWSHDBMsisz1EWRSfnOQkg1jTMYwNKe8PhIfc1RaH+DeWR/uqg
afsBQXMJGfRvkDzK4qaV/CeqdRKALA82004YcahbtiAXDLCUxTRNlnTUCioh3FVi79xGxCdrw5Kz
nWhoylR7BA8iwb6Hy2j/aJ8pX5dEZNT65fEeJM3FA6Xmbfmur7+kZe2a6M1HdUluE+QfDliSydQj
y4UsDxmTf1//h4mBVZjK3BuphuNdj7xaDcDgzUEes6koAtMnhtX9zVIVeYx4/eRL8pnj8v+ROhKZ
z/yziJYj0yypo0gyrjiT7QZKXTFrSqLcwqFJC5Ah/UlgaI/w/nJaWcJy+GsD7gcCuUOYHKV97rdP
ACwnEvAR+q8QuCln10OtkOXtEVwuWWO4mK6Ct52ebJxpJTedVFq1/h/H+/VHxJOhrPBD0s6dC5Wt
MqU1njOs6FZm82MaSkW03VOpYJYKSYLrvOLElHsGNABtAvxODui9A/e0LGcBRVyXECT/oqtEpHpt
f9g2Yllipn3Ud2o6M9jEA/8uXxc0NU6qDcYNutO0PCW4Q3NJMW/T2oX1BRqVRmo4Vp+q3YvOnAmF
YF9+6e8kfhpWGwE7ARBv5MsdV7PWEuM0okMtGo7EzXdfmgzMXFWmy3I0Ma73otZK9qEWalspSSLt
K/Cd00V6QdsUW4uvgcUtMWFUMeqLngNgrIL/kcbCSywqqpgxT3YvxGYY7XPJ4t+VQIp80hVae6Ok
uCxpE9TcwG+0C7YOpOBvwQ/0JPKBCSuqdlfRlptc6pwxg7Qe2Dno5BVrfk1dgE7OJdRUlt1o+5Gq
/qvY5llVMbnyWMvgmlp7gNnul8Q7Y4plCJWwa0Yu7X+fM9jVPSnKRlHOiHxprQ3Z3QazRfKkX0AP
oE5nhnKYB6NpntAC/Apg2uIkwrKexzGcvMnvJvKWON4L5kg84agSDn1cQOk3dz21geNdOmR1FcBh
0ojfbdf5LPKhrQfVOJeAER558c/aCvAQB4eBl7WkcnB3SRE6ehfz2ZS6aXsxHxXfJjaaJZa9qSIX
+1c42PvRFLAhf6l5bKxV2ujBRWZ93PHMqHYZhWppvAo8UKQVytdwL/1lmOPOHqMYKCwsPnQs/Ijo
feYc4D+zKKyfxd2U//eJ4srk8X2L1MY0cS1bMRoljql2keEVzC+AfpuorTQTXAM3YmrxyEBxHKOf
GT25I+Wj9qomHHifBHj8QMOlcAObMPpcVU87XoUOJz5LuufxR7iSGXtAbQ6Gs5xODyBvYx3fgnCh
rqoy9vuCVmmOIU/V0d5yPZM+rWJxpBuUHZHp9HkbpPYmhmPCupYZVXkFa2VPGjD2vU78LrdYVYlv
VSaTRXlaiLx7T9E8db8OzD5dKyOSSPgbiPL2zRWaK/O+u6DYvq2psp0tXQDSggZmWFdXy04tF+LD
CO707LyHJV0+n8y1FgMoUQlsBzIv1BpQe17p1i05TmbUoHNyVrpoYU09hj4OZd2dtMXTw0iSBnN/
NoMrgUVmVVQAt1/QhI54LCllGg+1UWIYTCCpGv2zSEu7eLqsQdH+xETfGucsrOinxp60WMthRKlZ
f8nZCk+BZVBv4H/PP/BtIynHORHe0TlEtVmd6H2/dXINCv8whRIwBXSjrk4XykNgr/dGQ/rbhall
47oUIJKOTl469r9N/xP59h252CiKVKJ2XMMsH73YLzpPy2TRIUzsgz9RG77SevRcRQ+lPV2BH4eC
x3gjjsIaDoFY/Fi6LlLXg+QxFEmozQNBhKRr46cqq1WSKgiB6LgJZH6l/+yAOb3+GG7iQaHEiAV6
KHIo82dAhA7Vhm02Pf1Ad2DHwAmvaz26e/JlnyaNE6CO0gT6JBCcqD+2EJJJA+dSAzaA7u8sENEG
+WKZ/2NriWVSwvALEdmnFkdRkOFd822BuYhNIQCDLgEQAlGgPVUkKJ/9uSUSb2PvSTCR6cre8o8w
y1P+FS3gxzu5OJfmfMte1ccDkyNvlpBq2hgrTVIQePnnIMYBJLqIdFPJPVMpFlIR9BE/ICA6Yi15
7ccyo63EucNKr0ygVDrhvumOjCaZrbzT87SUD0QTem6WhsFH7p/H7y12CieVL3iAAZiR07lx1/3n
nAgVYGQINze3FTcvpoq5qbZLwYk0r6rdg8yt4Ei+520wa4UavI51LySfatIQKDSOkZ2RBS2RR08V
Sy4fbqm4j6ZMz3IZ75gfcXjrCe/NEWdqTedWjjWwDNEj842CQJpODi2/EajpChzbQJqrgqhi23Ec
5Q3l+BgIfMgMMikWejfc96ZSfvmVlhdWixRTCT+qRjZRx9FuWtW/qdlfNH5FdtyoVtyVZe+mSMqs
ekNx/OaHEoQmOuO/TIjffu4z6R4191OTk+3hwhxSceLdGXji0Uzv7xzSxiaOlgqIPeOvTxFcWyJc
tAcuqbv9qemwmOuvRtoY+iUUDr/YgSZrLUUkC5tquCdlDLi8inmNIWeZRtSkacJC9k8nwd+blhoH
GKuidZv+XK5flArf5fwuUiSoyogclN4HsZH67HFeOjvntub2+E4/QgXF6s5kn0AYvqj+RiuFjzm6
CCL76XpLlhJ4R1LTJ+rQNVk2HdKp87Uc44K4j2bhmp2Z+jwVxlYWOTb7LSd7Ixijz5ZtcaAoq1S7
mjBVrUXPEnr9ZIq+Ove42vrcSI0twPfK2Nub8pLyE6IpW4UBfvXAdoxCMo8doUXmDp2GqeegLXhI
wPNTOME2VdKU5tjsQXZ9faWcdT1kGoDAz43RMgqF2Qno3ZGJWi2wIBvAi9pKDpsMKr+OVtn+4UJp
mihN91ERIM+s4+ynAQlDUhdpD8bi68/+eeRpvvX8AfTI2ZfEh5lNI0+f6i+IldfsouBG2OtsPAMo
APp+y8NutMzD49nf88sylRRbADy4G5yOMAWXUDfc4SzdaPMy6N9BbUW4x/yyEJ9u03D/1pi0J+b5
L8ibV63H9bEzaPlSmLJdNGTnAWm3SVDThLNEzLF5dASmXFpilTGCUcullZEoSnHEN8Qxto49wNSZ
B5FFnrhITz9APzNBbXK6bhs2SHRUmxih6J6nE3xK5rqfpg1LpcAiSlc0AGpHgDY3d5vNp32zPNpK
OuAQ4E0CO2SlOf6b7g2fxTHOUkklfJtRZR8IKnWprFGT0NFodBfCBwQI3hRSkTiqNs+qq6fftDwU
Ifho5MVyNbokoJZQq2/5CLI4L5ZNAQtx8k8dkAC5UGz0lK7hyGVPPvubUL30haIeOJBaf50mes1h
uq9vZePuJy47VQzm/wg4vQltCrpEYz9Dwx9hMlGb7DZp7It2X6E8c8waUDW4zVzaMp2wrFo2Q5O4
CPXc+B+bBUKVzPgogECTg6f0YJANSL3y5p5MBRIHoGXVhfe0vROiZyskjVUS0p/+mcARWg/BWYiZ
HLiAOKscsWqfJbOw4H5UnQYPyivc41gMQZA4o69jbskE/BVLWM0pqrzbzUjfKiyTo3kC8Iy8/tIJ
v3LLCXcv5oufSdtq5WGFbV9AebeEH2ovkCEHARX9yR3DAEp76U3engOCVn+KXbKcTzw3dkE3w1B7
WPvyhvQjXTiwnYZc8X0tVaOU8RGe4Oewco0FmS040Vl9QDaxyM78npQaxiCV0iXjV27SYsWyrB2v
5hveUMlUKu4y5KWXLRe2g9on4OHdQ//HHaZGmzmP2UcAPdxsq4z6I4f+clCbGea+Ip+qjoWDqP2C
BKlCKQC8If57KTpuJvMWTlqCVLe/tt4tqc6rcYew0UuXdGAZs0jV4zvRfa2lJHOuv4ZVfo+99mam
azTr0Xcm9ZALwYitHhSXokZvbM73eCBxYVWITNjRvEowGp+fkWfIA+e/s0IP+1eNukZZ7OcX+XFZ
IEp3MYwENVZ/wOXC4EeUd/+qvj0IYYvM6e9QBOaa9Sg41DGFxd5m79CCw3WhWv1/wspb4fimAs6r
pJmKYAloruvwzVANwb+o8IlUHmlGWqAS6ItltTz/6U5r50MvCicktyGSgUlSvS9lZMXSETAvnAkB
GobjGOqaZ6L9/nwv1C8AvyvEoZY4Q6DO88XQXLxSRRnJqsbpzcSE4UPaXqISNobqm+DvsSHs/f+f
drZNTtDbSnqaxGpnLxcZ4IYoxTyVIKhfemXr4Di9lMm4SKVh/XyyCQeQ2URREWeFbDmCZFdoCGuM
9UMRRiiWBhdvIX0xVP1TvytetgwYSsqtWmEmGr4x14iKABfRVuCBbLUWRMJf/QfqpiP3BRa+Zajj
lyFUeX+wJjs4ziK3+No1VOIYH95DM+RjWqhQ3881wd2ePWNQeOW4PIu1hGJ4pcHMT4cPxCOdo9ft
tuQzNz0jw8p5QfJ1QLsYRtE794tbSIBftdK1nCJYUThq4UZGxBAF0IWDlywFOfn136TUxTo7BQHY
ZCptNL3nT4tTBwv4gNwszhc3E3S44Gm0S2A/Rdn3/QA2daeYikOs19yGFghBODK6psScDSv+PdTG
v9ADaD8s4sZD7yDEnegFiBe3HHCTsMXBfEJUiKCYaEF0XlgFdh9mftqH659l0aP1cIZzNMgBvQpX
lnFN2ScNeAlwJGnWrXwDaUlEseMa7X2uo67PLlYbRLGthugbHGxo9wCBSs7yHv6kofo92Ct965hW
1dOpfVDcUyhKbBLvvcVuDqGnkjLHBcWjBD3Mq60LFvdLGF/CA9+nQG1k8yhGpTCdwkqx4ei00YEq
8j+TRf6fB0ApNAnOMoxtL93KojKlIcLIe1H/t+XuFwDJZhfXD5r3QBf70qNx3pCztDd+WttqLDXa
nixFLCL3Dn9j16No4sxDGP48cKkWYJBdFgr96IC1Ioarv348T28+7RZ/tQHxnPDPZa+JUA5xlseG
HGvV8rweae9imOP7iOl6y2FaaPlzuam4N43Kej1k95i0pUuwUqSdb6XFXOgFbtuVypv3rpPF6ZKB
mAXJkVkIOX5RFru+VCy1DEOGcI3MYuqLR1Z+tXmV4vBT+pjPELIbMy1nABTQOzN6sAsnD6CIQEsr
a12ye+lzH5Wnzc8liEUslpxGdemJejwEah8QTau49CJ64G4y/Ni+tv/luSkBOsPeN3aKf6g7fRCz
JDnb7UGiOiTPg9CTM+7+mZ5VsPjcUgQpslIs/1W8iQiwnPlZ+CeVVxjCwvbaHr+l11BpPVOF2G+s
/mSvNC/jzRrgf+sZEe5Cs2iequI45GyIfdSVeHE6Z1JLUMOX7UsBcYnpmeyqgdPTY5YuFSO/gZow
ruDPmibK20j77uPu5n3ZalRw12wQ+yXT5RI5fnhclphJSVy0prYXBhoKLjxti1x+tyOt7xACmziu
/1nygrzV6XHjcjem+xhgXja/fLgr8qLJwTwA0rtprgNbNcTpAQnsGtVmm5FLhoUAqlsszFgGjudX
sr1OmUaqpCdv3yKrGEFRK6aVmscnoTX582GXmXTYPbwQG0TWN2/S6XYVYlIU4OGkhFDSCe6rw9H1
nV0PIN6fFwLM2eYNIljQj+mclhJfU9HhtD23YzbIXQC1p5gQR84dmD3mlVCW0H8hNYQz4lnMXX5p
o3GkshsLp0zhQjRqhvBkBQ8f0fp63ASpOMEwk6ygYx4Tug3UJnDhnWBA+UD4rtLnA+h3PWHscwLE
ytLmdmc5KSWnVkxpiKCJuL8V/qxUfmkxw1BDz5LNSdf/AOmfxJe0lC/1EAUBnKTfWbgasYRwEK/l
/8FQtswGL90fWroI7dwX47GR2Lil8uGsaGzizo9LupusrcOZryOOxlTdkkTywPLEx8KfxxOIE3GB
1Xzgw7PgNz/uYkrD+XDM8okoSEUh9iMfT4MzmV/DJ30CaZcIOFRI7EJxf85U5CsYwvwSvYMC4J4t
fidEvHB/gpL0/i7/rEmtNoxeCKJBuKZknKWKnOmDGSwrlHwTT/Ip9RY/icuG9MwLviOyIkmwic30
OL7qQlge8V2MODLCjwNPgfpT4TcnCTuLCbphAsVU0QlBr1V7B9BXtUc98Uh0kcdazHU0FlqHVrxS
Szubjo4603F2DLSxeXZzVzRlVtiWtp/5hnAKd2c46oxXYt00pJDvIIYGJwkC6HNKrCKuvor39pF8
Yb/jFduFxucRJIB6FK0rb/CnztxNXwyx6DbIQMdi2JC9ntLBeJ3hHeNpKONKsQVJAbQLeRlO609m
6Rfbv5fVrYCTB0I2kAfS+80Nz4ygCZsNAMEmUQ2AewMH25FyPjj8ETKt9qkrDuXgouTOE2dPV7/m
hP46fRz+AK/Uq+PA/HKY0VgP5i1OgaCdykbfRsQy8tJ6CsS2awqquLctBPGOPfROckiWlxKVVW/c
u0S36AQWkOFi9AUyFDAbTvElCsr3hAE2EVGJH438P+VK9qcww337SlhFlfPPDt6T60phX+Bs1tMl
T9tzbTrMFpIGLLrMoDa9C1LWsYYTDqnU7KJiJcbhpY6MTEJYwMAqUtQFlF+LDRYCfpOBxL/+dwXy
dSRmYY06FgsoxeeibgUCRKyUeHa3uTlEx0ApEdWRfgyVDw/wZAdtl0Lbv+mLYKREaCZSj2BBQhGW
UAhINCNYzZDud0/ZOlBzRLJ+74DXQHl13yz384yeS1QFyVtdx+PmdrIZEB/YeBrqVXxsU9yMBIQg
ZDwcN7+5aEBdNsyK9/+BrDYoqKqnWcivzEOG9st2itO4pYvGxZHAkjOWWMUboxp8jPmBQuupcVoG
r2FqiCHKFu9ArAil3s2SwhsGLg3UzkpC+qIPXBA7T6Jnf/THjt5mWPYyfmWhjhMGfsHdQTgEm0tW
Eg7uUQL0yuNzaGBzXFF+eHzWqKwbWpX0RVkPhK2RqiSeKLSXFwjSe7ihD9aqga15OZChBhawWoqi
+t/HkMA18a3hsNYb8kg1s10JHijoAPny7dDzBAGxvmue1BvQ1APMKak9Qqc+P5/MUAf/uZH54MXb
7iQpFF3du1bys2WRF5w2K7w7CP6+0ZWoQ983R2TUBj52aeqki+PUfGiYFqzr7W7p2SNRU7B3d+H9
W2w7AQrCamYnYWUDOrmrfmAxSpUT9AjkeM61CNTETdU7uHBGHwwgvCAGI3zmJuf2a2Lx24nkWnsK
hUutuWqElnjVd01CFlVk7LlcQLYbYiDyk8wDBOhXS3jzKZvXS0XJLOC0CSTAl+VUxVDxHcXVFl5z
lFmp+gUs+OYrt0f6s7s4jRZInZnOWkWZQQyy22Qg1+GarerJzXz8BDveK0Pd8kuhIb9iwRa1zW0R
oiux1btn8iDxtev77fqlzTjgmhAcZq1+zpG1QgFCs8rw0FG8jP3wvNEjb06UxMuwja1m+GOMzrz1
sIp4T7sXZAVv/3zbDMcuzhaosMeM1y+m2tgqnx5o5vrJnnVGApFLbJ6JnMpUde60vx2Nf6D48a0D
mg3G6Na4pbNy4xVuaZOdae4AsLjxHNRD04Nmg9h4Uc2OfVohj68Nkv9ykR1hSnUebaCq1RCZ1kqe
sPPT1F00svmzcBTu3zdRDI1+Lmuym6kFd67Nl+VkKHfy7p9xvZ5en25o2btjxOijXnWkLhJ93RZz
eg+jhHKh8nDdvuByYUUIeS0OwKXTvxku2x357G2CWjuDRRV0k/jvZFi6x39p9c6bcc/M7FnrkSc+
VXe7pDT9inXwg1KDYgCbFuQzadoLS6Tpeziu6RW7hcopUOqWFHRfydBc43QlB2JdGgHcaBAfYIA4
nIVePou+bBqC4g6FTrpE95atNRAaG9/rx9C3tCug27E3n6KN+P2Eo1XA5lAxMLhw+JfxNYH7l2/t
EIv4VsyZmlvzafxi3xOcafuBDW57SVSgjq/n1+Qzi6+C3raCTr9pUyHSWoafhn1C41lcC5bgmOQg
0AbgbhLRyXjD9LMdtCdoLm0WoqAR0hUySXTqBARDHHC7jaWrK9yddD+IIVBCB0NTEuCEKF9GaTff
2dgV+vnMeJsyyqIhXrmVrlnkn/ieG8fMByzqSGohexzULQCrX77Ssxn9CkvrBov6XfPhgYlY2H+x
5wIDkH1uVEllS1tRpdrxoXCkxiAixb6QdLhToNAwcJXqt0OjLdReFTOCMdTYuhFVdT7YEaUwVCTj
KM3j5GGTW7GvLkqaU+lipsxW0JHNd3dC+LfD2hNJDEK3aKE17vOjrN1bRtQnS2rGGSVQ9GzcP3oM
HEoZtUUdtpJInL+4RoM0aGpoid8mGrLXPinmgDhKrhb6gTSocSU1soPxLxjre4N81vj6mNttOxpp
h63dseb/JipZEdkDTi+QpddCYS8w4SGRVpIiQPakUrEUJYv/LaIvrc7/8d4FzzkJlS8hp6DQu+Yi
YRgUSzMMwQ2F71eN+87sPrWATY/UvqNEdF8fWpNcMUKLdPXREDQ0es5s3CXlCFJwqJY9asjuM7So
0YNP0LJpqyaaoSKNETFGWiwmdZ/7lyZeB0/Xy/TLQSv9TvB4YhD7y0z0t0aEkb2TyOLlMRMhDevh
iReFZ37ntuHOit3vd8kEacRkQ+Tu/+pSgJ1D3eIjw85ihrv1I7WkeHRiZbX+XfspjRiPCkR8W1I6
R+9Sw7uLwER/7XjtmTswZiNYeeqzU1uUcr7nC8K8542uYHKoGrDkgBeOkII+mISlZ8IirBa7UKgt
YfvFz1zy4j2MJPoQz+x/xwBlVwbJs7iVpd0hU+ZlNnwZtQJjWpliFi9dgp1tY6agNm9If8P6Uo0y
1Zw6qReMazItTk6hFpS3FzwJuMzdWscw42lg2Oa5mXsp6EvyQC4Zqw10vIHxoNmTpqxXPEXsSwnZ
bcWeZWb3BgEew0gmxbPG5AXoHBh9kHyMkl/sV+RNy+/bNc0WIeHKqYjX3Lgk668QxYUnKhJXde+D
GghTNI3oaH1JstznEyeK0gGDEdeNy9rxtW0esXmHJk1n0OJSf+xexqaasmqiPDy5vaTGNPCRMbuY
UaKBef3oPpGrc5CWTGWNduRsr020ID+UUTBwy136IGm7JgDNOSu+Rn8t7xg97gW0/x7sGcF2oxNZ
XShw7SE59MWdexIKerNXY/Ed4qOjqXB4DDsKPsDfJ0EDyseYVsezelFjhiwc067mRUQxtPnghokY
ykHBw679/i2NrEONR7Qh7KIIZBmXo2kj2giyCtd0XrNgt6WX+GZcYGhXIX453EnQv2Hr6bMphTNj
LtbH/hDFDP9cIjDnwW9C4sxBmhIAVZlGDZTcNWwSngpCeU0xorOeZw//k1QGXQGQr/4KfxSql9Eg
+il+6oaq7qsa8UMAmsLCeUckDMzqkz8XFrGVUNmR0RK8x26j1AB0YIKOg1fHYQ53XLTEErG2YiMd
gDDiTDrLTTGVc4S8BcnUBF7fyxLbdltv5CWkbPFQiAuX9v0odI+LaD4TyX0goyIeXuN5zpPqm1aP
N7xhZmjR15UlSzcA7FCfx9iyyLzJUwkYqx7kxG+NfPpZcQOIWP9tq8sZeEWUiNRNKIdJr8izNwOK
QLPdyMxjcri6GPnTrRLY6fMZT4k+xe+oXjjc+kn7oeLauHbXE7/ZV6kIvq33sB2wkdPQgh62tOlf
o0oVv9Fh0bdEKIyHkDc9nqJ9xjpMaTTAMJkRcxf+bWlH61w2lpRyxXMNLQlmNW649cSgXjxW7zfN
na3U0CV51reiuuAhvY27ZbwVgsi0h0/yQN9yJFDb+zD1YxSzH8eMKPIXDT3gykmhNScdVTxq7WqQ
ZdWyTVEstcHV9YDHR3pLp27R6DTyXId3OQeD66OhU5SSjrPnU9BJrUYYP9o40q7A9CUUdc8w+pVB
2bKkkOJ58IRrSOhZu94kISqfh6J48zckiQg/D7pK6zk468rhwypTFjON8dkHoVPvQkaK5rI14c2f
3h+8YeHboPtZAOOejcdJYuoWHsMIPgMgHP3reGYCl6McAzUZe6P5YGuAB3CNdCdhvLYmW3LVv4kH
k6Ly759EdbgHk0Cd5Fz3n2lmKiOs/PFZbmc83GE/xIoT/fWIDcICaVW81OtxoxwqCrGXTEI4ushc
5o69DiqOyaTAOOtlVwRzgeaQO99NIiGqgAuxoJm8Z0gsoMSECn+TSIg46lCE/w07KWe/a/ChTqGq
7NalUjcVokJ7tP2H2lsWwerMb3ARrppynBTYLsMKA5Nh5TBK/nFLNcrNTJbClygCzTBs5yKbdRoR
rRbcZUIkq2MkVDk0d66ZAJ9nF8GV+5db/PxMlO65SwoCbN9gr93gaAnlQtzmmTp+23CJeOcdRk+O
cxA/8oWrse5McUVMH3hxXYkA130i5P3NYGcKkmOsCpjdE8isLSigbeMfWfld2g1WmjUQCi/HeGDU
BPmA8EihpQG3TdINYnPbGKbTa3/F3Mo0qrObR5hH9vnvQdXlHvSxuPgyWGG2dmfLq6fNnGe6V2Ac
zBZY2K/g6Xocky5VYhCF1v0QGpr4SM8yNBtqLnBfMiZJZi0Ild4ke/FrajndI4bmdJpJEZustJfo
NFzVa6hr2gAostex1YsiwvlJfNzu6cKEbSgYXCRwJdUrzRqUzcbyZBh3aPKf/74Nes45tCjIrQwH
9kzj5Yc/eJi62i34dQ01lUPYC37lHNo6BORfews587g95odCLJAJsqLgqoszuQzQ8xR7ZtUEYA9B
X4fse1nU4YUL+vhHHoKTd9OheLt8GKhw/MN0JLtV1SV/e0qRI6h5USJxnncaIho8eQ5mxIdohl7z
bkG0DFpu50PsxKDdaDYv7eH/HdIpJtpf0h2fbuzxMcNXQBuE+ticEsqoHi48/KkCPZSLImnq1Coz
uR5RXb/I0zHQuQsXbgy4+ZzudLriZdcaAsFWWJ/wzVc3cRrW9RESKgyC3VuBb1uZeZCoxEvZKPAv
hEAMlnIo5nzKC+y7Ili1RcEG1bWpWl5eBRThoNppHbNbWiXKSuToakLilv7dwDZ/MqG0C9iSXdCE
skNE6OUNX5u0wdeSaFoNvUbXgLR+SBQIumri2CdB/Ry9i37XiteioeERDJ7Dq6V+4NoO/TEvwyPm
6kISXd6ShQ5ymdS6M7So5MMVhhDI9QIe5gZi/E1tUZNiqz9vD8gM7VIQujoAj2XKncmN+9HEpggH
CyJLZqakrwjncejhX744LXcGn8qSIsJRYWAzIymb+6Ekyfatfwp4cfKaxEU3FT159TMmEKTv+Gkz
hS/BI9gzL+K5bbaRZDZEdTCnco2JCL6EW3xFzz2vdjIR4DB8dUsMtH0PxOzaBc6IXJTGvmmBlm2h
8AyEW04Rw43jNeFRypU+CNcKf7+9OmGi/Toe/FYhoNLdsmGwo68ZPb2ZMuiJahrHLEGIrPBJ3V4U
Z7ZPS4ahEZjoXGdOgzHw5fKFtjfQC9sUIiOOPEUPlYplHX3oZX8M95vbwjtN6dgu8dkke5fDmNS8
5zksEtLLaAvRvo+McwuXD10ieOUTdQjazX2ycSYhub8GUdp3HL1eJRGrf0e0CkYuN5KMd1L7s9X3
hrExdCL3KCZaAp7ITIpIsQiPW14iwDqLncOQkVrYwgp9newFimyjJwor5olrNLV/4oROyP596aHo
NlE0rWu4afKNEERw2WA+fiyaqbygbUTG1vrjORhb5qWHkNnlqtZkKyp6Bjn1Xhq3zgYbA5K8zvbp
APuKR9SdhGhavorKp7TuSmPgsTvD9w3FUjXJnJRXE4l6ZMPNtI4gGhI0f9aG18jna5FTw6zAcLLX
KMjIahffxRTL+L5Ch0sbOKarhkTIO15lBMODNLx34CeaoMTeaSpDOwtsgt+R1Acg5rm1DpQ4ZI67
pIor5TC2URybXxAuCahHUvaWXnbtbTv6Dt3pyUShaGgHRa1WqAlgY0g8MzYlikfIaMK1qjPCJfgi
s5FoxBRMR32dTJDBknaFC04HqimRoYAGcbzQpyjLfTszAmUBD1K/rhNS/DfB4VUSELPaxBUOln41
vtUZ6uGo3/eyE86Ekdgg+d5zLoMHrsSF6JbI/byPcijxKlcOIG8vo9icnU5pwLFdEfMi2qcVtCRo
zp6l6ozMe0x0R46y2arzE3BwY7v/y4qvsABF2a7UkNH1cA3/LZpvmYXrXk2SFuVGVAI5W7KPGDPI
b7fK5+lW97/YgSoZI1Wct0Pi1D6Qmq59SF0ZR08yx4yZwMKyZRkgPHlPz2aqnPEdhnlZ2Twv3bYv
d544fnSNP4ZQE4xL4qNRBedErs+fDtGoJEGyiUYqcLlW+3Gvpo7s5LWI5mdFabCDa7lyQQWLf3J+
wUVDL9yUGUkhbYUUEWfEUR4nP5dTlHii9aNRC8jyR9CY3j8tSaN8exx9vEu51bNCvMOii3kepL9C
GTuD5VAYJUjpWOescmfHNNzEzpqx4eTY7SREU8xGgswoWcu44zaeptBmt2G7r4qq1M3nZ8Vh4f0l
fti2IZUsojcuwTMwUZsrOlt90BqWyQi7BRpqMHyQ1y2rFJJrXUGp/ipZgEabXILqcy89rOfxGKuv
9I275CXoJRIfgbzYk3qaLRIHA1AsHtn4SVRMgDFz9HoYOe4zT/C45hLqj3DKNLTA5UIkJVHPn27M
0UeLPWFfc5nkc8NJAiGYsMxNGBE2psESZRG0yf36y13U+Oc1OpQg6DPeMs/l90AoAKSKFCn/F8dP
I9aA5AnHT/h7EAxBwS9ZWqdQKBrLmceCkTM5cMgmuvOeBvJAHdiMHfhgXHEm/rancNjZZSkRqTSR
DpLlTOk7t3Wisd+VU6EZJ7tsdNT2Kq+NvUiuM+bLwi+IoNY+/4uDOY+foWWN9SLcSfvukzGX/BN4
GPex56hAUtFiRZAPXYLq/cCPFRMAZh6U0tQgXJ7IDwnOrW3/kpHg2pazO4QNMzDBbGU9dAuv7rDn
QiYc6tsIqiSSsJlP7j14uPXOEtRhJXGI8yzwYJJ7+pj5ORl/7ExxnO/+7hh2bhjCurI9rjrYhYXf
mH6fMNdWexUT6rHGtgLfU64NjtQuTMZuFUqRd+fhAQQeTAPhXz2ro0RgN+vM3jV1KJkTlpsjymSK
jBaD4Dt8XOocPbK0MDMI9r6XMA9mpvrHUCyDZPB8N9sDN4HiMfudZ62e8btZyt3fQgUacj+96A1b
GHJt8BP9UadhctiLxCUHKJ05nBSjRElnwMAxlyQ8kS7hRtZbrbrXoQlHHOjIKifAcu1zqRbXcFHP
E2TkE1TNvkMRmQQDiRKyo3FxcNlp1A1XDPESpLs0+Qih+1svASy8Hqxzdiuc8DzZP+ahQ3hni/LM
2nOE28UMdQrG9A+WKLFj0LTnK0GSoBTh/JuXrgqENKq6jlQW4Bjs3L9CQunbDY6yE/s1O3LAq/Kn
dHdEBaDC1Y5OaBuu78BBePj7MIx+jtQfGDh6I4SbqfasG0p8eMAiMwP0sXC1lKqEoYeb0BBsg68C
YkgTeoLNrBC5WXNxon8y1bGYaQeVcBqqBYwRs5UxXw3MzsUmPa4wvz+++J8Fj4DGwfHY/Wcu+l8/
C+FUOLjhKCWq23L5U1MeRoMxFFx77Mc/IKha3JdjBkz2OrkKPdg14/2KhJi5Ohyn+cjoIg844Wj5
6krFqHXc9Ubzb6zQFWCNx7tv5CwVutpjZGBc/Nb6Gr7MsAaiGI+SSxQqp7OsAKhOeNq5eKEQi17t
jQYY889/+t9vh/4CgGHMy02AMBw4NbRNqreAI/mURozmy03VsgEVYgzSKebxqtk/C+4oBTz6EHZZ
IRVfUyqzpvONABvsNOuci5xnMlr++nxun2lyVoAe5505Q83C+0elNH/6CtzNTIH2Wz1jjmEg/VLa
GDY7f6mvSqjOlHXuJX0Re26MTHxElXeyraH9/bOo1NuAft6SjvyyLQLGnAgBLOjG/Rv6x/I6OzDx
d0oNaiXG4OaUBlPR9jIuE9R3+NIQUQLAADzNRt8JLgeqxlaaYzyNXGNi8o1vpSEku2E15YEBZ5Z8
URd5odcL20pnlNxmNSOoBA2asptK5y25C4eix/bkVxxDd7LqUT8HO5VFIWinuttWHx2c22O9q89B
STLQ9Q1MYcW4xIzh9QpHdKwjdf3GAHBdtW+5ZaGzSnYe1TTgCMrnzPrU3nRTayVn7u0G8JI4I8vQ
17Bx96TAnKIbZAZiw5XiYw5LGNwPUgErtRAMgrZXvFekLVm0AB4jyF164+Ifzg59mpbGpAjvbaUh
dp5mLwqTRY+b0MxPEya/A+oeEU0TLZI5wEFpsy4ZcTC1RvBopcma5n0MZwsZYzu/zr2xl+WYPYcH
n30dHHXpDtrzSB311vfd7i5GxWpdZ/65gKfJLgdUq6V9RAUDjtTzVxVvF3gtXTFNX4Rck93lQpke
uxoeFj7pAWWUkTXKQ/PpQ+YWzTb7lv0xP7hqzGfOwIDeTT3CxctXNkqcH6Q7xXFjCxkC8l1ZfF9m
dhEZZtaHC1cbnoijiLLa5PKrrSVrZ9DysKMW1lOkPMZwB6AKK0HtTVDQ17aH3XAN+DU7xrhl+29n
Retv/RJGfyQqpVRffYm2cvVhCowx32ISTMmNOKpAkQItq8UmZojwimNCnRh6cTTmJT54yJPqeg0w
k5Jm9KQUrgILpW9hIYuL3+iDAb5rV9MkDWoTqKzxoedrCQ35fH6wyQFgRdXZ4wKeNmONVpergHT9
720oDDCBnkK/5T5CLvp7tCogZxEQEIGXL0pv3S7JKF+3/9TVYyUypHqevBRoOTyS0qQt1rtyLYvB
rBubhHKwESlcCd+8i5hBaZ2K322ec0lXhyU0fTojnS20DnXnB7XJV30IRzsypse4lwGez6oFNkMZ
3zFZUHbHYemRhHJT+zSGVHNaJtR0SYJpUVbpL7Rl6Lz4JVm9LtkeokfA7yCLP7F2SUB1EMZw2c23
jIItKpb97auOqHEcKqhy65OWU6QDNhEsCVvxYp2P1qe15yfTh0Cr
`protect end_protected
