-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JDsqEZgrJdIyK67aBySLj3ljEXsCJ4XpecFh2RYnH+wbpZ7HrKGO/apuGVxQLeqyyG0BL6m+QSpN
ZDiRIgzlvw7Eo7L7LmKTJP1SQyIY8FW9VvGXNckHc0F5jR9YiAO9VVoUrnZF1gerh6vLmT2qg72p
MYgJWGiCuGgyFTr1flENTKQ0oRcT2o78yqMlfJvL3Vq8l1OHhfD8DT/uVdzxFsTw9bsWcoqZOZZM
3ZgHxpDRlyz19DsLVSV0NqYx/xSpNWH7WpNETa2EgztuyytDVKYGTVrpLwEfBmBz0bBDBt2eRAGm
bkUR2eUA25bOcRIVvPhsy632okvuP9WUtaSVSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
5Q4uFQqfkNosQgeEj/1/ZVUfka8HFa+/jtDd3Xec4fLeiuseTexPpTeskmdcfe6YuwuKsMHRTdoF
vgS6yO8pfPBdC1cOkcVxAVoIVBuPGJHrHQJRwd6XpzDCmDNB9eInNhRMNz5yxbMrPtYJsTBJ/nZe
1Wobzau5wsN5+wBY4HtBBYMv9/m/w62Zj73jo4orN8jTPCvR0Ya4yW4Qmao8bLAtG7I9kU51INon
PwOVw0pJ3jRaRSRV+J6tVLHufDp4uL7Sg746kD1dJcjqwddPn9f1T9wKA5OMJ4fvzTMmPqZmChF9
KY7K04J9S5rgC+DsbPn31LwCQeNnIOGPkrC9WTJWhugH+LxYmNTj4fNmQCQPMUER3BQ8o9i5eQNo
10f70VzSPwekvMm3ay6GBGv6sWOvYHn8PzSzbuBRv1W0zhFMxkYUKwRHDL0htOxc66b4/uTmoZyV
UkBGnLxckRdHEF7sOViEi6ePw7ytgeFGHew1zKDELwBjGnghhljFo7WColiCwlChDgrUZhaEtA+U
PpxkMt6dUnS9hzPJfOcoT9U/1GNVdDRqued08JwZBAAWL3PJuM/u3/Cg1X28CZgVRGhpG1VowBGt
PJfKRuoypqneeQhYQkPwrc8wQimAQrZ5o92Ud37FUNxGV/5HgTVTa57pK2D0cPuzrHtzGj680+h+
XTet18t6eCOTgZJpfaSniFgOZuoZQkb17KzLdRNOkHpKXQstu174GOs3MdnuIuGhpt1gMnqHzC38
6Yi3ATzecbSoXhbhyP00EoXdy1RJZOByqSnOWxahrJzxWMU/qyh8D25W/qIm1m/BhhpL278Oo/nu
mJVrktcj8ccY4VcYTL4a5zUfwtQchqJ2SpIQoBGWjcfYDwUuPyrGyergBvcGdYeR7GS7DQeNDHzP
d/1fFkC2mKaELbhY/alV7wmKH2bnBqpD1EPws1fCGmQIFqv3QuPulc2KvhWpdBLoD4R3r/Yy+ynX
7NqM423Sfdw733GeWLsBjh8tPvKlurqexvmV71ZZhq1w67z9njtqSQ2tXwFYDVdk2L0LHovGo+0b
84H6TH2lKUMVkVz52AtC8nlnZlslBdwViyoAQNANkcGHHm39ioph8bQObQOflxv+9Rz+Ib4zh6Bt
XoHK26lOVF2sBE6aRRa3B+d/XhOnzsi0FO4lb740Dnovi1Xsx6qEId8L1zD9YRfm8kWlslFsDcaB
afN0G/8g8kyL0bk6nIzC2+EMKmvAx+vTpSmmkB1sJ+WIT/wtyKZgIIDBz+9M77/gGD1EAjZ9hD73
HYSxK/vtnme2/os46OMZhB5yfBfkhI8ltYT8v8+d2jRcZsCAP7jpjoV/8YNlC5/bRHIUb9I9YT41
YiJRRXXPdNYeLkvLTbAgBGCPG6f8xy4vjCstDl6VrAMgP0LAKMleKvk17SfYbOwyFQg1Pwr5IiRz
eYtZCNMCH6QJaLsThHbKN8rZhl2LctBUGFI8DObWPtGCoa04EW34WnPLUCvpWtVV30AtjvkO2iFp
E2FugcZIVyAuFva9AIA81D8+CEr04J3z0CLR01C/Fjb+cc8v7ouM1sGobyRlZJKNbCHLJHWpxwuR
BzpDy0Kk/+zK78/huBeDQWfoPxN/PYt2XFuSgZIzWj1n53q2mMCxa56WH12x/95OzKI/wD52b3le
UOGnV9CcF67AXdNF0ugDiaunydYKU8WRF9ROYbKJhcRR/vqpspXvb0g9uCdKL+6hAeamEascRFd6
F+zlx8Jdct605GIU556zbwmE4hCqwM0JPZDqda1/KdQSHEDHDaN/z7gr1y1TMTuqYG+rgSwG1joa
MixOHYp3sTcw7zhaNaurX37LrhuNxN8XGfjqDJAdnJYsIPYD2KpOnPPynpvsyoq4TLcEr5yP9hQU
zkVrAgjjSIFygxIgCDcYhBLghUl88Ne+q6ELU23iBbMrzlQJGskMwc3zQXz+cfb7cBu1u2zaii8J
rdTSDojH1huk/xPa4HWc/VL546hj0lQgMRnJKbKSXmDJP//wTxmVNKFyTiT+Rjh3J3+JFiPnEh3P
YANcD3KxESW5NKUT1B1YyYXNJhPkryeqj+IcRoft+66ebs0eU3yCWXx6SV9r/C93wPoMHiTcpQKe
0EUw9mJQxbEauJ4Ti3Y+pgZJT2NRe4bWs2jq0xEN7FjMvo4di5CNwAbtMmOcaKqLAdDjWvp0g7eR
eiy+iMaeySJV9DnTTrIvekEIwJihw3qLyoeia9KTwaEaaN8zXMnITzIDL6wJPMYJ2Qpa8U2qSAP4
KvfRvlHnpvblS4/emmGHLedgksBdznStOwirb7qcSyoRaUIjhPgqGa7txwQ+nfwRhGXALyPdLVud
uCXBTKdMhF/0yikkSTrVJW4hT0J7Ie1C8ay+mIT/ocG56ujjoc9OE5yHHYvc9PW9jwEReqDO7cOF
eGHivQm9Lv3BBofTRQgBhmRofHRemzu+OCYqekAlP643/hkrrKnrXdSjkjguTpXc6WtmJw0ROLNi
vhjE8ryGL2Ii95bN3p6Y+zmFYNTp0bZIkgjNswUUsnWIqGpYfnL96w/re0NPjqKrBUHMenurKZMl
LMKH5VjR4Nbs2k/07DCWhT2Zii7eIPtMcigMYYlBvjdwcX7reO4O3rBxzhKkDW12q4zSB5n1bdd8
huy7fztr5nUkK0TLZXpyiJI6Fxq/1iIH2RZv7bPpn6bloS0Eh8IbQ2mEwTi2QUARwn5oNeUiZxVq
kTAPQNlFuNUT+3boEOrjEIGI+dNy14LtaVR4WB/49NRg87zl2l2OOvxX6rRlq7ciVu2Zgp8E0MDm
kQj8ssgNM271E1ra1E+Y55SvRhbbEHabw9yVgFGmTRWARYAHrTMRRkk0wBrR473UcGrNKdgvqVeW
molsF9oJE8uAYGK1bF1xJB+J0VcH2QqSox1vyQUO+hOlxgQ5vUCtp9k+iBXoysrqwsrLVJkEhTRF
1PXDzoLPRY/+i7UlRY6lQy2bjQxLcp3m98e00HQsCWsiC8ZUbWCxFNEXf7QTKz5AV0P+Q7wi3bSw
B89ypiYBLw4X4oGo8qWBS8AH+B6XcgwHUip8vz9fmNf2+3ahxEWyJBb8xyS5TJPNlToMiOu670af
g4hwDdTFC149WJZEpS1ooaez7J2XOm9tm5b0NST2vBVd9MMO8GPjRDCqPN5bQx5RZItmk/YEFmLd
kGhdLGNRAhnUh0WApz+6gNJKThSmwNtxZ5mgG8a/bkcrDH0upkdfzqo9gopsoSFGzGtSpB54IoiX
zx/PjGvh6UXJevx0QYVMmXPNgl+RlxZaRpEcodaeuS9PJH0vk9VutV3di++mn8DJP60Y5HtatK3X
aoY2hnInlm5PXxxonP2K0Ol81sbHSmc7Eox1yQqBlcoBZTQoof5iuppqATkL6y7JUmYhYZAkDCBN
Cf1WQISkYFWaW3SFTVMLZymZZqEZUdrbGPjsKahhDs40nglb3Nh9Y/2iMYf2wUzyhyg6jgBcBgkj
lEE34SZxg0Jy3PgvkrmK6+JTV7sKykccb25lUMIECeOND66F8hx8/y+ZWPCsKLy3nQ1huggTV2+K
1bHBm/43DDVcx3Y1GhSeVnxFCfGZOetpqRa3tmgrD5yqzUROQnjFo/0ntpbzl6XO2vQwFdEuG8f9
S4SJUmGH97I7nmmI9rmrRlhv1aSgSjOcGKEVH7h+2kj4PU1J6sVoDVh/ByLbw9GxqTV8OBZGx+eq
vzwafUa4m7itaFUnzwOh3Tf0d+Ug6q8SCXR90JYz9e69ymd1PnvEV9rO1S4PDHpBn2WvWHfyxaN8
HP3GTJb95t0iJVQ7IInoKAmabzTOSjvpTDobNNOlCU6TZ29iBgrMkHZIa5Bptg8LmQPj9e1d9iSU
LPlG9Mda3iZulCSkOL5XOxxOjaH4ojdbEn1aSUZY3M5jMzs2fRFGHPWcuWzc66yLMge+Gyc7KD2t
GPhI+6UJRPyOdAva5cjsqIREqcRKn1zsJl8potxBWoNLWzfIDBu+V83h+AWbj2EKqgsgbeNINjAf
7IqzxCyAuGMJVuXHTQbdO7iywExVt5cGoiJwfNZEvCysyKpuJsE7ETQB2UykdKoS3pUSkmJj+hSF
Vdjr10CcesFZZxOc0qfg2VN3dFHWPWmoi1xLZ9HI0cD8+Koc2T+DOyAyfLoyXxCPGjx7iRXhwnj5
lpeFn4AnE5DcdhfiGg9Z/9srqFbW0S8DCdrQOwFve2dKYJsI/Z1O/jIkJrKIxAEuCrFRof68Gl2+
bA6o5/PPNTgC+UEN9oryMcCSS0TJT7m0ozY64BIFXJ5VtFC/wpvXWPlGnkfeAQ3fmmjeAQXD44gw
2Q+kjDBvEv7gsWioUI3vuv9q1IGyM9FPJ529pn2cu6RBOoBGV2yoYOQ9ClXbNX+EGNeli9fl9Qkm
6AZA9caV4hzXbApe537Ab5gfi415DEHd5QGV5bV8TssmUoFJG5mJeYPGT+zLQzvYH/vECTCEHxg1
ulK0gHLBOnQ8dWX3HxWOuUejQAKVvAlePvacItQ3eF11C1CUCdU5IH/uNYgYem+UjmGn3cW8bYJd
bR2dWeMb6mrHmGdp0ILt02M5TItOYgJtTGQSp8NTdFmgiWKmW+Ly1TpsdbPFKlDaxx4ALEbum3nl
9KEw5qE0S97V7OfEfqvNwvHP6FmGNJlZdu1GscOKyVBVd2E9f7rCCZnndcIkx0A9dTNNzp/Kw5z7
ZY4P+MyW0JczpDVBs43Mh8IJRzJr4x2DPkNbbzLrljuCNDQs8D2lAA6MAx8ncxjCAP220ymY84qD
eKH8au7h5zeZr5hqfCo6L25KilzM+Z4q0OwCj3m/Y7Xk1Tqa2GiT3tiaM5CL4ZtUENX8tbi61yFi
xEmRqcD29DydH3RGWRZSPL48lt6XXkZ0JsiN/EgzN7BPs66CJNPPO1tjlvvCdpRJxDS9mNr9L6lE
AdTx+fw9X+D0ez/xL049tPS4cJRFctF998rRFjOzWSAf2XnExqY1wIOQVRN540wCKB9yVMmHbULX
joerTzhwAZODuf28VJcCr+P8dcA+6gyAp4Gajf5uulvItsGjmNpB0zXuY5OafUjA4uws9kJKgoHk
klOC0hYdqV0axOBh5tPQAFMgdimWnuelDpIU+eG+E6aA96GUBBXio+NAy2rqqiKWVl2YpNCz/8jQ
FKCi/9/9I4nelM2akMAtyZI8NLtsxmzb1+Skq2qtkWaYQZCAIpRwrrbrDQPdELKncIwKYpwzAMYZ
r8hGRuqsQW3QaFDy5/h5ECZnIiyciUYF5rSkmfH8HRlZmJ5T6jWVueZtJqvHDilcZUeJpC7TNGoS
PnRhlAgoCIxSweHqKFjkdwR82pHnMB1hNVFTd/n0UplPuJlQciJxU3uJhrZHPY5p9PErUTl3furB
9rvT8krycea96Pn6qtKH91cfnUuYEpv291XZkjV+59DfNfMjLLUd69KPgi8f/vFv9EDAE7nq/E0G
b7o/xPbohLwJ2KPrJhrpMuo0w9MagDZ9r2WyZLi5hOdNXUv5q0ZotUYKkuYjQJzZfMWD7bLt1EY1
TTqP/gLIrBGGjBoYURagVv9k3rk2ucYzr3soECvarRXN1Ds6muJhEJ1gb9JwLOCtkBDON4YhESLu
Qihrz8rnDAbjD9FcDCO04aSFv9VkoHeM24B/4hwySOJP3CTcVGPo3OZ0cJZDwkyfzWL0QHUZwihU
4mVbGVCZu3ZV42yzYZYsfvB6YbA8r0NGr2NgeQWsOiVf3DQp0dGxEbZbYRy09yWKtffY/QlX4dMu
H1FJT87Ctbm6sPBlEaCmO2A8ibvvwpxWl6G6dWcKvo6oJMq5og50tCCMYZUSgiF/1rRkBkKcywGt
W6ww1B10BXkwVyctJX3LmxzZes0vG7SKHwWexRwfUJnd2pxWhpusbM4PK40ft7PUUcA+OieL1V/c
98M8oVYpb9qcCz2h0dZQnhAEA4O5CYtbzX/OLJp1uPBtXUPIHy4ofmv75Lo9lgdZ8mc4otdtG0Ls
0eR1lnCfS4POqNM/jKk80LkFooO/RHw2PfKoDUSExPuvJ11KohduPggxmTpnOP5vJRiorcUSGTyd
Y2oP7IuVoJU6Q0EqE9ZS0UHurHzW4qPtcqY9F1wJiLPdFz28r94gCaR/m9AOt4lJIhZDwYfNBJSe
0znmpX3I4KAwh8yiV7N4dY9rFtqtUZhffxmzp4UhdDbAO0cl+g2Tkpk7WV1fUN10MQKwYUUYa25q
aADINMmohmfsHDqtYovQ8WowjQYLKhZ6XqQg8+BoQ9CSiOmPHKpVd34HsZC1apjH5BzvluQxSOV8
8AiPFyphzOlTGUSOdn756kx+r4ChFrlYLedE4+s/5FiXrO9IRxD7LA+9MFGEYg+iyJ0/TcZrNA1s
CEKHlRUvOV8WAe7HAgDqNus37izx4jFYxp3jdfMYsqMrAaZUM1L9hUHmn+LRcg6Fcb7L4GS0y5Ek
wAVMokG6MNQdj433W/R3IvG92XOmOgcvqFQ5j3QyBlgepE1rt0IkHRVq8wFxDbXSbjIe7LUvgzrB
9M1pOUPgRZA3FgL3XjMFUdx0Xh3LPZaDPdjqQ4Ycuk55aIv4w9kqs5NXbH2kIYykBt6ymbJA4uca
fc3GKHHQ5gus8TccDW5bdoAtpXPFETglOl5ZKhJePiAa12JNkNjruw8i3vg5VE1/bt07VuAS9vW6
0tmQjsM3xJRk0KEz+Qn6FLG9mu3JxvGdkhWyW0i726lOEtN9s7fBbOEX7qMJZtfbeTMPhYiaGjeT
UnhCLMdVdhTmHfFxOM3N8SRpJlisocQXTZ73xdNIQm9kpBcUQrpGgXzK9imHYQurzTNfG/W8nqcz
hG2bj+JIxjna4lIvvICr5GNHiTeB1GBZWOZfWIWJN0aKqaKK1MK8ChBpkruNbK2hpmyOfNZ+cmGc
v3U4anHNmDvXD4PlGgW4Rg6RG2CTxh4n5DDG6k5ZSbMDZ6vO2fa8XxvMQEI4D5060uQvFqFv/HMK
hz2vkMFR7Gv/bJnwSDdPHq6/DmE2C2y2SbMlwIwwZyflFrP0yk/HEBNYCRtHa0TgRZgOjB3ylcB4
1BuTHfFlo8OliqU/Z9czWNwWroLBbg5wpmmzQwtbgRkPZxqG66EUqcKlXTu+YCtIxENGJcBWtWbu
W/rcm31LtxCwob8X9N6IzFMtig3wR+3ZP/2aIGig7vnC1pnKhXhF7WTaccB6Ss6XfnDz2DTjGiS1
zg0Gyaw2jbZczBLF1tel4Qa01ckPL/JEJ3n8svjAu07vL76Vtdx+XRj2du7/wpSfvexVSF82KpMw
rCDbbQCQdKRNRz+IfUcLWrx9+MfY6iCcQloZl+9BIlbs13+xGNda1lUjUnnn0ObIh0uB3l8xE/Ri
Buc9FSApDpaMNRZTfD2xruRzHey9LG/2I5P7a0LxjfxheEBRWYOaLvUMkvP3lHVX/NCJj0o0FjV/
aawHXx8ITeKJMAL9U4p3P5zpa1ewqDH4fGIc15onJjrry4hctGud5ffiApXvwguE/o5YrlsguzO+
JWCoevZ9BcQS/EFEisuBANLP56BCp6jRYuy2nvLgfBg8ENavpo2wuDSzgfTeOSdy9RIsRmBLlJy6
o0UEYWxUmOLY16cycOViwKA/I57g8nerKTE0NVr21xGoN9UiyHZQ8iggqq2Avx/UnZRvdxyxje4u
mJkZhBq3m3aE+8TrMEumbTEyiUDI9BR9Y9RGXdtN3ud+xsKv854TFMYrlhkLOsn7bDkp5g8d77u/
575VC9nWClURE+de7l5XfplgfT5ws+ELlrHdZeiwO2SoL8hop09JS/f7RrIjgmwFV8hXV6n7waUl
I+hefZKCv4dPW/qUcmP9svlNutG5cllHJy6FrkV4l2qTKRVG9JL7qvqBShfHZIz3+4XLWKnWrYYa
X3HPetsV2V5HKoWkVl5+OcPIwqCoV9ruLrsNUQuxqymrGNHVEGIvRssJHQtu4F0XzW3IYJBjgy+Y
vwiPsWCte5BX8Ntp2czW9HnbMx11oL83bjDA5QHmkL1322FPr4eRcQu8HDuyIU44wM/28yVvfJRa
BPM3V/vlgh6u8XvznL/bS16LobnEablc1yQuu06/ashrzH7VeRm6qPepHKeEjl1X2aIusk1nzXse
XRGeHWpRNaHEK02x7Bib4RJzzLHybGInpBGlJDz5LroY+2YQjs4PLz9spPyhzVmN4qnMoWdPwtFH
2FxHG7RScw7QOz4jyUihJEgvjOgc/DF31Uof9Mt4neE88LB+66yNsioudfa7MPzYKcM8hF5rUUCl
J8+q47ohbPio79XJIfMS5QTCEaCxYUmHoikDFtfuJC7DsxdcbT3Nq0k01I7U0NhlguBsVrnlO1TK
u4h4NLPVTGDAH6HRtVon3qtVZa4d9XwINk1jzIB34+UwM0/l/dxSrsTpdYwbFe+hUvMabEU6jNqf
oyqCNCwghI7UrMgUoxBkqevVLtWzlVaAeQRy7nwwQtFgJp216pWiikqMvmx2GPn/G0QwjJJjKyI3
4HesnA2EDQAN+uwxA4lH6tIGwuhAdel8tvwa3Q0r/wF16ZEzKUb1UD6B96aYpx5ZiclWgLy9H4ff
dH6T5iOxYVle5+ZI1y9juj/BVG7DTEzBFjplRKw34/GWFN1Bg+jG25VKsKJ2pYP55XrIsXN/TAf9
afaXjsjtMtjd/AEM3Jn8vy1GnJDRfbOrRrXvdajiEWeQTQbZzs2H5KO9xBII5ppyo5PKGg31h2we
hlSNBE5fzwhKQ2Bf0uX1zZjkU6iB+3dAQq7x/N9MGm7BuzSiMggkmRxg4BS841MZ2TIXmiQ1AbpG
V8J1EuvQcnE6MOpWxQlK7IiU8Z31mY3+1YsrE4eXXr/vzQaC+v8i3k8mA5k5sPxTILf8aNypzMhY
2FCC5eZLK2535TQAqHDc2+JmUKDMw/jncXonZ29wPqN0T/c+9FGp8r3GQ9pqOKcpnlueewy3E9fN
OAQmBG+fQAdtO8ZWWCDiYfocQdeTRTRZDabbHMB50/Tx4xv93X5BDyo+OdIV02dbjLUBQgkjVfAK
nOX8a5J7y5dEI0/d+PdPR6xuRTEWkh8AC7tl16UfJZi0TisGDWdMauIhMvXGgwmM9JMijOvWNpfx
b52b5eJlsuBxTqEW0MRCEk9Smjog9G9Jk6XNhLlINVBlriJH+UURLoD9XgOMD+hRqvEi5KsLtJoy
IbzuKVBfk/XZAn5uduCltwD0nD6yjRTsZ9gAFHA2B7TNmdY9t9ReYlFdH36ad5xlP+Zx4TvyFMXD
W1cvaMaO85kEsbiYLLhmt5Vjp90MDTZR3iZO5IMHUkzPBdIgvo/RkFA8fDIuCQqHjMMXqTeF86rx
LbY2U4qREalIy8z3mndacR+dFsxcSkJm4qfc06ufuumn6Dj6c7Hz7OunRL9XYmTgk7CGICsUJPyr
9cwcUz8yUQW6MAMhTPf4SjHobhoepZ/yIQ3vyhOPD1g+iXzJ8NquqhxgGFDdmNUsTJefLzl40ysY
SY7GgqPJ0+FPe9V7RJc9Sq4Hq8AxEaWqgPIGnSokBGhzHdj6mqCGD2tkFYuLFYawjfOFFrd4qSjW
O+b21wlbtxW+PPRpYoiYbuxbKrfxyk/JM6dqArBKV7UJNSuGGsEALy7gIfGsEWGrLm7TigbkQ5pU
4KQQPmhSfY+IHobs690v8mk2ZCYUEbiba54Q/5O/+sm/2qZc7ehOccid1oohAx6EOKCXTqFFvgTZ
BxnVkJpltocBpZgs070G6A2cEmXRsm3J/p07YNNOjHe0mRmc40RvrFf4YZM4OO+LKWDgdcE240+d
Lz4axK5Ti9gn3t9j9h/ajyUfCEtjcqCWoIYSWoNPH1DQsgVfmdqfCDdSoVCCr19M4C2zo1Vm9I/T
6VBFDchTge/97ZjjX6QkTHxxhd5ie4sWZIw9Xsa8DpAB25UhtxP6iesF1tFztGvFWMyVAMQz+aiE
iic26yrADxqDeLzyNeznGHb2eqzioDEvAfusgb0mAmX7yiUO9MONLyR2QNFTsJn8gq6s/QiO6imD
rdUqGs7gCJA0pq2JU1GVN8ODKppd8iU51op31AL50pFXN6XKz3gx3d2qEkerg/2yn0X6fZPEmHIZ
gYK+WPw1q9+mfZOr8AFXLTnsFA7US47sqyhDUJAY+xFm/Bho/84SRlOj81oVQASyzr+oOxGz6ZhG
pkzU9nw63p9iqi3GuQV5AQgT0HEAFcDuliF+SN0Wn+OR2bFYfwMa0HxqTpyUqqm+UYZ715GKg0JW
I8GPsYh4KbUX7nZ63x5QSwPK/WklfpgeOME52+0kLnNZ7Wbxt4CacmNmyd4wSD7zLoT5EDvWvqEp
mwwp9LR/DCVBlD/nrGP8LmkfWeZFASD+3N7WrfnLrshNQiYOp7y3zn5avq069bVE3urde59aqulN
3+fqgGWiHN1tmuoC3v47qCpDvzC8ktTpkkrpvUi4gdoTr8hJ9ZZnuOdat0EUBtUlr8IEhBCSBeNq
jxgjhoITsR0tsXsTohUyZNpXl15BLKwRM5gwpxiUNzHty6X7f5xpUx9HMuW16GtbekEEO8i4Qznm
MIZKp/HgDOYuAk/ekx5Su1SO8IIYz7qZ5+6DBPoAEJsAvxEk74MphTYNBU7Lt/YkGcWbyCMqnyxg
Vg8tr9cv/oyQk/UiTP33xlYFxFtYPRTNO8fm/70tTwf7MUYLZXRRq8SYOZU1OQafL12Z6JwahUU3
1bWXJhFmuHgRhMO6ccUr0fqpBApTQPVkkWO5MF14Hos/0+T072yyxU2FcvPV7l+hBUi2Jr1uwbto
t1gV6yCpM+BTVCWBsKsHBoj4sn1aL+jomJa1lWeZ0G3OlsukMYmLEvLvB90rXg1CiluCt0kCB7nc
eOF5kkAoqYzvDmXrrm/sK5T+/EiDfySA3//HaF8Cvwyff/TWSN2aVm2ItSh4gm5CbW5GcZmpgZXU
WOTxiuQVeivSgXQI1zKXibfwrmVYX9BxmSIrjtqpf6jeduhfkN4tIzz4pmKouzmLfFYYSrORfGNl
qzclaHIgjQNGfUGUTQfSzcin6xMouVnmGAwty653oTsm8jd1WvrKmHZOR8gntdTHg1jU5rv/qvP7
RSZ6uj6gU+lcnpGuMNF0woKXlDkNwKWHqwV2B9HbC2nIdqiz3aCQWfuMZJ9avC7CmfWTCOE1d4HQ
WjFRmsygu9XRpnsSRXjRrt/5k14CK2bJ5OUltRF91cRakg6d0N8mp/xBzOv9CIX0COTSK42VoeP+
yipGAEy3ARXOjFb1TMOUE3sXO0AH1EUwoav4Y1A7dqDN027MI4H3TFj+A588y0tKMylFNCtFiuiH
P4U2+I63cvJjS8McC+td69Y7X5WkpbBp4z6lyVokv9yUC4z9oKr1k3EOQjQPvOjGw40JuxigLqqH
n/OXY7/MX2mikZb3NWNlFdx6m7yLOKpeZLHotF9YI+rHSDh/G/sNm/vSwDuLT4y3RVK9ew55u9Zj
nUp5NObDuZ9c80y/9azNiN3rScezDC6D3uEClLXI3cWbCZfWjUApLrfq5ahG5j0GwmHUs0MKzm8H
vv3hD5CFoDZN+CwSQPfFSMHcY+FKHEamLem2VBCr2J6ZANdArgClrsIwAtXHB8sLlS3lRrAEpZEU
RAbFbLG6tm7b5krP46NAKMIKpXuO25rzAVwcI7qH3QQjYTIXt7H3qOL1P67L2aQ901NCoZsuIetf
AC/2v0cDBHhuQdWMICl4FRM163UrsBkHBuu7/EfMIARmIR3n0x76auBjhrs+gTws+F8UQl+p4/sO
DCzovf31aiIa4MZAVjRdbkhPso8/kYMm84UjapO7opqDRnCTDclkR+k6+57ONjGfIdz6Rwhe5YfZ
ihRzfEQCNxe3L3s+hdHJ+FnrWhI4bESGHuX5k5gBya71FMlzT77FnllFBs6SNFjNj2BpMzirdr4/
0o5FQToIC/ZEwUnvzZySrDKBwOMBfpsDqFYOh36lLqXoQ/MGCJiqZVvxcZ3/HdnGHL2B2rwVdPhH
pJ1fTr8PbMvCyF9RehAsoS06KVpLoUY+jAMpTvLXKtDHMe+1xge7GDcBlUUdO2vl+9KpG3Oi9l8i
6xPgKG4kQenHY9P4T5mveAetRuOq/mdnsZGF+GW3gjDyqdPekV33yRpoCNIl/tDtbEc7K8F1Q7zU
0EVRyiL0mv+/crlr7xIFCPYm8yK0PpNNUpf3gqY7fVlopNqQHhoNbMx2fXC79rjDxAAzqHYwc4az
Crg4rhhvRd60uXyC9vc+wVGIRQWfVKs0/woizA2jRbUzQt16ct1W2EE/9CfscUZboAvaVpbQSJkw
OCb5dInSNlpeQGOYDq31WGUlJ4uwSvJhqtGCEx599OgKZYqAGpoqbOmy82Sx85X5OwhQvLG/W736
m8h7ENglvMUtaY/rgOjop2KbMQrf5WNuDdnKY5yniWokrKC/CBKq6L4hhhIqnbs65X3BNqmqOuHH
TEWstbTJR9bkuh5cQb1bOSWMXrjct7nqXwrgIUyYyR/W397aNMleSahKkVG5M97dJYst5AYTvSCa
g5r8WuqJ99mwjTYndaoQHqGA3H65QncRrJlZWHrR7iU74KdUViqi2VExvsm+PZLvjAyIslNUJ7hr
2vCqP594CqPPd6Bs9SVxf9xPklnzbLdce1Hwb2g2vp4IBFa4BblD12mvIwkJDaAKbb+7G4RRqXxw
4PAtpvlf2gtAGZmM9zMCYYF7H9HGKafY3Y0jtgi9R78eUcBlop2D7RhUpYu/g6UUaCxGqa475y/r
3n4T60XXKQ6LTD4w/d1flhe6RNCVlPPoOuPr973EKa4oC2l/J542XkN1TzrLVaz12E7/vA5B72Uk
JexUTn1dAj+D+usm7LA2o07zJdkefTizzXjPSFDqebD2YwfNDOh/mBZQKvyRvKKC3KrHwXgF7PXX
so2uXCPE7mUH2pPUYTUR9ThnLYuqa02YhNqwi4EBbBxg6+6q1957XE4Xeqx4JIs2QJAkOvp+JoVN
zvMFZq+E8kxcaotp9i2o4MxG3j+A+4olAhrKTlhqyNMNyOww+mTZmL2yBMQXCPWg3JRuOXhRR53e
JcwarZrsZFlozcCoDqePREgchwYZPOQ4vHQnObblP6Ytmbt8Oi5P6oj8Angb7wSPXxqNxz9MLb+j
vZFOtMAA44c6tNmih0k9VN6exzX7GnKx+Ixkj5pkqk2PygDF4bZamRY2DXL58Y5gg/z/C3Mav8jQ
02tIu0G5T45vGpuj6botHVZd9H6idSRaNkkGb1XE45EIY8MRQjqx0NVyzAtvTigZgwEf1WGrRWrU
XKMBSnOKtghne5kFC1+fQjXL3Am+kB+M0Apk/8sUZdVbyDt8oO6unHeJSHT8M3PPFzVx6xGFTK4U
kj+HT090PnI97rTdvQpjmLGZcfJ3PQh81VFyHb4ZN78MOG6LTNfBJfZSCzF8fGf73vMkhbPiuZQ5
b7SS8RPl5+YQ4alZkVQwpZd5mkKGqtVsJNQwcY10uZ03l5HcJIDivCtE6u8+vQACdnzvp70rQwOd
fnQPHXooW3V4kn+rajSkku/alM3N1q9eQIWvXtoM5L62SQWSLI3dha71ASbSwCjFZN71HGkY3Cyp
AUpBE8nVf5D7diQW2R+OFtSaJDF4aRMgWC58t432MLHkA+S43guanVmamcrv24rxWcd0DuMQaMfy
SUouo19lFsivS6J5sn3RVFFh6X120S8zSYxKvDBKU4J64X7W1rWO2NtOzWNCtiipSdBhwMUmIfTm
FsRhr6JZtdR/eaMumiBqV6gCq7hnFdtsj270jy3359yzXf4akyDIFSgFiYgv67FX2UrS5HzksUfl
x6kYpPedlnzOv+HoNZMoS2JN/faP0Zk/NyRmGTnqx4B5sz52/iB8CgTXBgFd8qNzX/eTCxQpno2L
+N8/sZK+ldl8pH1DIZYuJtXrwBJpCyN5lRgul56ytufPb5H27BKMS/uonyZFEW1gK+tvyb7vSbGW
ASHJM4Do3vV9ohNocSeAXMBGLoqSVE8tKt+L5DrbOEYwtvwHujEGeCWXKa9yHIw89FHsLkQchYv6
1SKKpFn3MBR8XPG9bVOzP6VlLfDWLMNwd/Z++OUvTMzA5SIeeyinI05k9MDxyZGS3Ae7tWj3J4Eg
P0UQ5D7k
`protect end_protected
