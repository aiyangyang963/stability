-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UaTqydtiW/iV2b0UceidymHImZOrJETiN6Xfp2B0l89lmRDkQX0FmTKmwkXLNdOviyXDknVBQgJ/
3BCIQuOcoGdkXlblVzWt4M0JKo6x4+4aQZnR0+oNTu0PbulYlELX0PKwZ4e6eR6Z1EkbWEZEOBF6
IriGeD+mUPjGH9EKX52cEUjE/ncWTJnceN+hm3UU4I5ISmzRsp91VUHHL2MLrwkPklFPRW8JiJ2E
3uE7UgaiphSzyVwSLekcwLJwHLt7qq5GFc38QUqOWTcb9hgdczgFlhbPVQZu8WW74eSfWxI3cKwc
qEWn8GuwZJYu9TORVw1LjxO1snLcaF9omGHlFQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
RgwnOeD7p4GVJ82z0g4xaY0GAYU/zECtV4pUWtwNn08/CGYqO/BkAef1L24/8kxZe3V4QAhMy1qL
XYYFVs0Uz+Ycs3cZS5k8r21N14a5Q5wdTVdqU5qPdMBI7h7uRuS7VJ/XYfMT5CqnVAtMGGG0kbQG
swGfyjnkMgU/aXA/Xn6QVkg+h+7OZ6UgcTHdXSzRwyOsZ5ou0P6ENt+xy0MjFW6vCPdwuQjvSgKb
S1mbwH+H0XbpFd4G1poOltpQZlacfaTTek17+coPwJXgCBysUjOHYl6Gd2LsD+rVeITgF13lCLYL
zQYI0vtwSaKH4n7gCQ7Ds4PLAN+x6WKX442LuuReYiEcE1oVOMHU/y7iFAy67qrkCw6dHfckYuBv
IrkzlVyeJKofoFKMj6ncG+D0gyYWtsaLrsCdNAj8j/e19Ze2xa5SfetkFeI/dvnD7KPchd1hu3By
EwaYFPNmXZAEJQM9ACBCg0km1Ndnykeqs5xbHjD1G21mWugP6fn5wCQPA+ZtXTJ6Js/jfGMDENT1
vHlgQGmAcsP5LYuK3ZCklrdQoZVYqllofaP/R3Feua/0p4hIGPzRpPCxTXxa0l0Y/H6IIusqcmJj
MzvSI/ss1o5kNTCBmKwrDWU882yDsGJLwVpciovqoY1KjKp7CPGu6b4KlnNoZ+K/isVpDteFZ2UC
NU1o8lx6kjhavvNG8vXSwoBKdNrd+Ehf1teD6AmvXQG7hiQ4TwH5/HbZHztA0kdfwVXk8VfgaB1D
R+5Z5+G2GYT3PUu4FPzsRFvMZI+aB7Dsn1elgL6T1+helQMMenMdJHRee2HusTLUNMRyJaKG3wKq
jtgslgoHxK+NZxt1YsS62oJBp23VxNzzRcKrl2WOqifXRTNkSa942x21Llods5lRc+eMwrmYN4v3
MXBy06gWMciDGuIfW6olUW9qsheE4BExUR8Qn+xsf6HjJza5N9erK75/39I1gOkcejn+IOI7VXYM
ncasqolQqA3allk14uFtTKdgLuKWdbgZfstP29jpcb0wm64SmmKB67+UfMf+vyy6dyvtjStzu4U5
GkD3U33exorxIZu0HE9s4aSZmup04bPZJs7u3gVzMS6ajqY4LN+XskS2TS9ZU+8nS+N4hr3ZzCny
QbuYpxAe6Qjm2U8A/hny+PoyQVchchm2C0L0ZmZkYNfNrRNKA2P/bugJjdMA/TzLAxTFkeu+oid6
W7ObDpW5dDqvnJiXmU1wEaThBSGwn/nZWnVJjqib9ceWjOO9pRWkunAWmhyfges52kP0JpOvWrBO
Li07AH2im0LWbU4Gw4cEZKC0Svw0LCqjCBaAgBbYBhK3ybYKbt/bBCtHbZY21DAlN2TQetofdpTv
c0SbAE0jyjQddddczpv12cOzSqG1mYeMCEJFkwNZcSIPLSvJ9HKejBmIQdHq+AW+5pxERvvQtbZf
fohZr4aWQ/VIYiVQ1qxVVngu9FHwRv0YIst8EYa99Keox4tvdIpgrLhSCDTV6Di8H7syrpoHn5Q0
Ak8MHExfow56+QznRTahOXOBl4pJ25w1OdTTEQJalsi4LWnFneS+NwK7W+yy/d6dQCXhKyjEspTM
/yg4h0Xfbp7sthcl4/xkdIerdr+BvNXtPoAUAD3h1cqUyM2e9iL8ybTasvXPDH1JyK6Yr/LN5Tq2
rnz3Q8pkrG4R03pQSIGsDuYaij3rdPeyI+RsK7srcLlAORVzYUoy0Ga9PpogOd+pAHWz9CPrn8TC
nOfS2IxLPIRhJZPRgPxbg0YrtNsrrG3asg1q2LappElAxJAsWQEQw/fBFZJ3KMVjgg+JoHW8Sbf5
YBaLhdDRyW19ek//DzaUWgYYMQd9RZxUs7Tu5YJVvcxC6751SWYnMw6m7QYyNJWHCVwTO1WAN+xv
D/KGifeJf2ie9coStAQGxeY9H22TIlVhXrxdTEi9fK6014SyWWVRmjuO9yeoGSNI92wMhmpwVK+E
eOY1YHic+hLc/Bp9+19gkQdXQfLq/buuxhhXJzKFDwmBV5LKA0Y1ysgZ6hdEuOOjZT3B5Ge5mG9a
24ZpmwhcATuLZFcfnd7UcmWxGYiuEStE1WbXBx+MDpchSrBcZtTkRpN+FOZ8jQc/ViWrGmuo0yzE
24lBNU0yCVgcYD7lhQjmbEbH2DFd559ZglbfZLXnrTI0v5/iXqiJeU06Mb1eDQXFZ7adGSNS22pf
Gdq+ZhVtvmbN87DWMr1efUQCfNekHNCZppwImKWEMqxlpbSf65zjgrj1BDPGkj3fp8iWtLo/RVTp
KuPNobBXTAAJt17nmHXRc3+WBLk2udOobNw40mS1p2jZ6bn3T69WFFpE8pgZAacESzWtocrS2qop
tX/Ty/CIAIOqiCBAI4fy1H8Y2Mulu8nw0A/QPhiSN/PXGh/VRe9+XfNMpVmq35L1h988HCIVOUXg
vUrwgXXBeViyxcpqcfooNFnXL3cdyy45YD0nOdB6gcd1kJHvVW71Sx/DBuYxDwJX6y1hP91TEG3h
KXvj25es86wtEk/+QxSlNneldWIfaGWsepRA4gseYmbnt0zHnHIboMA9vO16/eZTmOZazVF4qbIr
ML89LLUU80TxJQEUAIhZhPBDisq96dzYY3Vaz06Pd28/5jmAY3SEZ3RFYMTzDJ+KnOsRV6EVVQ7A
h5cvP6531z9d4v3DoSmc5Mlx2C8d/PMAU6H6Ktf/+fFFMooNAaE7fVsF/qnDIcSGmHhT3Y1L5sT0
eqk7+LS0xRKhpRiXRiHCz2kxE8cIFw50mz8ipkmB+qUx8bLdN45q8Tse44z9S4SJBY5T1uYium9k
jqIs79UdsKPVCXgs/kb++487K1NTDpuTPYYHJRdts1+KfRlBd1R4+DpE1vEXmkYiMb86bhNuGPuP
LYBi/1IXE+dZgrPtMAI9n4L4qBqDJCC4RjcTAb2bZlTDFhjPvx1pBK9gWn2BUCSs8ipg5BktUKlr
Z00JYq3PZdKxa++9GwoLAPC1QDIJzjytVNEU243K4HfI0j2VAciiRqoxIx0RiVqzkP3ezbga0ZQr
apMa5TH9/H1xUgDhqTQ+BD0MASyccpXET9cfa23mWzQCYhEsMr8jbPsZnIWj4KNiBmAweWRSHkqO
JCuxDt6bUfnUr96cbOzalWTUbmEFnnIJsRJ3dCadj5A4q55lM7ifV/+egCek/tAr7G7xsiyUR4be
rKvuPRyi1LgYfNKP9iqPjxxL+Jt/z+qEb78bQRMmQu9dBCssRm6git6RPwDMSwqUmtmwjSZQmeaO
mtTelpC6EpHV1oLacFsn3OefGgfzif+u+F/3944sx6Ejt46qCENISxEJmOPK37lZHrEBM2W53zbq
gUvJXo5wfjmagYHnBPSTEuhSOCnT2ki4QDzpP1p0VbmNeNhWR4yyAf8YVhDbDIHCsp8s8Dt4DMFb
iEEa1OhnXRaUQUuJynl7qhtc8aAdXasSsGGjh8OyF8XMc6Dhak57fbg7IINrlJ8gUt0jnSy8aQnR
sEatMyFx19nq5qjI8sXkrHpsxaGNwpsrzY0RFA6DR9xrHVPLggSrDxF4DyF/+JYp8811LYGFaMS4
FYPPH6EEkCn4PIiM7n1lDrAByj5GlrFYSnuve6Hj3PrvpeUopqBl5l5lYJ3kNM9eUp3qZdZVOKiZ
YcZ9jSudLmfeUWign7xpoWS9DOkzKgYM/GbDIL8w9tNYnLaJSl7399JiGuEyBiZin375l4CLziFb
upuvcOtXJw86H43OOloEMncpwikmcbXgIH5IaUMZGnyO7AkKk2z24vxNBqJg6lT/9jNsyJA50DoF
krJIetaMru+zbWal3piVLGch4oL7Afu1ObLy8gqegD6D0lGIjDm7rmh9wT/+1qFNUFrY/OMAtGAA
23c3FDcumOE5tFV20mK4OmoVs2ZzcltaFCwDDIx0b9C5BJYJiP1DqPirISpOe1OnD6khLN7OHOSO
cY6Omchh0cEqb9TvrJwSzb0IT1Sdqy82vzwimrqA1XJl8lVxDlGEuP1hgtwqdwC66sNjWC+cM0/s
+cVEiVhEjU+GStJmzdu5UsTKMsu828EO6GIfMHsvH7N/DDj5yjZ/yCXuMNit8v8TxKQ7SGlAmC3W
60CpQFxjEgEc41uDUmYU6FX3RLpvBsD7BiDEQlUVR9YBSH3f3/uiAdwu82fgTlrt4Oo0iQHHI2+U
BYEvJ5Orvdpmtf1J5jHnkEJspnuCseJQaAnWi3+G0uutXyLlctaG6SMBr2eW4M+1E8ZHYtFXEoTA
qWo7g4fe8n5ORHRA1TJCuXi4QCN2hw+6x9FxSaG3RwloJ6tsZNEvpTSzbmlQHAbMxiWqDYq9Zh08
QI0vPmA938et8avxcQgVSwFFOFp5Ju8NU2g/eHCZ75hSFTKOAQA2BK/vimlShrUlBSMS0qclbJ+t
wIEAUoTjecTUFZgBXZiYpiOjwiDe+3a0RZYl70mvWSyNtl4X3ldvnxSM2++qdx6NlND0+XdEp1cN
EsQfIpB79jcYO0bSj8Bw3nevJbn9GkG6kigwOSSiDEMBuY9yNXc6Ezo2R+fCqUD1VPADV8tR3ADR
bw/vYdbuwmmcw8jjITzq+NSMyCCgQNLdmwmT23Ve/tO8GmgbAM15+QV1ldj7iwJxdWfWS7OAzY2c
EyOJ9C51reRbhKhPkozdsZqeTnWXlI4ke6mLHW/MOibzKpEDXM1ENHlAVGchAA3OH+Cv6WxMUeHf
pKXwGl+wavuOBEG4Sea3CtqKh0zyuo72JE0mqtAlOVKcs0o17D7Jgdp7h0+AWibvj1OsqsuYuIg4
KlBKPBfX77iDaIbdCFeJOil5MRTJVT88tuOeEe2wi377FQ+cIiBl2aVJolnIvcbaR8JjnIzBUsfc
RSHblcowYtXr6z6oMLKNXTx4lX8p3+m61kP8zs6wzq47HYoOR8LbOp6/xCR8p+4R6VxSWcbinUE/
jeX5YrX4nDzJ54erHPDXqPAygix/8kiUk7nydPvqKVkRIGLQ/VpVSGOOPLHEZROM/dF+P4vI47Ql
RkgkKqQ5P053XVVfoIDD1wbjqV1gjCYZU97jzNdVW1+b5FY3GsdwYFOgKptKSQcc73VZTSkFAcLb
Wh9xEtLDkSU9T2DndAPz1NH8l0YJQFazKM5CcsEl5njmTBhBb9FEi41F35+sGTE0YB9rApj/1M9C
yCwWByUYEyQKK5ZXJ/ecrrc9giFQ6G/SWBU9hbhUwc7a347OVYgwMuowbHVjCmJGH/Dsw3KNp/Gf
/57mueeKcaG6iU4/SbriAnMHstvn/XVdEoo2Gf5/ZZUl7BQEo1cKJp3eNPArk1Yf7vxUJEBNSnc4
873XAnveAffHiteitditb4d1ytofxH9PceY74mfgY2Y9uLdcB0JYRVC39PED1Qg4M5+z4ofUB+cb
AxTrKKwt8uPHTOiSoL/c4MbmY4QKROMfcdKotcSJ9jitNYjKqmb34n1tzxx7CK06kWP4GBVJdkNa
/icaKrZylr9ZkFGKXdMLOEt7XQM9HPgXsjsO5xynfVKNwC6PKwz4nBqb2mdZfXjBkM5pd9/g5bHP
Dl0S1603wO/nIJpdcNa33+ft9q0pJ+/AoaSQvIgXs9OHl5I8URrDcPlSBRiIj71dryjcIskPYStD
mQWxx21VpObdwlRZyr+YZUFW36BYrsKWlsA7KDjoCSuq7xPonyKqMR01pvCj0gKVGNroSZmGXYW/
4RoZG336Fbu5UIjk0xbe8TwvjepPzdt/cCSGsfmQcEKye0qbVCh0nKdC+5x4etD3fq6r3zV4rpct
/3xpymP7FHyoTPOk2iRw26cMTG3hyzFz1QPhVfRD6d0tpqeAj0hJLvsNFWFU1S9T9eWbo4e9r01y
VMnh4tHarnhwZpfqRnFBSgKWjnAGkPFTOBbHQm2/ARTQPQk0LktiROuSrCFoSYFUdXEkHbXyYrwd
y35t+IRzP35CZ/SfXmeJkfHmNoV8JHTgZNOvqUnNo/eQh2RYP+Ymw7vm8nlFaPc7LoAezaNREsX/
bySFglgRqCINUOQcgRZ/yCzd9LeXoo4Rvg==
`protect end_protected
