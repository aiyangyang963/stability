-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bDDUlVrG+4lkSUXtsYWdIaMPTXYxOqa4c+js5I24L3LXNQFSOtIHzr/rscDM0P7n4e0hk1MYGJMG
4SchHg3E6BHfortQ2zKdhWMycR5K24BANiiFBfn38p4eQV3LhbDn1BdJO2Z3M8CRurQK4Y1DZbSs
cZjJZKGYuz696D+nF3IywqUnZKqvXG3apM+4f0erKTZhN9Atxn22B+erYQKl1EMmJ0LIcE7GsDir
8weGx0OlB3jnCQfJyjm7B7V/hVfdkRcG+bcp18CL8NxF+P+GQMF97mR6D7eHEAvPnk58u8bii2En
dBX2Yw5iUgxuZ/OPtsQcD4OFyK7FWWt+E9feVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
KX5JWT9aB3Qr4svRsvClI8AeauRf5Nh9A3ILQglWF2bU69SHdrLwgAk6vmQppm3YWD/qc+GT6QzI
+O4M7i+TNIGVaHuLwGD21tZW8hGhVkt31cNJMTRAZpWeeAx7gDONQ/8c2rufTtkMGnx326x69kI4
2MXcpXPyKm6jlQaDYqGML4frxDYHLPQBu4M1IeMi0h7/Z3xCvKIplR+H3eqlGnTScO6BjbKqOop9
5LXdAaqqw2pOCJPkKnsZHF26sCq4wIQgMF61gslCuniAL8AWq92j/HUzOoCKG4ZnjBExZvAzMqCg
Upe69B3qENTkFUaxDAQZIk2oUs8y4iS08pdO88WYmo0ab3RBjuSIwuZ1Cd8N5xULYUS0yzlhxtfD
Zdpzsi3yj4KGIBDp+g46MLO6HFGIe+t3RPTMSHpwTrznX3DeH334tqSexuWcBdlwgwlVVKhRrx6w
o34Nivo3ha2tSBkNT9pL+ZBFmVG/QAGcNuXrQ/Z+mmKdRw8diwoTDx+/R9XCMjiO9EbN6mUcqK1c
y5qQlvPjqZ4oi8sgB/20f2nW+JYpUp/9tusWfY6g8ohqdKt9qGk42UnTwNPJLuQ3QvPcoEDQ6ueN
1Hh+qD/RWSE7b4Ywlzqkim9Nu4Xeyh+EgLK4Xf4uNA9Is1I+skbEU60Xp/+7HtiTU93NStoJO4BH
wi3rD8M2NH1XbnavzV490Saizd6KJEYDKCLR9oihc8cEDAj10qgfPHIQlmlKrH+gRcHhbuTbP/fa
LlmSlljNPE+eOrru8jK2EUbz/Bbhq1ta6O3D1X7LzG96u6BFbmGl4qqP3lL8Jijs5uCBp95ZGWdE
j3Ym+/d7MULoP83EfsKw/3kFeq98FRsooDUhCAsG1qzytgqnyxzU8fFmGOZkNDE2I9RjxWtwNJbb
lP+YTHnCfpBFYRiWuVD3HGbbOLsUfj87aqW46XLdqrg4vLXD0wW4GGoEdowWqkf+CUsyWlDTHmlR
DCX6BQLfE/9JOpqnERMggw+S3tDFf4QbmZUnfL2JFe8Aqxx4PIgxBk5zAaUGrR1ZLQ4urvorWP+M
fEq5BCtjHbZzQm31j3QeFjL0FCKfvwUlEpF/sSm47/xPRu4A+MrnX9AMxyNXXYzGJELqEE9yX9xG
r6OpfasXTkdVkLcqRnIfKEUlcT1iynORGryJpvYs/4V8yS2RL+AIzzY9tLiqiVGhXBGGF+7BpB3n
DN1U33dag9cJsTDhqjYs9naTG7Ic4OsJUCULg8LFhItKZnzTqxfGz/ntVCD1Cd6fzx2dhFhABrLs
WTWCmxKFOCTJNsLVS98JrNqBv1E1U6GkwPP5Vx+N0c9yp0zjNX9FOgfhdhgbhweGoQQ1ip4JtTIn
jI2KkYPbMbOY14oeC5Far1kSJg2FZ/15Y6f+3JI6whwEy3C5bsQOoMgmuGTaGwXbBy12kbW3ezcS
C6acZCCiinKQ2DHpooMPfPpamOxWdjjk1eoTtbADf5gvpFmNAh7FqUW+8ETzRHtQEpwKrJmwVqKI
ac3Zq1YIKFCOpis7k/5V8ZAj1kqxAo2BHhO2prMM9Fiqai88XQDrzZsnN40j/cqr5rn/jFErLxxq
M+VQV58w7SFrTFVFJRV+ZWxjnXlJ0tFRgJ+Bc3hajRLEQw1i+OB2PPoLEG89/eWAyU5BLC+wbYE1
y8gQJUIaGuKFHmyRcTF5DnUlBd0ObVgyncHoGdfA1gpH5jGGDqfQbElMXq5/FXEZM8UQ7N8Tivqi
r52EZQwkr4zlFHgzAwlXXXn+QCqBc+7UwAnJ7kPtqQru8HcgQxOiEUGXGghAecw+srYydGwedvjj
PEqqP8kvht77DJt2+XmeDSaTR4Yj2pjsZSZgySuMtHKb7htAMYTxiVxiGlW2Pq2qDVkcut7GQC54
X1NEIlCTuBcgD0SfDk4ty1e/aJmAcLDuEsPCJXTfUIQkotQhUKcKIHlxyP39Z2NY5jvJjH4B7rXd
PDZVw/0P7OK9rmMb8XbTsWT8u5CjIOvF8MZSvafpLLUPjmTJ8ut6RZ5zggJY/F1H8Creupk4mtYq
XXtsfPOJR+0Usml+UCEwYFC7ck9fvEZMCtBvft9iN5rOCwuRD4EcEC9xo6oEYm0u8KVl15ACuyJS
lEc+9xcZ6GX7wU9foDGhagZ2oKQurbDsLyyK2ot1LNSNq9KuYOC2m5STPZQmAVwMaUMm03asQDku
Y9tylSnbHwkKatcIMRN7sSfzNnzTngWGxU7YtGBE001OwBXi88QevJE5fpf8X0xCwcEUw6osoZUx
+1O8kGraei2A7nHz6Z6BLRQ4c9NJ12LrBsyQaXTEI/t71s6dvD7dcyVz4b2hlh1oEV8G4kiS8gMI
dmN5KIrIj3D4oaIVI6t3MmMcGSzLrGbmJB48fSbrCfviM0N8WjhoOfyMdpQVwzqXTsmW2cxp41yM
DsU1b3GjftvTyatIv0SvFPRNcjXcqfHmUjRmM8M04Cmcla7xtk67VApp8l5xwVAbI35IZwJkASa3
2Ggm6oeSY5BjA0ozyfE2J1eBCuU4wLLCYodd+6djlX8XoNFuomW+PVGICNYXFzRhDW1R58qFgiRZ
l2+zf7DlrW7IVw7QYfztNfEK7BuxjwJnipXSz7N7SonZyNl7N97m1CTPT+cfSWATXLIPc13Tytfa
ZREwSgmXEXzFvFwXbLzpJHGSSBkRGHwz4BrQWTY0lv49D80o8IMk/h1ZcDbM9ZOSmyTcHCblplhi
uHWmfatNOZa32/pCa6C/X2xLAnCwA33l6DxC1ikYhf+1VV+7eb23M9RM1P7tisCrNIJE6iGKwF2r
XFtMNT/UmHYMrXSR2+Jx0CxvazYveqATRRSnNd5Vhz1NE4UgbQiMMnNidB4YpgtQlvDRee1bUxeM
wYAH1Ee+9q1cAytNgHr+UhBidCc43lteWMw7fJ6qfmp5CJkcpwwTUPE3kCDD7BoOaoKaJAItIu8D
rdYCKE+AnnYV+039a6hGDiyYa/NyEHpT6TQbADp0IObl16MD8W/pc2c5hmI9CptXSL/oTUmdEgwb
T8I2OAjxa7Y2Oaq2MzDIQYTVg5wr/51/cLRcVQzWLynscNS/KrrkHbPYf1aEAdCMQurqKdsvQzkq
MW+VENzdPRiKTxdJplQ5ZN04rIJpbAwi85h8QZ16lzMBOqQFtRulytPvwUsrBujsuYht5GUCT1h9
HxSCxC7cYu0Sfgg604qidvR3OeNIOdIWxYZ6u9/iAE08QyX7bUN4cy4BEq/EqYoQc25WN55ZMg7u
dHX4WUmulsw29iGl8CA81Fin2wJM3MTDprTMsU64ds+D7MxWIFax10mxm9LoSOkcXqQ5qoL8nsb6
D4oDkwFkDYZzv8aIBWv1i3kvBNWF0MeZ26Hx7tso/BYINnVaHPTBpo5pJ7kePLsJ3i+FyX7y7p8F
qcIuKnSZHrfiSApegh9bYNmWQx7JRZ6K8YEdmalFuA0QXuGNl0n8yJbL+scWi3kieF56XusIeNHu
vOKmCN06cfHHLM2hfbvw4dyN3o4YvxabzwaW1de3ix2p7oRIsDJ5yCfQHUjPTETUG8Hc+7yB92df
mw9h6zSWvKtHhYcIRGeTeqnFIsRXwKxtWo37oai0NNxiyh3E2Xd8GQD247aIv5dw/hy/DU901wn/
5V8srmPTK6BMcalLFJvq4W4EVJs632hzDUyrGN9uS0czWDpON4tf/QbJZhzMUnQc60AEj/2lmA6o
UXNuzNuVUNHl5rfkkNB3/MoIr+q4bMAryioHa30evNgPpZS7CagmLgoIX0WzhLi8DwKX9j9CQf+w
77+gi0D8ALWoDixBqc49a3wAAAquJKqHCIz0PboUsKAkikmpMO6fqMgPyPfQFHUtAQxXiJoIXdhh
hMpFraRb1CBFVXJE4uuseFS4UzeEgBI/u0AelQ0CoNlve/qIAUn/xrKe0wBOp+rn3hF00uKKBcel
B6x8T7obeI1pNChcR8uEB9F93XtaomSa0x6/KfwjhwaJ8YzJSUMxokObEvMTzVz620M7jxek4b6L
WfCL+oJpnuT4HBDMdu95m7WbQsBRS3fFXEpcT/Dk4eGt/3aUxSrtARbOtcVMO2k6fPNmseBxU9ok
32ykovarQAvs1hWdFRGyB7d76DmJmt9HbbWKU4znSuzPsciTUSTdFxHnIKn1RohXke9h1y7obVyh
QPL0Hvwvd5iYOE0ijBR0git9MLfaBiAwAcfr6Kvj6bE1G+gMJS9KFgoBHzCeJgkYpxAVXMkmmPZi
J6JXTRHm4IgBmeSASwW5Y2m0iWCbijcfCs3lVRmuVX/++ehC95jsJnDmTkiyeWWK/LS6Ha84B5M4
y58QlQQHvubZc9N3u1tH9Wup4i6xbD63Tpdl5O48vXS3XgRVmlYuTmDO35Njl7C1xSoyzueyJGU9
8ceAo/r4W0/wp92jJWtW4kuw0k+yNmjTIWVwFEpKiI7fhqpGlgpm765QAhruLoyFJlQ8Y0ZNJHLU
H3kVTBb02AqMUuzPk93mInDijuVkR8nHCt88IT5m2Ogz2OnB2ELvXeJ1AQIpQJr2M7hqEX+ySUwb
i7ZMjskUhAaEEUqKFu+6VAN74gDMFHFiuwPKk5gtnGzu1qiZIMnk62hyjVcz/72XN4u7JZxsK6Fb
VNnwqQPfUudAgeNriPatLl4CXyoyvd0UpsyZ/W6GvAN9X7FkeUZoSzI8l0tz+Pp/sKkLQyRKpnKa
qmjyXHFYQKH4LlQKVjIDK11ugpcIplGhA7lVVnXWCW0v9edksmWfQHLgBJnRoJSh6hgeDI/vTV7k
jWJW0kI2EnIon6JD8p9CJG3Oz/YsGnrIozYv5K1OY2ONxvOfUh1dOzo5jEkJ9evYzholpc8yErHs
ZcoB9GFPpm44yW8VdHcz9SSpVue2iMbzE2//enEB4/D9WSgaZe9QCe9H3m+Qm28822x9JjhPqERJ
UJ+TQvVLULoqJypkLxxU9k1M288adzLXTXtQaT7MCFtYari8rvqAyiDvLr6C12vtuexDr/QoQrCF
CZX1VU4ToEMc4kakoVVUtduf2VlB9D3nzqCSbK8ROmDrGfhlDSA6E0Zs0L3WLo5Naq5l/DKFItsj
d333S5H6YVUsNK4zKhZzA9MgNedQrZGWd+xboR73wkz/w4MECqp85wjsiAxDV72JuxKiAN5c/nVe
atQDIcreAV5mRqPIeC6UlQmjxDd1wcjz28OgrtcSBzguAVT1S5NSp89VX3I6ucnlIoP+AcVfHpDS
tKlo14WOt57XfFIMIOnO7fGgIPCP7VHCB/ToEojtvgNWrzbYRxsBGrofENp23nmsy2w0VOUnyao9
+zft6zI9gNlrtesWlogF+V3yOVVfOK00ZaSziCgfNtvsadoOoSO2cpjgACQPoqvTPrB+H/V2ovcI
kaHbeIxx4bY+9iiwmbRjbsx2G2cddwVRTUJ3Xr0DILV7VTn+zIhLiYRXw40+bdK6pkmd8yFAjoa3
6F1AzeXrlQPQ+CdFX3X4fOpIeOQRW531EYGtncsM9HvWSLlxFpaa8ThuO0dOyOJp/ZkBBRPPehSn
oK707wI2K4CXXZHgrdPy4GVUW3D7xNG30jrBAn0ubXwBtFY896dYaZJc3nK9PKz21Pruto+cFnHj
R0XvcllP0+wA3NY7oLo9A3FCrHu/zXsX8UIj/HbIQJH4sFPln7o7Q+/AMP/E7chDIx8jan6q4ugf
bViSe2WDWpzAUs97rV+hpZRdUdy5hlgxlze8Q1Onun2Xo7rvms5sxD+40oXf/2XEY+3ZCKW60B22
TgMsTm0BKdMN6cqxTxa+7D+zWIvaSWclSznbJ3q3u0FUk+G+7W0EGziEbQPyDNeCDOe3KeFEQh6I
BRAzrJdjp0tqnGIIXMorw5c5RuTBT/1hA/tpWbZSu+E+Tk2bhRl9rkQmQt/vCF3KaNpWM4Ebn0Yz
8Z+QVpMYXKiwM0+J6hIy+34n1x45MQIfcbDDphy3GZP1/oDiXid+/7NFvMMgF1OH+Dk8BxAo3bXv
yrplw4Npy8jf5rpoD53+AzIRgXVPrnI/n9zcX0xrd82/mNbcE2+/5fafjkJQacFw6le4QOEyzFfG
tU9BKQB6QRNid+ZTWkhSYFbfXwNa8ed5XV2h5ArVDoave11iu9/dUZMT6V0wSUvM14EV9oB3/Pt+
v/zTF0hL8GAwZglw/v/rl1a7rhlUhZmF7HnfW9R39LZB8izn/DDhgfwWHZHZldZ/WOWvuA5T9Lvj
IPWNcfaU/QBZcwbR1t6iSnfRvf+tC0nPdf+S/vVxwL5UWSHIiiGZLXgSFCQTWbprq05zlueXn7NE
jDCwJhZQyTSKO6mN9V0djqydc8vuFTp6kmAYCyRlgDMQGmo10wGSzge50ePnGmBMWgpohjmOkKXd
Ni5MnZv260ppt8AQ+7OwaS9O1Eu8qHyJQ2GRgnD/bsTwb97NJfBd3CiQr91aHUbj/Ca2c2pOl7Hz
yN/x2g82ZEBxFgZlOyB6bhKyfRO7RzbqhK8aJhqBCkhLhB9TXlXrfS5jddAeKwS6iYMS76vlFHFr
9FZ2L+TbHmsidju0yrRon8dFhCLsBMoj2/Cgqfz0FdVNykiYMTTzaNG/LN6o1g8U13UFslkhQH/H
Ywd8cTvKlRCVu2pCayQkd4xZnfhrg9++vmdxK6plYLFD+a22BpzNlry3uqkHAFw81zFNuCUSJbMl
OJY7Jqj5QRyC0ooM8SlCTp1oP+GHD+vET36KdCW2qzdMDgEXWMs62nUUtLA51cx4FSUnQL0qknA1
SYf/U4KNGl5cVhtEk6XyhRbAt6z9+R+btEGygQzYYDscdsgs7hv5zV2b5MQ1TzBABdC9Gj+GCZCe
Q+oOk05AkRi4QhvB/ukxs+T2z7znID9TO6bQQIeR8JlJhoAX0pNRc8oT1IV0CedDrgVSj9rT26gW
BtSYXQQPSzxsaD6bDfu+/Y0utPf2UDKtgsfJjhKHwa1qKlYOJbF2LAk9QpVsDlnPFzfYClo0Vxqa
BxSBDVCPZ34LEYpmiAP23VAxz6XMcFsUf7cwv22d9WvuwfOVFCkHyJwAaTIicBqBESaGnm4cg5c5
K/UL8WPG6PIuvwupShJLIjNzuYKwVsh7lhlCkQ6hTOMeDXrB3c88dTD57MQlsBxO+V45qbZRSFLU
F7nrXIoBiArWT9dJT9OA0LPIo6/qfP+B2vsI7AabwQvAgP3jhvsxpjtsn8q+jGXr9+Br6SvTQXH5
ccHBITnA6n4d82MA3WfgCDqLmxPhtQ90zT2Kyi83cSKQAi4UyXV8o0T7WLfk2UbvPgGinHa19BzF
Z96GHT1a62rScUlB+q1smvO/WuDmRasE0/VcgisDkIzVquQ9GcuqaqXQfgTOIvPebs13w5yoi9hH
pieVFsXa4qw02Uqnfjf1tm9oYrLxvZFxGW8f91u9r6g2BK8MvgY2MGcdMZQTTv4imNz81LoWSCSt
6dcvQKjqG0KQ4T9ZZFCw9exCLNwPSFotHgDE82esDAkY0IgABBahB1wiPDBabRHp+hMSGlTIqH2t
P/DIvq8avcOEmy9Sj/BvneSnu3Csc4Cu1gpw5eoCgcBhaOzpKB3A4+dWe6FY6XGEOjkiKslamgSr
QGR7GeHnEdWInWUvLBiQezNtrXLASG7V9XB9frQT5/8Cj4qjo1JZR/DaN7NfvGBDsZzB2KvNTQ3C
ZTeCEaDP50diJt6Vz7m40XqkbGUW3HKu41i2NmVHVmf+b2syJL2XHtm6MXw+r4CUsl22Y/bIJHOm
3S1MG/nXAopFeHXUcJ3v675oK/prV9ECJUYCb5p3AvDrNxc9m9MYlzSXo/QHMbex/pmsecsqbxLh
Unrm9h3frOMHTRUEasnhNCAjz++RdhyKZp0UcjhkthSjwVN2q2RjK057R39Frug0aRFPQAxDqPaD
pvx+3i1qZL/e8o71DyvazoAOWxloqasAEx6/LeVqafEjLLrgP/GsHk44JlTMw5FE4CFb5zIre3wk
22rcBQDqKsZem8L6ljOYVWsik5MvPHBKTHUp6WcY3WmpgoKiggKUF81tAairk6sfrJb29wYZHauP
aLazUk5JURqVYNijVm0kYMyo/yn32VlBBs2A3lTD0YTncCserWvlm94ZgALx6ByxPtkbXlQjpNR6
t2rnKxSHrzKUWIqmsyL8Pk61UE3wWGLXMpQwUARtSER9Lvxno/BoyFyZ5ie/tuEA63r3+J1VcLog
FNls/cR6PZO7XNfRwaFLB5/F2HnZPsgcZWf3D8JU6z28pPjfH+OyJQWkTjCFnlhu9hpNYd3wJWs0
DWdRotf6RiqtE8M8hyt2q8CWENXyNDn/xFxqKh3W1nYLdLU7Db9OP832Ma/YRfyepM1yFe8hdadN
HOqHFI0FeHu83z+KGbcoOrERf3s+lXVAwvTv69UnEGgdLkNh54tnnObeI4qeZNHVPzvIOwKcFHJX
IAOGMfbmdx9v4T0NbPxJz3bHNXesnAQ/hGQZVB4HixC7nCEhsQVs2wNuxFJbB6p7i0HWRLRsT4bz
lc5F1P9AWLRK+m6Ko2pntg84kPfJ786zTO2wEdg1a/dcsIRttRqFfVs8PJ+ychWOGg6e4b6CCw7v
PE3BxjiDqLdMlP49zaUKmHw+nUGrgSasTG8tDIsaPHv+DC4B42qkqySC89G5cAH0K5S36QvFH2CC
yxuLOkY4wz70pQTOVdwJhVYcEvbda2Uh+NbvUdijl4Xb2Kq02yZSVI5sx/CU97n/yHxWVqYZFjDq
UYO8oiucRPqrSLfsjhmBokaoZZkq51gvrtmU/BDQjYik4/SSniM2xQYgFcFJeBK22ChaMVbw0lDu
F9I+jWxxi/IZo43NCgpkh4u0sP+t4qsGubjwv8XP4M/1WzTTQmPPh8qMhK4TH7WfHn74yLg7HCxO
cxXndtTLqm1wjxWXjEoV5j2xMs8NRpOfdmwLYAS9sLoOsBf0R814ZjiEbGzhWUw4v0w2yjzkigVy
4R0uCL7Zhs4pf4A4ITWfWXsVX8Ioo3v9WCSPuyJvhJiFNWNb7ASf0mUTsASjTYCUWCRqCC5xptLp
jElFH9CBGiYvNG2dgJ7I1mu9ma3DoAC+SE2JVlky5rNhmrJqyDh/0ZlyFk5PCwPTfGD4wzqQONsF
1uD0E75IoULaWDT9o+0A2id7vyPTtE/jGb7yABPftFEh6y++79KchT1DXek5nc2I7O4RomnPueIY
I6lZlWXbJY5/mPbVumf61baqrykyn4s8zODI6kg65AgQ/6Z9C183fwAKLEy3309zEXFQI1eKX8Xa
mMML/72y8qgyfKszgQ+nb5RKS4rlTBvrwO1KmrrxcAk8eVgNVMLktOxWq3CYNzfMwMUGBnKkopkj
bscHMKi9t3V7I3FJhhShSYDpCyNdDuv6KfrqXjNyeACLD8gslSLXzfyd+6mtuXbTyA3wK8yqZWa2
L/zn7jhFILuMmzN/2CZBh4y760cWlQlQMvUryMoQGnunl7kZa9XXeyJfsrltSXjYq3uUeC2IqmZh
w8c3IcchX4hdslx5jv2bVJASvOMGyh3PRyxqozAqtvpl/kTbrphy6sewbjpAbWyYhNK6482efI9E
EnoFpYoTOgTU99cGFNppiLYohIWia5qcvL58pq/fdDAvgVipLTJJfoCqq5Ioxl48kXcjowmgUgg3
SMDTDssWG7ZGsx2ntLpEmhovuKVo0cyuY4ZyPjgcVAcKnZ7XJ/+2NGTkSvmg9mhqKyv9MMhm6/0R
aCEH9kFCUv1frsR27iwr6ROyknR/TXYODWk0yV7tvUI+dHJ9RVbqnX/z8A8g2KJ20J5j89I2x1WY
2CBlQjFVbwO+q6VRT5KqaZIot1Ta2j1veUdWrFUuPc+5wQNbLf5EV793vNO2RRV9rFga0ijPMQJv
wNFJFr37PzdZA5TJ+AcqAGWZMyeSIp/C+NIUa+bmrx+3Rqqfv1bFneU28jJJULnp5wbt47DbwZfC
31JIF43LtLBa0rR3bs22OCG+ZjfdhdvKMOOB+vYtY3kjF1kdBOYL/VhX/EdhuWkWGpG2Bv6wMbZf
0W3WvWzpbyqp1YByTnPp+hv00O+NjkF8XHMrAqmwFJ/H9W4f8baqLKklPmzdXa0ROr8I04OBDC2s
sLdQ/uhBGRHAvLwqgRaO8b306ruazi9uCZyHjtiM1gV2Hp4rj24uOJJRyiIBhSXL/DUCAhzE4lMc
le+/rwm7SOk9HMZNRjjP8WAjQ7cLtNL7tXriluX3dPtOd4jEOSvzfbZouBpQN+3d2wWBkw32cjyA
Q7I94JDPhyG9rCkj10V1q54YftV1NdV3JfnKBHdYx5iMQYukmff78+B/U9yKM4ugKIRNT6JCrOZQ
hIfzfIbUuWmHrmt18ROc7Wsdvs53NZ/wAJPgCdp8hA7KDvp8wLRIyolf92yjEeC7km79qtHOX6xq
ATXQqnDURqmkjZH44WTxU74Q/JQKOUw+c3QzWNXN7BmbE49pgfyFK4dLOBzGp5M+b8BeLRjUoIuJ
fxQZT7ysS4xbDWMOL4JqZBwGE9qx6NSSslyy7Xfz12/WgGD873S4kEcZYFQIv2TRb2yCYom8JcUr
opXLhqURoVjjgpqLRwUpWv98pwstIu5IpVszitAkx0GKN/eCXZaiGu59/enKNupt2mbr3xvkIIDy
5ZDOrADa9fvxTO+q86XRQcSc5hjxT3zdY0N0cLHu+0qpwAn2uloMkwAJevA/5p5UGrUNynZEGeU7
tYhbbpeeivIPva0pgA6/21RmblHXa7/ZzKWlqh4IozFEHDsQX6rPW4Nmjmp8lArumf6hlsO9KrSc
HqrXAuSAAmr+PboZs0r8uYw1+PDiMSXF8YE8A0p2NAJSTQOH91bqjGyCmbLAVT2KO4ySpkHCui/9
PpG03jI3w7e/1gCMDMU1vawYEU7GtSBrVATzfzgPjl5Gki19fFL2FsTgMcXInMJGu0NlZCvPOuw3
Qa9x57LHizXS+76Dd/HGPJXMa+EuEHtHYZgnT8TAW/vGY2cVretD6K2t1jxjq0qmKh9PfOSN2ZYY
hwqpoCuAIuavVA2CEgbqHHCHJp5mrT3eompA9APoktA8gliF9j+2hJBtU/gUREYCruisrm9eD2w3
/Z8RRTpBxpYH7qYDJKI9GIN/LLSSgC7+4a9MGZ8fQtAxoSh3cd7hRocS1rJzxFTgsf2idqucuVw2
vSBxU4+y8fKy4LH1AfdMLIfvSchQ/6SH9vioymttLmhwHY4MEJBpMhzQLIHMtVxvjbPP87ZvpUxv
oa5PuM6f4u3evkHFmwbuBsrilXBsvZCTF6UbC9iFM7KGYCcIF9oy2sWY/7IWfS7w7qtrZYV8HEy/
XxZyjrwngaYHay1ktDFpt3MEoYpJuVO4BHvgHUhd57x0b7y4X6tqTPyDmQRAULyb96P2cFo7x4u7
yb/hOiH0rIoLBghiIBfZkMgtX785fCrJpXc50SQZJHs5B2uFZzl0rb+2BQ2paIpN33MMxqDVafp+
OBqTmDEFVDoxyIo8ZZyXqynMbZIqWFiLH96cA0mVmcN3Y+ftZ7gZB+Tr1JRuvurHnVGKkx3dXhZU
9ih6x+j/Tmpffk9Femy/Z8zaGwUKlHU4PzZTrvH/iG+PWISjp8GZVJSjPouY+OD7lOpX878DrzEV
KwKI2Z7uDwB/MIJgDedlJBcF/gBq1QpLvD4NlUNIYxTjJ8qPQ8pC7NY/Njtls8XVhT29vcZ/xxus
2TgpA1uxRuq/49Qx+Z+NY9F47Z7CqUxZUbU5kA1Ig8FMCNUJ+W5X6ntVP8/NwtEKzkCTRWALhU3I
kMzqHJOeaLfaALFUJjCI/dfjKKGFiluNTYgjDTH5Dom1wukfjvywBVPMxDV22PnUWmaM99EHbD7q
ABbAZo2SxdUssi9HUZGcIuKZOl5DxGXkk3tVESHsZ4fV9lnokTELl0WZsN2jE2Tc+TO2OEeVllaO
6M7aQHnVgBD1XO2FBlPS54r0n6xWLJXN+9hOyAL3zARz2YArIBbvHh3j/W9k3JwPqrI1ZrRHNVXY
JxqRaHALwxRCHRHvOGX35UTYW3NM8DZCbln/EwN+NaphF+p5N96BgG+DM/Ax7KJBsulk7iprwHXx
YT0n6jlGpkXuTxlQOxtFnOEwvChb7OFGhzilkSxXAbtTDu8CPyHRhRh9zgoy1L12d+udH7cY3pAO
0V5NiNmdu5/iCZUiMpRBLnl1lYz3xjFAXaMayuXuXgwazu3S3NkvozszcwdMJacppEj3HYWNtxOe
zoBMs+FlboRpm1tXsp+7UWKxbBu6GZ9vZKX63NowirLGI5mihz4GWCePDDfTJmN+KTD7XbA7109a
7TVwJgNvbYwb6ym1aXg08U2RbNntn3coUpIwrLgFxWMEknZpKkVX96YhOUwBe/B7NtQD2dNdeowJ
+4C8fjFRjaSi4QK52seXNoesWyE9nlK3jpFBE5lVkAcLNJ6EbrbyOiggSmHVrmUu36W1cEnvnZ/h
ELQWqmwia/GzyztkWD1hlIZhhSnFsppvulS308m3MQg5VXRZi3PstAMRmong1pM8CqLXwlGwhK27
J90qhnnWyLToM49Xbo2fh7STbChefjNlhRdySZGp0octScaYyMoZTyTdWyqQTMJYf1fnoIhjlzAO
JfQ8DGBbIEnh7169L7MuWkTl1akaAG80Qi4Nb81Jg9k4W+/L8FPSzbKIYDn/Oznr9VEYnr+WTOdo
EUx/SbxuRWLiXXgs5bb5z8V5EpR3RgQdpsGRMez3FYRuUEkYZLHZCQJJx85s5pvBm/ciRXvzfBUZ
2eEu3VX9SJKmn5W2qM854dOO1/dPHTZFM2z42hJpAYq3fgoHkp/bJ4quM8vX8qQuVwTmyIgmr/KH
K/FCQi91ge9w/s/bQ6AELdDfEMreiO2YdxbweCi03civDo6mmCb6A8S3WPAJx92uSWzoRf4tfW3e
rPgZOa4XUhk3LMhN9b2x1MLM6hdce4xTOzhOmd8t4rfdRk7uiIZXyPEI3cPh0MYARM3EjkFDp647
3ihf0gAED83upLUjaGEmexx15Nf86GjRSNiU95CMYj3npROKzvU0D7agz9a+gTo+K2Lg5UeN1UOg
5xebSJ1J5uGOcS6o5zvob3B167y3XhaodanZ7cOdP+UFbV3sgVnW67u+e1Iqe0lEZqRrP2KBC0q5
ooK53bVyrt/1dZ31HyGxVqU7XFqOlXsNDxHgyYOKuBxNto7TrFgXmEvaslzOFxmdC63jMHDz87Dc
4MU=
`protect end_protected
