-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nejJDQgmy0J0QBbKlPunXF890N4ODY/nugn8OuCojHAClMXixY98KYYjwZxdFPF8EhCVdx7qH98T
ljuVscaKDp/t/l/95QknOV5b7AmX0Buc4p0GeQHcX8ff8AHBQzPatzyUAKmS8psen2Fxpsw3BDVa
H4eoFi7IOoGKHQPi2c9fFcw7h4KHgtoBQJVetY2QzMjKBEnF5I74VlsJ4I0m/EPGjouYyn7j4FRE
tKtEmY+AcVj5TRbAgOfIKJDIa4u6u8gzq0AlMZfKIgB5UFiU0BMNQB8SE+ThasgGzFHwJ861hrl5
HYOzfDFBadmJV1fQ1e6iY9r1JwsHO+eFe1dXSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
cq/Ii6y7EXH9pB1P3i+6Rlsh8kys6pCiBnfOhCgvdIe55CX3g7MjR1D8LR1RMcRlpalQxIcHwMjl
gY7le2Ee3qWocPdVusPa9RAOboDdvrEEtwFyeCGLb0XpEEcJFOsxVpNqlGoz2XnpdG/yGMmNpyl0
1Fd0DJgpMTthcntgl5KCx9a6sb6TzxFM6IHqA0G3GWpZHhZ7MGIqMaUp704UgRt6lnXnmq6WK6cH
Y+UH3Ku41/v7RePshtinve5hHs2PnSoiK5s+1aoQnLuQkDTecmQBGNJIpuJxkiHvfNsSS257GEdX
A2ZTxHlYQG6cfza4R9N9r0AWdwvokMpMTtrIi1OU1wHZb9DsEEx4xBN45NhvLC+017bQTsnjwJXN
qU03YR7lthhuVTRhFtAqEUTgU3Xk99dFmRB/qok7wQaAbfXNJALwdi8DIe2krEngzmRUrR8y1flE
sPTRYyps/tNpU3fAc6iG/REfkAi67HdC7kXAqkAz2Elb/70e6uDZrJMkCEaApiFp8I1MOJtzHt2a
/y2tzkwOI9/M4uApiTVPhaLrNiC82Cy9Rc3q859rtNE0uU+fqNZwhsjr2GYTDufXKy46WkQjBdt6
xViCX0V+B/5waoNPWyIVYckzT5frVV+qAoctqyAngjQo+o1TVJVHTFLkqQFYpNBPZZQ7i0Gfpfgn
Z2xGin4E3KxfTSlHK6UyD4xs6he2IOlS/+t8nP0zFjHknvv4Lcd1ARZsOrWhGz0xsiVVh0NP0kes
WbfJjpOr7+9bt+jGXpW8hdFOSR0A2BECUUoOjRkxF6GkqcHLKGz55mWNtApmAlaY278zuniwTB1w
CmEyXfPHI8nqssFjXqn+n2x+PfbDljrt0cxXl0QgQUiKCIXLSwYhPuu5ajj0FccfFConBYY+It86
MckULdo/9ocleRDw2uySKbh2C9yBzl2AO991IeLwK1x0ObhfEqQKDzva5E7abSEkhG7WjoJxKmf1
43kpxdJlmI3hcMX7885BbR+yjrMKDUYkO22n4H31hz5avccsLCuLX7/u2+mdGv1SDn9Dw3SGS8//
ALV7ar/pZNqS49gvxf4xoxgsx/HNcnPtdPqhIyTmKrrZDtIzeZe/jVHjqIu9+lzRYZZKPYaZ6R5N
+x8sFwnE8c3t0NMgkvY+voW5m3iKrd4LLDROSJcU5q2pNT0SiSUgK52nFxqfat9vEFyQ64Zqs7JQ
v9WuRwUwGI78wSCEbzxuFpBIgJ2nKVG0bP3FBsvGFo3zd5rP1HV+zHzxDdHCupIg4FJ13rg7VIoD
6eKlRiIA0b2wWmGqEtcVWy4zY4IBs01hOaFptUKyo7sG1HCEuZJ0zHLMoEI7ZQTWctiSSi6h0ni4
g6AuJdi9F4Qux/aoLhmwPRD5SDCqatc3Hag6SB1k6MMOwviv828AL3BNcH57XywLKyn4IWDajtkJ
gOTHjY+Mq9Q4pdTyAeLBmK6oQ2wcMizt9Q0Ctgp6yZsnyOmjfxRLXlbMWISaNYCvydBA5iR7Qtw8
sQluzF29BvmpXq9uW9uGUb0yKulyppnRAxnkta8JKuUXRoCmMNVFVEN0mu3pac5yIO8tfebubzSG
t+aUtoqvUT/vK23RH3uJCvC/SijG73/9t3H7kIN7KmDKHuu5VYka1tEAkfGuzRMt/v4TVmCdLJ9I
3eMngwzOghenG1tbzOpCuJqov0Zsl0LOaTduu20KxGlLcHwjW5ZyMLuhD5nGpR5CHMYTa0M6D5JH
j5iAErMBod3oHbO9+SRn/voBwSCci8O1kY2gl37SE79kpNAgCicDkn8DYMb0AhApd1KT2wWNV7GJ
vXWcmsSHGX7+axuQzXy5Ui5VkmpEljE4FhZ+oQgrGOvako437by4ts6En69/4Cd/CtRQbeZcNMJ+
oAETgJgSn4RbqNfspw30v4gL8+k0IO00/MvMHPklfnPMM0XPzRF1e80+weDEmr+qTX8KGUyesvUl
IqxpZ+QtG/woM71TeTu5/8rOhi66UBeuBaEFU26aB7fvK+DpHeQet48VRmfZpR1W+7dEIxpgM+d5
ajlF948G4dHOyDSqG/OsBeX00BW9+lNUNBN8S0Dr6lva3gmj2699I50/kVbXeKTgCC3+rz2hxXnh
i6YI9Lw3t8ITxTaUv2XhYQFLyu1uSbP1fCF/BSSv95DgtDlmXKdOLJ/+QBWKWgBZFA27bHGOY8EO
SpO2fgGy+b0vVycRRZYmDlcv3Ll1jXiVOdI4bU5UO2ZZF/Kp7mnOY6nheOPMTrxAvwn6EKetxsRr
EddBN0ut7E2IoC2ASmMz0fS1rSoalMz2xKh1rAjx6UaxwdeRw6Ll4F+TBSrsk4DGJ4J04be3fF7f
gRlunCIGjQLLltA5Gj8fayyS4ZsTL4KnBVuokXOG+mnnJukdftPKe8VjHAMgDgr7q7NjYZv5921a
ovSpKOHNNu9TOKq5ACdKanTPQgrL5BQZpL3zgRmMY3uYR0vTr0keJeFMT278RDuKn/LP4J+GdIxG
dYpvgYcJD0TEEpIKF43dQ8ppCfmCFoG2m+igIAxWMZ1+J2mrDhZm++nVeu9o4MuXZ+oI/lfrAZJv
1RV8gy4v9S3CSITnIUTcpwOTw3VoZwTAfnko1nEwN5JSGFNRpWAMqagadDzC6Vf1UEq2Z8Pkncuf
+jVt4IN/XcFCYzgz40Z55F/K+aiW9ixNfckPXLai0ncaV5t/hku95NNuZwV4TRMHRaJGjxaDA/hH
xoQKwFvZ1BQ31h2UOxe1D9I3egbprFRofg5ByeYJhH1HguFc6meSnlIInDvHjASpXJAvW8rw5xJ5
Z18LFKrAGiwa7e+EG6+qH+kP6QwAYt4lX8PjtR4cYQct+Cx+leRE+Ut3KNNZZuv6K5plhsGT2FXA
dzdQ97HcdK+Vs6XfXdWEC+7inX9S3isc+yZ7Ze/hqPhQBkc5ui8SlybISg+1kPIDldnVSCas4ybc
gOk7NoKFnLx2a3Wn/jse+60b03YpUUr/tNM6iJEorm21qdyIktgQWT08JsMpY74HCo+5I7syag+o
N1LtUayyXWWJl4vviJR7R3udeWSDVQP9RiY9U6GlOgrwHfUBqDmg7U4ZDnFg8R5+pFrKqgnoPMy5
yPYRpS9HANKXMbjnX4ehec+ffS9MDwtxJm5E5HZIN3s74hNiukMH3WUpCLEJqce8asdWT2v1riHQ
fB2ox82kIrPvNUFinpHQWIKTyKgTrdRY2xnBG3DthgRz9ayImvzPGLzlegoE+cjGoMFw6htpuyrD
LWvPyhRHX3eLAEmz07ilqhidwFuajvfEGs9h9ISSoFh9o6JPncQO0WraxxLlQ2U8FxyNf1+jIRFh
B0eRcDBXfOmp1WL4kLkQ8JYq9CrCfDjFt2DokTLcbzkzLEnsXnGxnfsGWTcZbmMSox1L4CF1dOxs
mrt1p35ObfgKUR7e8N4IRh+XDEfrWIgGwLXqkyGAEeLid+kAv0SxDdHqZXcg8bSpu+kGY4hS30kd
idCafzKboqlLi1f0C6j+afU/yJQudkIe6EyNaTisWpF5LzFcvZQDpr0UDIXyV/qsXz9N81ogbIA9
fF44SeIXzncnzNqcR2j5f0QX21S+4OIjUtrZB4+4a4YzG/WONNPhX+NsK/bjGWdWcphGVx7KGuG+
Qfj0pmRuWJy8SxSK56vdH4ILlKvleXT/CFFXwiHL02yYdob6bBYaeFrjSfVr9Chfj8UPqXfHO2Fe
NFp9id+oGM/Y1ORzRPQ5STfFkLx+O5YxPA067UE1pQnMtAgmBkhSuATACk4x5/dQnRpLAUHfMikW
Y/pASJXueRs6+6Pg0MXiLUdbnuXALqi59wsP3Yq7tjBMPg1EXXIDInYdPC4IOVnhUTQQWMU8xLhD
BoYa3VOfCmYfW4EYa0LPNezuHUE4XQxCPmkaqCd5irQxe9PdsdJXH2I6K7DMijCe/riSufo75zuD
jbYrhZQj7r8Dgc9cEMvuupacCJn7oJEQhV4oT0cz5xwQeuJdwzZKSW372F4xQ13VuOnXR/1E+cgH
Rv5DQgVUhjTWTu9vnE05mC6cj8oB2Y1OWd+/xZ/6V7gx+OTyTQSd2UO6tmhFgfajZ//ot1EZuiBk
y2ZgXwHeibLh9da5hiT3QlGqV6pQVDZ1N+FeQ3+ps8ultYGDmR03ocO/my1Ak834xSpFoQD4PSMz
tWn4uYnGOHQsNWFuOzMu82VRX7xZcr1ntH27ruoKuBJfXnWRQS8kPteWmhaBbM6+YIJpvJ2/Y6M1
mjhOrJk55bTuz2VNfJlQtmxZFOjx7jbL6EB7T2JCVGJEYiMz0wbP0wTcdQmCM4GH9Ou0Oe4RcljX
+yC5HBcdJiuPPtYl97D3NdFbIUyzpB/vYw2vCZdaipSeOh5XsVBIqsyJsZmH4r+7nPO3OjQESREq
0c71OHD/UohzJhYqz3NUeZzN/0a0HGkSppBjFCQ7YTW2Z5rPHg9ucm5oHJgapMrFCfF1BIk9C7d6
Pb+q8WAPhbQpX7j+bsFaX6MLBTmG3p6C/42nAovlwvRjM6Ub5yfJnzbFlbuQtCliRIhg/WRwVSnE
KCCDMOso5ICRXoa3AekvbKcvlBxz+L7ijTuwOPt2WM1wHUmdlO9le4s9O1UP3CCTz97HNoWZHWTb
GiJcxZmAr7gWOhIZrKAMAsh71YvNblEMgdPVEukiWkVrZ/5/d62KOqIB3mDhqAFa4TxiuqOwZUl3
jeljUADQCz2lxaMO/TwtsOcYgXHf/vLW6O5mjMHl/inG2EUjlRmRGogvfAOHw6Vf1OuSutFpgWCx
pFUfIRWPG8eHNSPELZVLhah0LG57E0vk54uv8Zhwv+ufGVk603lrjde/rTR/gP7x/YY9aTSO2CBR
rkRBNcW3udqHiEUjXEgW0QpVy5ULikWLqlb+VT+IEMhEAE37Iai8A/bUDqYc5QMW9Egg8UC5Pe+v
har7ejxEFulwSpQIQI68ho6wLbwBtif8+fUsdiX/I3Q2ZJ2B/Q1SHtcSrDKcGqa5j83JrBo87Dj1
i4Jv59IBgKKf5pNk16iNnN1AfnkVQL1o93hPdynpZ6OSz5JVj+Xj3xcNXGPIeX2tyopk5InmqN60
wZY4mwj+2UIQhjwLoukj+0jprIk8f3ui9+UFPb3FrPomDp9D9FMSoRIq/aoTWF6IRQRPvOmLdx8e
UXygLIKIG0xL6mXm8ap6yKDM13sGT53WlJuw4lEALsGXItVrFJkQvYEVU7Mq3HK7EOKwS4nf449v
UwQKfyH6nyZ/LpZMZcRkK7g6U58j2VfVKN/TD0uDhUL4cIFaaXWNaFCYDgByAcbrNBi4A8DLPCPP
g/fEn2S5nXqArbDa7L0IBMBAbV4VlO1h+Ql/CdMNttmh3ofIbusbNImr1Osy6w/vf0iJ5vAZOMkd
93eJ0PsId9dg89MxLL89KIgactoNFXgJ6ngvAaWABVLqaVjpJPlEaapBsPTKcfXWvpB9rZQiomGO
TFn+h+Eo2CR1LRtAZlYE+ap7Y/YTSfHfrFPEiwQCiIatwhndFX1K5puiAngpO+rl5EYt+1XhvjO3
ONgLHL3DPU/v3dXW0TkNTkltqlkki8TNPnTDTy2tPkCQZtCcZ/7oFEWHNQ+QCKipny4bpEvCtB6b
aXe17WJY7yrpZ1ZpVIMcxNDyRYuPPsJWBcNpQO9LJgkqv7XilFHJDDm6Fp9S54RvzhKCQia8Hj16
20wy2FY4iPaTAkeu4RX14XF/liKRJCwlkTJjLkNUkmwFuVA/3d6+vb+7NnQAypcULdco+KBhURuM
gtaMgSUpDQd6KR5dUDDqE1xpa6Klq3rOY87YG3x5juMLIQ7IAMOobpJNFnJTDz39P5vgqrydB9Vr
NHXSQqc8OiQCCg6Nz0LrqtSB3EmAXUQKTvuktE0Ue8Q9cJWKkdgzTzoh7JnWSEBRe9tOQOx0J1Vs
FzVmQVAtpokTk32rAVLeexg9lSYyFmOqx1X+eRqNq48gHDMNZKHkCISGib3h9WYtsPdW/VnWp6rF
ZUA54XnuQ+unxmiZc+adEtGcFe/h0RARh6jII4VuwDWrAqldXCOmJhWia1MieQINP6CQeuVEIToD
0/B6iJLtVnYXHGGt0Vk7T2OkuE3y8WVYabF1w2frnWqD1Xchaz+7mZyGHRc473UImznEOl1lxuUF
izQylPtvLzypc05Q0l/iX/k9/x5nYvO71jZGOLeU8vfY2hZRzsyIYwDRhP+/u3QYFJ3OOPWLBQvI
PjSHFqyk26UB78KzI74YlmlyOlRZk0WIdKVNG8M/QdBXb5GPz64Vn+l2K5PEg/7HdEcaJ8eg5Fj0
j8tSwC8shA4egdPD8PGf3Im7dCqZOsAdotX7IiBGBosG0kUku7GEWA3h+lbrSqmOBhXA5HV4fjrp
mO7zv/SxJA6EJjlAweIk9cHWjwYh35AWXk+O36B39dKxsAcScfdLbKSMgqqQtZgWPBUG1r+RHFaG
f6XIrOIz0QsnaDsIytp272F5R0ox8gQDx0ZdmV1aJpwnaZgkdDC1N3FXqAC9218dGQz6pxgU2d3K
UN168HjmavwYc4vzdy31Wa4rru2waNspovdCIds53zopDbubFLccoKO7hYtjYbqg5Jskndyym+Qb
O6RWLm83IGBj4nHQMihoxRl6gYaURQ7W5MvLI30u8xl6Fx9Og3w2B+JzhdONfgShSJdYaa8mua33
skT6ECCYJahTqbUP4qvugMWE1qlwPa/TU6p8pO5p4Zx6oTzAVyKF0rOi9/PrvUOQq8RFS+TGqJFW
pi/6GBDhH0sxMR89bgz5rK4Skylg9SfgDdPtIAhZgQUiULK386nEGzg2lQhfMk6RaTIC1VXdC7j2
zjj6hkE8BvyUcWndy47BL4uDpojU1Gpz2SZH3XS9tp0z0AGh2kHrnTMyCzL+rXx+aYMw8mYA5RH8
/vJm4OGE+dsSLayUKyGzsf9afHkA1XPYMRvDrReikiHyyrPJYkDzUT12pwVTvdlYi6ueRzaAx4KA
6G5x5gIk0GTFa189ETFabIJITUDSBPpm6fTP5W1S7lyoBS+1waUm2QcOZeFxUd6C7d5SRrhrICDf
DjK/RJwjn7S7ItxRmxXaOLk2ve3zlir+SVAdTqunQc5iPshOD+pdQs2+8xuZOlQbrDMFFaBiDfYO
wFohMVBrkgu5TDg6gyA7TXafHnlqDb/asq/2cWUWjNaTY27bYEryCEe7LNYUpxaOjQZgkmoqTOLB
xBcp9prgF+y69GvA2vk7lbwiXp/H4DAFKQpVOytf3f2xGRBjSH6/ur2GnDf59kZtQvng0vLaPFWL
Gn8dsTnrKPKrmn0TvU6c9oHWdFLR+Q4DglmZL5NDNgN1+TK3EwxiGXMNHP8k1o9UQTkQmP2GHMlC
NzOup91VSIHMMETxVC9Lpz58UxlrS2LERgR/HjmU+F+yZmslCdlGVep2TXTktWcbkHzOPPLXGE6x
26MIamaAC0H12nnZil+Cytv/QAE2IYK8gAjiNpFh0zb4D1YvtEwZ2aExhHPoKN0nog7NkuJN8C/V
hWyuy+0ABRWRG3P0zIenrTiZ9e+UyBSPEXt67a4ejr8wRg34aS0urAT9r/TS9Ifio8MZPmt4eiSd
5n16hUSj0EWi7RragExeEWaScfO8lR10rz8SJ8MkBelfuxIP3HH9re9POSeeOKNBU7yLpLDLmWBK
9+RplMoJfi1lTd5mVOaK4wScRl9DHSF3k3hZY/DDDmx6hrmO3VYEiQrtd+7ZcQmXhJGYN9ow6NRs
dE4ghWLuclAF8/zBWPWkufuahMVoJpUMPhJdox50aZuN9+xcd4ZhC7Zh8MnTtsNkMN3yAny7vpUU
SWumjjhsSNeR3kEFKuPLBD8cmJXkml4+co/Eeu9E8Hl5O3bMGnW9kpqFqNya2mfuBLbd6rvRdYE+
1e3z280uQ9qRc5wFr0z44P270AJoqdIkmFPkYoVUgU148YTPPVnf81wT+ZJPCfDsKAGSQBFL7scj
7Z1l1XboLvhYkQIpK1S2JYQflmF5T5v001jl3ZKMSVk696v+vu1ZDYfH+YBpbZ+a8X+/Zh1TFpwO
H6JnRKqGYZcJWkrQphv02hqBTcxEnvJvq4U2eZcP9+xEx0bpUK3otzDjNVBYVYHCswJ2ahOosFSz
42CClkF20EnBu+oPZt2NlI7eZ+3tOcfJK5EAMtcokhw1P0UCTKVP9Abr+eE1fzSW7IooTbKTuw2l
9kx0tDhXNUPQTM9KweXGAmATyr0hD5Va9GMwG+2fdGI2mvvnAO/5c9lu0LqI9ZNF1UP5+5tkBZlG
FuORTzvihZArTNxJVz8ziDNQgS9lBEX/CpEMAw/d91nfH+0guwhRJP8Cpyug67BnDL3EhbkEe8/t
MUeExLZEeMIoRVZ2vN6iBOeZbdQUnP1xL0oaX0SSnrwI4YLd3acVL0ZkKSHcKSM5cEuVHOpnj+wB
4vqsgkOtWhs/1BQG53K8NJoRCHcA0SKbE+4A6azHNB4F3k0elrO9bEpdiFCwA52HtWbt6VPEAn2G
ZFPYeFf+38gsyOyupZGqtBWu7uko3Sp3DggpvqvS4dWdBVSrOKQQZRcNm/jspZ+PXxESvlignL40
91zyAVLkI++v+mdreKforq39hG+9yoHIpQ9J0s3OoXOvIQcyuD/U/1Mcm8agvZbXa/Xg3Z9b6QME
Ejd+rIJesyRHk94r3znOfdvDW7rCUCRal4KmlqakiVXUz0xeyHOfFU9tohVVqgpW+eG2J+lPMVON
anSVd174aVl53XwWXnuxTjcUs81bBxCsqjeDwF5Yy3QtsfGCK6CyQXKEa1CtktuNEZnyyBS5l7TE
kEXQ3uGYsHUkX/DWwqNewdt88v9+GjKFlT2qF9XmFU57bg4sQ39ieNhraXehmp65VT647P0bj7+T
WPl5WMdOc1X4xTtw5hXmiwhWrvcSWvqjHVQUrW142MTJ+ZaMeIYQ9iTVRKDVIrZnjojNqskuhNg7
wHbbjn2tcC0wFgvOAQ/jsSgmgAB+eIXud7yHiNMdL96C2OMXMPRD3CVEFmDmElbG4Y4solDj3SrH
7U0n/hFuYb/avem7DOmXWEROxPIwGbzMsYpI67Sn5lBxNGifWxQFD0y+/eKqZfWrYr/UJHRuz08G
uC2CyR1G2cLIxtg8ZHRLBHSkryDONuhfkiv0TL2XtABT77uplA2PS4JjG2lgIQoSuSRRfEy0rNBh
x8bmAgmOExOZIYbXmnx+IWPMHJG2HNXVgmvRz47ZD72l4I4oCxX9gPf/cMytwxmltvCFn74SxadT
NwZ7cx28Z+cqMdzTp6tkbMAmDFrag/SVcsacsa9VSwA7bpkWvKBHtqSDV808IrEjFGquZNFu5qS4
gow6uKI8vPooQf0XP8cuoXtMkuccnL82Q2HQ0S8qMH0a543rMVn+WMm3GPlGc2e1LrCbMeD2p0b9
hH8L2+nQcK4IB2/dZwIlL62E7PWdDG1gyOfHwRL5/r+hM7rVsT1/O636Aj0VYiBNQR8DkbGNJiru
rXdGbvcaevw9ZRNnkEPk8CP2Ydyh9lu7z8eXMHHKIEKkYz5FhrB9cN85TxPrGJQBbM/RnP0PKro6
1Dfy7miB8Me43WJAWOivanEogmYAb/jojHPa9NrNWrOttpxFzFAn8iqQC/DBcq0DifThOnpyRnkp
EjUxhQAiTXgNWjwbl6Ox1cdACzscFFN9yxW6R5Ez9WRZtQXVWp0oeQH3FVFM3ykfUZEIBPSLuybq
md37XHrbwl1KfeKVxKosKQjiFeVsJ66eyIPfYXqnE6H0bJQwbyLWKe0PG7XPp9kbsgLvMaWQg2S7
Jj4qeiTsvW4T8zHsQa18+0GSQzIKSmamzqbftiEwtqYXI2171LiaBOxsV8TsySB3lsS6dHKkq6gz
er/PgTNR0bgeksR9KY1mo2GElNcYVo+pmw8Q/Ffu/svQxnOCZDE0K5TCR8SrCW2crp1k3GT3YTzg
Y4Q+hSFL/QcycGqgydTHq5vu7FN3TU1jK0ZoHxeL0yVr/vn1Ot6w1PQYqpr1JKWA+8B5T0V28j+A
XYqzZr/0bEqgnpWbUMXLsQZR15KYli5rgGdmlj/Ie+E46Ox82/xoGukMm23vQI8lxdDLNz+PyQAs
jC1fYLqM502YQoh3WD4r42HMbykd89XkNZ9dofkkZoXimpAjKid34sYIrnJHfU2YcqyeWLUBD+v7
hc6w9/HmNM1hOtLSIybzbd5dq05fE6jSs/fd8vnJorb7XSypS7/vA+jW6pkTgZEC8wvkuFZhvW0t
z7Aucl9QvqZD9DWNK1GBsDbH7JP5104p3v5V7chAgWwzFyX+GHsa/4nOWWojAki+Xu9pr1IHKYju
hawjUwIMN7i94QnhQOGkCWipoA/x79mHsjqcwp+L2uQF04GdCaDLrfPWKleMfIGs5hYiibwo5ffq
MKY04CPxSnWnE3I5FXNrj6E0/TCtHMm0duINT1SypcII/zIiHWiHuf/50l8hqLlRk7n09NivGaZW
9WljDm/GCqmN8poDMzFwrqVWp3DuRu/WjsaWNLm4GNuKmtdJ0yhxWBzyGWVKGrpJNI1/FViPttrO
rwzgUdrMUqpHkt5oy2uW5R14gOKDVrVV7Sd8w4bJaL32iIVHjU7uKaq/3y1hn7sSOzATMwMHSK2p
qJPFC+bnPhy1M7Sw2vHWF0nnKGtJFthtJZaoLwa7RDqKEcY3cRtO+fvtODMC08KwAZAv4nb3DKR9
DCXkCo9wDi17p9aCLgR0wADlK8Wg/ByxW+oB3Qr5jeAAQhinfyCcm33lyaTSWCa6S6laPVZ9XnIE
0zs5BQ7sN3Eo3rkaEtzsvV5c97mcdqfcwwPkTlVxU1SakA+b0IpEoBAu792RopPF+/Jf1HzTN84j
Fcm14xbnZPPcWCaX3WFIykfNdPOxneNRXAxS7bbOSQVfCUoTXWbeZzCsIFJzwDEeRdiXj7mhTGP/
2jK5rsnpKbwgGMaXFd8THiCA6HCK2bGPOzb2YGE1hWQ7DaJx5hd66f7tXX7keyXmcxOV7UW+Y8AZ
ZM5ZfriBVzLXl64Ru/tdFwTcrpTIiztoNalzrIHrXHVBOo5dm593wekZOuWOH2A5+gXC6uCfzPaH
M+6TWA4fZaoHQrSqZMe9EYXwvdCLv1D8qcnpX5aRtoy7TXrZux0e429cXiSIRb9YzBoXPJkDiK8R
N3eerJCnBlDyqPSy4Z1auOGsxf1I8EyNeXvBEXmaZzqIgj9mhBHI3LJpWGZC/wSNHEfAQ4u0TmEu
P3lIp012bmwK/94TwsrHO97E2W+KkHCmVnnhsC07RcC7+h8geo1WEsZ94f2tyzzWTEUB76IihDTr
YKqI3XIkeS607eecFvUzniSxQyCphX2CbQqCiX40XWmNsR7ZDDV5ReoEuxKy/uUjLd4kuIGerdm7
6Dj4uHJPxOlCYzWBZQ46z9E9ufR+dic5eITF9GPuLul8bMOIu4FOe6awFGym7ULM9oBsbTD7AYlm
0l2+85UAWqe3inMpZw8wnRgIEl1ezjUWqDghRhdTc9ROMWjeOAPiEUaEstmdW6xmUrPHhhzfSvNC
cDOi3ZT/eI0MGmBgdhVwrfmWs5QHPzaatVfDPY1at9dGwEb1n1Tl7bKkBf/ZGd8peX/yfoyYHYbh
oSf4mNe/WBMrrCyR/W3ZKlULRhMdjIPRgMXWrNqwdk+/Ada8Wcx7/ECME5mx3cNlErVyRAWLJO+a
lXeKjuSXt1AuJpjFAZds/FJTd5bNYqqabfjT4KA+RPX6T3p9Z/DcO+/mDPyBYFXkX7qP4NT/DerP
QRfucmTWqA/x1guslOlrD7YL5QtfEwFnSuep000RM2X8aLULwVy3PmjQKrFToXeAMmefxsB6oqUR
svwMfXDqNe741F2PY9nqGn2sBI5OMMVnvkirJPRBJ4hDxfi1SBMzfQJZ7ZZ65AG2Nt28icFzM1ny
K50qZoQ02QAlrCtToONJdEsjb8dJiyDHpo2x8APLjWx7Qa/pmvXmeBz+cxxW9ez+U6ypiZvffKh3
f70SBupvt/G6fMbvppbewFXXuwEoIl994DrpfkD7dbtBu9aA9mRT+ExDYh0LyYb6fQD9O2XBvKKP
hSZdf8NYsLg4lOP2vyYaCMRX96ufpa9dACsx0tqYX/F3RNj3NABUktuepkvWzjnHVeOxbZYiROHZ
IbuGBxFPajW4pIpIhzFIhU8/lM01cJNws7Euk22nhW98/HD6KpPRVYX7FUTd8+hLHHQsSWZtzR9O
mO1VfXs81N7GK6mecbsrSNgdaFBxifPloRzEXQhz/hGhFdENEFD6XA2VPuJfhAc1qD8OD2IQnTpQ
BmL2apKOF4AoMorZusZFKzKQDO5AfdAGNeTWAEsvHS8Qn16nmhD199+RSxQlHRSNi0rgRWxxz3Hd
QV/cQQsyKo/qFXI1uABqE90I7JQJCkbD4dkDEBHeExQSaPpFta8DtlMl0/OCLWd3yLzZ/feZDvwq
+RGa0fT6lYQ1NrJh0wxv3dVHfZJx/og3pWaMZDsGQXwGBudaYXBmG7OTy+DGnIfPxkk3EyB75YsD
9gbzUpMqWg1dxkiTInjSnb+BQtNbfbFNnT58LAdfiQzNrWnR+Jl/v0dswkr86VRMwqI6teGAveII
yEzpF3497mJpaTPI/Rbi8r63D68LcDUAvaO309BEargArve6PLvcbhf7Odxjt8WR2xQLClCCZFqk
7WSYW2Fb+PuGp4kaMVwiUbuPMt6W4r2FHQ0qd/ben7t94VSYEhkJMCNcpKdrztXt+a/JuGveqSR2
6Q0YPhN8vgN2SdKbV/rWrL/phKiycn8uuJI9D0p6KcHBFiAXJqUCpiOM0hvBbpjVM/CF6NMeh6gg
CDMiLf0AkxjUgp2fXsmHHgngGXTXx2ADn6WG6Y6qvwHU2fGr6kmdSsmWvLW3MMeftZ0lzKMBalf7
MwoNj6PlHmnWYE2rnslZEDNxpcWlzs2InvcmiXXuAPMwWE69Bgw=
`protect end_protected
