-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nsdAhzm+HwcxLVDnwSkIJwIAc8owT/tDXS48nPwDZcw/h+RAOleqPlC4sBCwukMw3vt5uJlG3ktB
HMv9Cje9hqQrIJ5tbemmPrZHEnNleSelToe8q4N3SVLdtkTF63MaZUWnTjsUpQrH4Z8JqMWT9+wc
L4dHZFq8ov/rYTyy3E4eTmHE0pFYGqSY6ygHjfifI466orAbpM0W+UsFHX4JItPw/W/FxS4CZuiR
ptRNEgok3+G0xE9DNwP3uJBpN+yt5IIJAcoeyZu4F/L30cSZgCQxh6an120VQXLU/02xJpU8hUXa
2264PjGv2/MsxEjteNBJopNO53N3TzJf3LHscw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
rSJu1LRRTi7Dnfh/4OlmpHRyDvmQV07hwWnJKeDFsQxtruZ+xToeV4iVKpw1HDqosIWq5zTJ+ri6
9Pj5+HyUk52gES6Q/dOjROpZacgH13UItr0l3dQnEwcObnxXFaPLrW1WFvVw11DtYgeLAejwWk0c
8GvCBovqeYRAyV6i6nxYeikuVEcCvEMeryx9xoW1tO1NhbkFhr36zP21eJyPof05dq+sFVrwyH2k
qP5HL4h9/F7Olei+WlKQBzbChGWOgkc5dKdqrGpJUaH/4pHmCMlfwgzOZYDuArXqHBuWV4MtjlBO
Bu9T4cdiiRXgZO82zKHsy3URYKW12gMq3JGnEo78T81k1NUyPKggi4IqaKeU4aCPfCW3tthTuKnU
LNXGFrpnMM6wU/+YnPR/UNmgbAFINsPmksi1ezBniU4UC5C+qWU/7JaIZ0NvpHorbJgCglF2GTH6
NTeZjNcf8m54l8uwcjzALw5HfjDkLly69Z+M6f+SIAhMvqF3VrYEw0wyqdc4KelVvHqzREBVEhrL
eHRllEL9KGIlmbgHftk8hp7b+u3S8qfAuslvq7VMZK3zDuP0izPRm8ZadBKJfWrH++zdBOaF8tCE
rornZEt+xYlGPu9qm3acGpOysBMQ3alYUsTQtwbl2+Q3yH6cen+o9KUsH85/aJ6eRwGw2r1u8Rk8
jg55IcVU+9Oovn+NzAJxPvEUzpOh31c7Nhcwj1D3zUFcGQOCGn/DHWm3pcTv579JqN3lVqqGXIaJ
J9EEcy+PSjGEM+y+mcC8KtMmuK2+lHfeuWD+CHH3SMW/R8gi9V+wygV8eulG7y+vvPXFr8mbPxkK
oaOqBakOoij0zi/TnOJSKoiwEzRBzRDiz+rKLnLm5QW8BK4EBXyOUDYgN514XLBCq7aG8sW0kbqQ
CmoJVASVA/aGF6NOoKJ8rTHBq8x+F83bIQS6yF0KhknieUOp2Cmg8/mjp0cdrMzpL9pfK6Ul7+WI
+t9XydWWnk686/fnE61OaGlPLL02uBhyHi/HazsRFhu0ASQr5Y0kNkWxmBZ2iN1GrljZug5AV8l0
KNqn+0/0zaIH3YOx3jo0YpSunZdzBDdWUsqwKNrSMiqnq2UzfCguWQIrj+qJy9GghM5XPA7A/EaQ
na7Se1hqRDONdJL4NEfesCOAhcOTT6m808rSTUF3OrVg/QRXpeNOXhUUI9xJXIJong9vIH4KbgU+
ZvdLMMHRVkL/rx8eWh/6k/L6SmBcYCbg8xlblSGITtUo7fZ8xn+Im0GqWFkkpNfdE12HxKKfqZQ4
DPMbZafn4sa3jAR29lLrtAQOpRHsy5cOjedoZpFcLRa2c5zRqtPkvus7hVCEGzmW9rQsx6UsZexd
aFmcIABNxTUQ5KRSHv3HDvJAodiHNWXhRM1j1+njus4nCmw+tA5qLojAnB82q0p5SRgV/KH8Ljyh
ZvaO6UtiOWE2NxpYXbJQRx5gKA7cOe2TN2zHFJATJQHnET7jCsd4nJQtLLZqTEbZVkA56KzJ5Vch
BOmq3IVe4YjTf/j3Fu8S66siXSvn+StUR3q5OUW1p2tifoo8E7ZJzTa5/CxuAf9eq6ou9575hf59
TbNcohwxfFSyrZUBHMjAuOwMT0PDKrSelNot2Aj8gK0e5FUdjMZ0DrGU/w05Fv8B684KGse3JeDG
Wr4TnB5HRyYwmqoHlOWl5l71yYOTIaIvmNCnRd9nMqNFjZ4x+GuKalhzBGn9+WZl+V9UA32Fu4cF
eAddl6F0Df3PikV7v0tGz1OKP0h1u/wIStHBKGZsy3/rd0hyjxmwy04dlQ89bqiN0aLi3u5Guh8G
fYb0hKef0uaBmchO/fEV3tDI5VuBkVoIx9ifs4cF1FDy6EVuhAuK8XCITVPSjBOH9Tb8fwdoJjKM
IzgsrhXGDsEQvqGzA5Xc7aI6FTLDamN5XDl0doHNAmKbAzwEwi2Y0CGhN9/dFPec5U4TtBaKpsM/
pfWsqrkTmSXYoRpKs3HZtKyLQtmOOx4q1OtKRG+2DXF9tA0psX9rm0uKZyWWM3XfBK8BW4pl41HC
SeEMl5wLoRgRl7FD8R11nm1ebXvJbbrW3qX5wlPAa6jULafxZVKIdZ4kf5L7dhlqrcf+4PhQ5QxI
TvUShapa9B6H9j6lvO9lwGaFRbwsTEn89UmMTsclWIiEbkPmroA4Dx3RUAbqdYNK6GRnaji77nUR
I7fAr50Q5b65Nmx0Pevy2rQPSLogLYHnRmxRYep2N3kdlriezSR17b+hLpmgIDOjZ+z2gJ8awrHn
Fewks5+jsQ66sU9OqQNzIKopVRyX8lceqyuAkEMY/UZa0AWGJS4pvRLUZT3+otQydzEoltWAm5xW
KhibquSInIQqmuHeh6pe2QxVA/E9Zne64r/G4Es8pd+58yhZ1VULqmzh+2057LTBLgDB2FGywGux
Bb7LKGwVsyBM5jHtC1bSlus8suLhq6inNfamr49Ic/flhL9iabraKZlBw9N2Wt3IFJ+wLqPF+Ha3
WTg29teO5r1qIX+/MvrOR2KPK+NGG6w7V7lEqPf7R1SPgAMsXczyAoj5ybp24Pa5FJ+IXq2CmIwv
pH/y/D6CUlJDw7On9NVLRlgJMLRVuxV8vldnXdB8+ze3FoplhH+p7QDp/Y3IbXrKPl3DyHpuczoj
JUhxdn4bCum1NDFz7VSS3HiiXkldTiPqUAEQc0AqMG817A+QGX7RaE68naOdfQ2GZvOG4KE41gY6
1lwbqjUOMyZGV4t6P1FYNQbzUogvdOGU3Ll7ROldjeYHnIm6cv99fHgijf+gXmuQ7RQxyKr5qJC9
Asfwq3xNOt5M/09XqVkw49AGR2LfiAt2JlS6R6dTawB+ke1l1mnpZIIZ1vbY9FFD1+ysM0RwhfzH
byauRX5TqDPFSp7oCNF/xZAOxb5S0VgrqWiTprUUwQ1kB+fFZEyHTAQAK3oZzC12dQYnkMZxEohU
iISX8RHMlLpjgkgAE/vBIljZTKhaIRlQYFKGlJlvNgpe7ZyOErNZeivr+3ZpCOIo07GhDjobyVsc
zDdjEavSsbfoIaceL4mcvCXYvLZ36mzCV6dcVNo6D7DXPw9u2vF73lzYENQzdViezvUH/lVMjzJ1
whW0bQBohKj55FplHAmZkJTFzwKHlnpikEJo30E9IHM5xsOoqEBrkidWP7T2HlIkiW3gt5qcVy05
nLiy5JQpUpedUX35g0nTnCslQDkrxwZVnBjClhrAgQwJVz9D7R4seCiI3kriV4lylyQ4mo6Gj6Ne
XdsuQebYsd6V2n3w4Lt6lkC8yzEHUJe9d809l6ETAaYEXWkmW91znQMzQd7X1vuaVwQfhIswT6m8
3cykk0HXquSQCVMBVL4ngR2T9+3bgdCCNjLx7PVh4joJs/Dh4M+iYdWW/IgIqu9bGHKm9B86COwu
HfvOQb/yccod6UBPTdFbux074uvK0apEdouLjdryUmhuEpVcXimovBw0NFVojr8F8v9oNZdyQQir
KUhW0nB15IZjhqfLaRDbwIefEPWAb6G9W73W87pGgDzIHmRHF+MoSOlLWm3SlAgIoXLYCG0iQH3j
WeTpiDWVqdPqQjbdJ7xFgJPqRw2es9QtzxuowYdFm/DZNyWl/Qutmk6raP6dAjBj9yRTaCSOT2I/
qeuwvWrswn6LoFTO+pzC3IS7uBt1kiyRXjhdJnVxVYDvhG3cvlDjQVsTS6z7qPkY3vdIMqRXpdUe
X3KympfhVk1Po9bQ9EQlrkbkR29u5XAoR78K88vNSmEoPSL5NIiUXOtIHpRZcnZJUhGgwIiY4Z+M
xZC74ImtejLAcl05RQTU9gCtFCLOsD36AyMJ+o9E8dWf29HHimhsd5haO2q/Kv8fXTYFSfNA+tAP
+lOWJdu9H7Du6Vgch6rwFzcdznP3b1OjFIvJ0SC3hoR7PjuRjgMik8y6aNW0spnRlycDy8ac0SJT
dUXDpe3+7tFCudxdySPsiQrpDmbaCFd/MfI6826ZOa7xMY0Zmcxj6RwaXodAnQH3SosAzIJ6eRoj
9d7H0u8xOcyusm+q2lg03qD4z1Hm0biav/BJW7l/KSagmaP85+46W8E2rE9/6fbg33/s3AFLYqcx
aoSPi9bWKtmbuDNjwTTvD01pWKFDl9bfF32twm0gaZZp5scb8Xh4sVk9GEsdgUxoSZ+NfXB0OLXY
CDqvbs78pCAdwkjqrPPby3/CNgSTFW984g1uKCZ8DsgA2QqZ46DQQLQ9PmFsioCVMCvgJ5/kIDXY
53Tb+K1nh9X9ZOQD5mLQeOdOI21wqkMTCCiNzofotTjb8exug1hiiuFFGfSRaGORnL/vlN+XZeDl
pfBtwwq+IXy+LeYEJs1FqMnc+fiYsfIXBNzb/AzCe4jANgT1BUj8NA2Sdk1ok6OFhHt2+9qljL8n
hZ9KpW65G+4FnPxKlLOB8AFJooTbB0RRRnmkPajD+NHFHuI/b4VqyRmfk1JpuIgRFHH6Qneiz5xA
5ufZ0vpi7ouzbKej9vCGOGv/97F2UYTWxeuMTAxxRoO9+qpHZK8kCEkr5OHzDADuMqambsyivN+h
K6hKav0CInFwt0YVxeX6+upAuPHt+dyKuoO++uugVS0RB4zhi5ijiYb+MWbyyPSkjuEHbaW9jg1X
0APOtB+/s92pq1MA4L0xn5Q+/OE/sri9aCZ3s1v3wn8NiwtjjJhWZcfQGxe9EP7x6eBMpUhBEdiO
cICX+CYJ1Rmt9GQrK8uuyNNt/+Bu2ar5qXcOLsXroj8GmW2k1cQAJd0XuVRNzVGkmEfeLpouGhUV
TnooljRWnj4fA7C1gYKZ+GKefHZyn5Idu/RXP06f9b8J1TLuDauZKnHTinEx7cVxRkn/aOeNfRSx
9d3dFZQ8W3ZvYp6COWDOI4nRebZGeKMoRhZIutvaFyq//JyX0jTtnHihwpvRhZ6GsYl8mQgLY7iC
PzSRKZHT6tVbPuFrQx9Phqm5oY+NyrgL7ggVopELkGMbMyTJvs7AmlhmGTKGU5Uo/C0ajHDF7F/J
fuqVBWjxdD8SYs59pWyFqnRJze/8+aOBwLOj3fsfvVnYPd5nquIDGZxlzUxDUbbTr74rcqjNss8L
G0xB+GMwhRCqz7S+JeZAvohxxIoc8yaGgzZH47sLdLCPc2lV4JW+cXPeWYqlGeyret1DTqd3tSo3
KozCAbqG/qBXJJzJH3MZnvqh649itckHoO7aHGTBEmBlgJKy4aH/Mn+uM1KJFyLEDHqA5kPou1fO
Ft7SaoU48uyLNDZ2ml1AC9SpD3S+NHc2Oht/O3+9n99pRBAnT0Xqhw0KS7r7LeKPJ9dN7hQ10OfN
M3Zvgx9PZ5IU0O5Gha4+VbCdOhs4UnIhd14HTZioZfmfEK+xK9iFzxXcqkDz7MUun8Pm/TF3RHVR
NKUscyqrdTdNTJJqZ/9aI6/ZvU73SqgyN3gkEPqsBpoOmSYW+ChkORWRBEJeQYoClD83zCkS39/z
1N/IzFpzV5rxhj4OO1KgWSthhRfh8PudMUO0EsJG6KWqO55s+A3bKld8KcTV+9cq9jUvFn38h/xW
KVrGk/VeFOxgCBAS3SMUpHNDUoMm45aedb6KuQTGVrUXagzTwuOMsrrv9eVxSI1lwSTJmH5OuFXt
9+lPX+WkmS8M6dE1jG9ghpXnX0W3yKAwjxQtM5/yW0y+jAzlX7dxKIL8kGT4tDhESWvJZLkWIHrh
Au64Xsif5+0ayvo08J0UcOrIfydQOiGVc4A1n/Se9rkhd2Arc9e3sRrK2CHNG7ChHJW7LfmdtaZs
IRafnEW+wTslWS5AgTe9Pr+OkEz+A1YLrcH1qR63MuoB8jPyFnvraGJ/c1k1aSbcM0rVvRGvmEVu
q8hkxj35qGeo0beLUdVIeHr5s0vBF7bt5Uodz/SdQAPx8ss6vNPkgD+YpT/GNuTndvWrhX0MnNxm
C+hmXqgTvQ4shmP5LTLk91s2Ow5PZ3IZXFD8r2GiyUUoeNmTy7GgXbNM6V0DDLLPiX8q/e2zYHDB
Dn/zlQG2JSHkJOzxNxSdS8kyyADCTRI/Rbup74bRqn1m2GUst4qjvFs7yPNCEc52S5Ztm4qS9dxM
XL4JtNK932611GwHWXJjQOXg8DUkM4Y87YOd9ZwoWLdt5z0gdCS+3BXtkzurIS/r5O/BwGDqP0tE
JUa80H9Ou52sqw3SaupytooMs4F3oGRxT0l7TTPjhpFIx40pW6Lx0XhDbI4rLRY1kCI7sSKnkMdJ
u65MZdZ7Iqa7vrqFLCQbR0jlmUWlVkZbz0UzlrrqmigTGohmoBRH8+rso395hr3JKVMFD3ZIBKzg
0sLXoKdorEVmNZcva9OxrsE3Qrt7cVTmMO9+bSZ4ck+182IrRfV11p6kntM90iiuQd7DdTjpwS24
tP0qLPJGLXd0vN0aTRYJ5eji8AiN/B0GntNQgwBtsQe/ATzQuj/tQdqm5MhzNdFCiE/y/neHvA2w
dpKS8/bXxdK1N1VAjclgMSgnxOUs3mOFlcyldm+15wN55NlL99SWp/LJt3EtAUqULPbbaY/Sj+gT
pITZDI8cfs1RJuuw0iLHDUkrpxBFOKhkESag9hLtn4S4bgul6UUZUMCvRgfav4NSZa/Hsj4jiYJy
/gra/TxNkTvlRT7+UcBLVIYqAfznnoKR2B79JoXnFsano+D5Iy9J9NR3JxsHg7uaNGVOv/SnbLOR
HiofRGNcZWKV+idaMtRhCSYnDNg5p7Whjy5bUrAP/DoqGtmlRLpf1ACFmnKwVVu+P6zzZfg4mJ2Z
2I/V/Ps3P+ydD3TV6htTxjzqJfhGJ2b4xT6rN5eKWBR/LsBIgwPe5eBhdyPgKzuwIWgMSDm9DrAN
Rzdc4QMAwWrpVOQ+BRdfftZx1UDcv2NRKgW4CnNlsSN/pZ8Pn/u/7Me8DkJUFfSW3au9UXoJzeYk
wMI9rTvDUncF90e7tlwWSemyg9Y2FBidSQMJhBc7S24iLexsQrbrpXN/2AIbyfPbV4kMz8e70F6C
86dkET7lce9R0WQ9LcH4zn7Wx0TU/lIL7kkUM8l440TJICbCNPBHlKFJlWCqk3mHUnlO2/gV2ZJy
Hvs+M8uap8quvlMazunzlHP7lsGvjktyN5gocnlr4jHE6+tzarnzzD+4hf++aKusH4cjWd/wb5Sd
VikyC0KVHYK5ngl+GQmUGM/mYDeCBWAQS0nCrda35OZNQQ/xZXGPT9xtccJqndzf1A78iSir/+wP
vqmd0rxziT8SMpzJQ5XduiSI8jaLUnbj7dR+z2tntlwsWVoi0jQtrFzwiigA6W/oPRLxpZ5dFI8p
anjff1GZl/XUMbL7NrtAG+npSlQt52nLU7Lsh2HB5J3UC0ObDTwpR8QaJc8xKQ4jvhe30y3DdKZ7
kIqlfC1sdhkW0zYHr047m0R9IKdIULWowEMwU+HzYKQGK7x23Vd24ajVCfWQgIlfTs/pgx4V83K7
JC8eGcMgEqdtsv9zsJ2o3yRWdfHeGW2VUEJpKwR7aQnLAm0iteH5mIPXBJFsyIkJ/Z4HktA0/I2G
uX10dbCdlq5Db7EilqYLNGSU4tdq6VgujQ/C7J2tqcnoMol42XkP4JK3iDi00KF4FaKV8eq8KNjm
uhV3yOwrq1kiCr1cWRzP4NH1YZWpZ8ZPgEn4Cus/aPCrzniwLv5HnlG66+4f8YiJ2LN/0CA+OeO/
YWRwAtoqbJ2G9+eRYLY8RivVKup+y5EFUGfGJmpH9ATWD6OFE0JwofY6oRhE7WBYr3v1k2qR/tU4
g6MYxHlAbtDxRsK2Ut4grMw+p0f/39FKLzFQjcWq42yHIKQD61Dbd8VDs/MxLRvGozV+lgxiYrWW
0PHAn8anh2+Y6bA8ljG/XwXXyVAidgkCHRNO6b8ipaRClFNLd4CEG2g/tv3eb0j+OM/MKun4llak
0GJq8BJ3ThMuBYPHH1u5EgC01MBfcBtT1Sqv2RSpD6tekH/MrOPx9NKCaxdjTc/g96KAwEojahHm
sc47RZWbeclIHZg+C3sVSl6gJYiWw/MbHQItWllWzCLUVf4avzqnmI+qbdREawCG5KTy3MZ++k+H
8j7kBx/MhyYrUNgkAqIfqxrP3OA2x/VQd2Uw6Yz/VYpWeibGSXjx041Xf2cmfiwpPj8l947LedC7
gmHgMc/rhiiE48RwgGPpp2O4CtJI7kUcqUSsuIa9tJSRwx2hEmllCxepzSfy5kMwOBNDxrjqdZAQ
oC+N+d+enVv0PuTdA11p3Tmmv8MldpC4Tmt0JQ+LjYh/PdGtcoyIPoWxLpwUPv8IOCGuDe71JXPv
OIFWdi1+lfdFvQnU3QoBrycX1nRuz6LOXw0MLVxUPoxVbnvx8+CFTzj5iipPGZ2zNSF9zuRKmmlR
Qad4i8ppeKtsNh4CYM16WmVBHGxBcA9sWibgmS4F576DoGLEd5dyY1zpUWLW24eJMa4gRNPA1rHA
j1QEDmSKqzY6pKgsH31ps1stJpLwAkUzjnIxVRNdAyYwodq+NglTMj1HRPj23GiBYu2i2s0SiXP9
oyb/RGLQKEfLRuWyPwaJWgYGGLU9iNy6dNyPHp29SFEV2wZvGGO2Ds6K9FkyZbBJR9BeqVtOrv8U
+ehhhl+ZF0EIMHNqYWFNfYV6TJF9HvStu42YKT1kJxQTsYM1TeZ2/Nb9LBTAn0GjBwGrWN+mwzzp
7TzHk5aUN5nF/XFZhfgJ9PtFtH9uV2BF6Tyw+ZQWnc7RL+4R6xbK8bwVmCTSKIYtpW14K24Be6c3
+k3uWY6lQGwvXEsjmTcXP5f9wEw/yFq9kHzMTw1IlhpBiMbas7001pKMCI7Ydu8pfZlsanbxDgSf
TCh6WqHaU6I2uc352yxHhRJPRHSPx+TPczv2/M019h55Z8Pr3/t6rLhLKyCna/ESkJzgoa5zzV2i
uY8ksh9v3JeVDoQe4Dqt6VdJscJ+HyyaJk03v+Pk+p7McFkFTK5CNZrfhkPSoWq3RkaBqLtp0HhA
oZo9wKOHzZh+JhMIxH72AS/c3+EUvZ1ov2LGOcVF8uDUDey2kZNX5+T0jnMMW3qM4GgcIL8tms84
28DXiyK4dZPQrbI4+pJF4bn/iHqb852V00MkzWHjwPdPVRLG2d3tZCc1rS0jSAKFNJ5s2FXOnp9R
XkqDlVrODefhKmPyfpC3EskwCS3/PbLkdKEK9yg+Va6ThxtfvhWi+T8z4FJxmfRnD/1nOm7cSa4A
GqOXTe3SXaPyzGTNuKXTmwGWMLl+sohWhp+6LV2mpOYkTu7tVj1Yzk2IsML7ltj1s43GbINU/Ice
PYByComCS1mZUU1jMxl5QSCisELkFJGP0Zoem2nKsajVrqSy81dPbEtK8SRtYFFwV1yZCW6NAN09
GsDneO+V3bmGSxSAaWyGnxC8BGaRuaIuCg0L/fC7qfTpXvqRtrzREF1fqAHMgaKDtdFk7dxOpROG
7tftojGXI9pCIURhtOyuWfzazp0kY+e39cj3SzUFoWFTEwbvHPvEMNv9oWuHwCeNvTHaQNBglhyn
X2JJShABIKgydj6eWeaCeGlLBxqXmd9zCo8Au68qQZu4k38a+TNDNghpm9zDVyWFbV+56V+KOi8b
qV5J5QvA5XsglT1xEpJSjgRQcdJO4gMTst4/jEzgba1KH9qrCROOUf42ySWTynigNj4Vmm7kPuJL
za2jBawySPUiKcW1hfJTNlN4tM6T5AaBRKSVjB7+3+KWPYp6ciDm/HNHAw7ljpEOy006XaUrPMtu
BXqEr4EHdmF1hmK3VLskyEHCmWOW9QHr8p1a7uypRcJwRvYiFcFJKQss8IzdoJ5ZMpDw7alAlNzM
zk98CbgfYnTNoHkEgpfNmLicdBieuWex+y+vU/0XHdg9Rnogi2fmR/gRQi1RF88dQ5T8N3/Ep7Lf
SpOErgML4EOyDeyAmuf6kRjcq4ArIkLnwYd/GqtLGHumEfoOSwwSfUOsP0SzSuVED04djSo7MSNK
Oatvpd4eibO6nPp0Ql0OUCdRFOaGGrjwmVR1hsiQiRHVKfFCzmefXec6cAKlITAhrr2FtG9SkJ8X
oi5UIS4Vu/8VIL97pomD/byQvrVEz67xOP41oZKMbt6sLafA+VjdwFWM884IqwuXJle2DDEUOFcS
2V6b18Z+y1ihpq+sHhBsrHkgah5xSMrP9GGxARYLVB9+hGwR45+c8yM0VymrpzHLmXFhSpBYQqJr
cGq1JOG5exNFimkdSe/0a0GN4mJufLtCG7rONDLiPuIsqwSRGSl/CvdgK0Z5TWCXxMzbgL0M0yIU
t2D65D2g9fN+iqCfGaHrKpz73gJhbIqOKpCTuTSDqt2nltKak3hyBIeg3uD6OS3UCh+wG6DOL2d2
4Lufj980bd7Wdo1brnVK5n0+lfPAUJX1Efnp4g93CTsCrdMq4PfcYlYA3ANcnKnMl0BUoNg7Lrvp
Bwzj258QvPPfh47C7sJvhDm3KhdLp6z9OJm/k7e4WhvM56iqFor1+F6f9LimqK3Z+XkZrBw5Lxao
M3rlVjvyaZH4uQrZTVs3aRIruPM2aBDjvqDevK3Q+daTSP9r4j72as+6pf2WOn66BjzhoYIY16Yv
MtAVTNp/1gzt4OcEECFPW1pqjsL8AfyDmCa6l9Kjj1gAL71gu7x9YV0AefK74o48m+EhLhfz/FTR
yPDcxz1SaBfoB+W/2rAW3ctSoxeSqcer5TP5UfWg03CX+JNmy5wV/VdIkrKMOPTnlnUr0M9p8eEL
Rm+O+T1QTV7ESVBwiIQfVcINS5sapsczz04sHyPng5MkB8tWtU8wVCCb60kl/AprZw4g+GmImbLU
O8Yw2yBl8wLBapL35lso1GQ0ZMjBpzvPQu+wBqdZkPFnVt+R/n8vikHcnIpVXql0l/Plbv7GyMKP
tiAX7oqEvhslv2MpChd6U/TANBCxpPUoxaZ1JbYXdX7Xsc3PQod2y9JDYPUWqW5PwGdSksasR2tY
pKWMECaSDxKfjTzuW6+FDMdkSFR6oGeKsmLerr3+mzgeI8G2N8v735ViNmvxZx8zTcVQE+qU+fmG
uuAnSL99ZwMN5/TdSWQ5xKw90vgjypPPXJ0HPI7fEVKGOxCWDrJI2SnE/cGuM2AQgNhLaFvJBf/i
fWNxbya9Xz+qJhlQzqaXLc0iS3hvDpHUVXzEMTqDIyESC6V58fikGt+la+j+8144FPTF1zCSyV80
n1Ap+Ozo7qpTRMphRH0fPeR8b8T6lfKho9YkDOhhfEXoT6dQYJNpsHOfpz8kJtpLUCgZgFn8UTyU
XxlwfZupONXey4WnvkXxjSw5zM67qi5orR3W92B047TtIrogl0upo3knEhbXYrQKJvEyNdaxyO/C
3KeUEBnwdZlpbmouHtEZ/QtpK3ZDkSg+4lkzU77y6nksjTDbaPtU4PT5mBAdf0dtsJW8tWEWG6D/
U3csEzadkW908QnNCZnxf04EwZE9dTDfBr504xFnTylPI6V++HT2NtC3vTM27AHnViPCT5V9Jcfi
d+6t027EeuUEdfM8s+8ZEnPY8QbJnlcJc7OK0znPrBE1NCdDd28iVtGE1DCJninfQGJ8r7voNilB
JcWSgo2/yZBUYksFpKbt0Rw+PD+hAwD3AZH2XICWrVQEc4bbTYyyiqExrkOReiiyafLmJ8BGC2Nv
YI8NZeRCEiw/ONtkyxYDTsTKGCxjfZaNrlLbDvX3AtKPBiwxOIDiRiIXf1oSxLVkL/ubvlmf7geB
7CMD7ZxP5lUA2xv/vrkVBnYQCoUQd9DdMg7aZqvth0Zq4QsuX0IiVfV2huLX0aQSY9+Qmo6jmhZ3
Q2UZdWmiPwRvDDnCaZdRltUcmLdD/kcpjW1d3fmC8bobVq1eXiW4jGwXBKIidJdSOt/m8RVKGnPH
8k7vc0jcQDvID5yhKb7Dc9wBaGmzBEoIVCw1VJln5/9jH1XxbgoRhrvP22tBD+cD7oRR8g8vnZdH
QDVRA9gSUNRCd/oF78r3mKZK3XbVjcK0gnbDIh/Ac2TJFRq8z19mRmivABw57aDAuwnBqnQwxi9S
IalxDSvu9oXsMd4JBjYXtNCYaJNPNIlhjoh0HiUFtStYXw5tNwu8iLx9hOk9zraPo6CdF0QdZhHJ
PC7VgXXWOTF4/TpbVyHJxFReXhebsaAwUx+/2sERaCArBiPuZxz1hmAljWKR+c/1X2lFkFU27oL5
8N6M+7eP6Mt/qvVljtqai3ALQHwg2M+AuLFlEn2U380bjDoG3gElS0wTPa3ltvr3M5tvkd68j48S
aKny2Gk+s4qSVgMfVj8vGeznswTNblnPsZiQTZS5mEUjUZABIUO8015WZddy0Q1RE+SOc0DGcUWz
VWh//KkviQjlLf1yI0gJIt2jHV3nHBJYaZCVreja/Y48e1P1EoT2MCJKPiVILEse8Jz18fkvohPV
uxTdcto7QmzuFO7G18AQPDOwsNpryFL6iYHNiSJNphURPwiA5GZZ0O529pkeRj9xbvZnDf8JQm16
NaZUjHMwilT7w6bANYeFBYf04ZGuTmRsF/eiXgR85leDjZP9NT6QRlWXjbUTxLVlCwFht/dYsIqE
ccoqqgLiGoMvr3ZTfkeGAs5bD5e2q4m5s2+nANERa8ad/hW+bbD9wIiuJrf6IIR10pocXjDBbumM
Uq2T+X3Z/B5yENPne5s5XJ1JnmhEfClFfHtJdXqa8pgGVmTOTaCtLU/Pft2bq/4t8e5x+4rU8m8k
pO/bJRojOdw7wv8dlmCmtw5sdEw5EcHn8eiKJCNiL0te+3A87g+D+Ta3wl/M1zwJQfMPI2b+bv/d
CR0QFQTQPNT4lWQDr8aQQuAq5ECU41BqMtY6SKXpsLN+n7MfD89UestxxV/OOJQP74PfDXFuQXGm
ZXvNRUr2bHfcbU9aZlOCjrYacMi3eY72LEEAzrzmiMnWgyPKcUT02QlcgfR0bIowl+P3IHs/tYvO
hbpHIIoxwGI2PyrxL1trugkNbND+/EApry5u+R4l64yTh3MDKtFolOwrx/086eAqHqMmVOhOjvir
PyI1rwQAH5Miu/1hgBEY1iU7/BdJoGPb7BrDoLctgqjilb3jHEHtaNWtdsrDudPdMSu9oT/pA3F/
O59wslH7Fxd77ingfwMaGJy31zyNuB9UCO6TWTRf7B7Emy0Jqe97ed8KYEu+aSmRCMaZkfhTXPKT
DkPB1GX0QSXV4hACzcnLepAMldamRARfszw+JA3zApSbmwz5SsgFjz3ZcWvoNOeJcKwQBV7GKReb
gq8zw+sADxPJxZoBmy1dkWtwK1SzUH6aaMLs0M/Uwt4GIBCR44u7Lu3D+9SDbRRXjEFL+x4Secy/
Br4R+jWF/5FRSJ3z5LGj9iMlNBj6NXBsIijPgFy1n8ECFS4Tari6+aEvUmyB0gLIDrhynzY+wdSU
m9OStHCvx0Bou22i8depdDCnk6HHZCuHmmNb3r36SJ/SiLc7RjyfRyl8WHIF5I66WIAQfHDzWdNO
hO7rIjsEBhMVHC1VDBag0NCcq/DMSaxGE/w4xXyQfln7k+zx47gmr3Y/0wfe9GeWs657c+O5qSig
kKD4kkQHhoEdn3ABVjCoEPGoAP8LBpANfrcyeJpE6KWvkbG7QugQeKcMLFsD0SVCB1G8SBrCavJX
dXXiberldI27S2DTM2yB5TzmRYiVqOI1v0trxbdpXTUEr0+/lxeSebr6YB8cET+CmJNaigpTQ5xE
8Plq85QnhRt1uFVkwfmeDan8nnE0XLRnKR9SVPp1EcvBXqxIg9x9Wr8c3vADm9wWHZ7U2zuGV4Q5
+96oLxAbMdomgytqKskiC9L82TfeN283mjLtdDzTLWQiFuvZ0YHJVUnZXK6pmR5gXuh2VvUGUqHj
VhaD9+Ls8cU7iOQdSi3YcJRG6XZZ9xLq0nmDofCSdVzkubRueiZ4p6hI5TOuVCFbTjAgx8oE1PdB
IouH+4Z7MPlcJNLJlOIW+ZCCLSvRw+qSFGyf01lM1+9/WOzn0IPk879/14zMC6PebDQZn9z44t3d
6uwJJ8Itoa27RpHPgdHL6qs5Py2od1oD/D9JIRYivEKqxSov/TU0VpYeL/Wyi5ic/eoAWPdZz5nv
BhqNltyXiIg/glVw4vI1p1HLlAixjJzBx+cVa3kUztxh3aOa3VOzgXz9tiTC16k4N+PnuLzbj9mM
ZsmWnyKiKBoIkldqamIoumUs33lL6wHfwoNd2HEbLZ7WZFwOon5ZhyR2Qv6rrOpRO561NfiLg4N5
V4d6U8HDuBMRjGAZh04MDoEDsymcb7iCcsrLmgEfLnDhexp6tJ/XaSml+Zc4uLcH2Y24TRHCjSBP
0AtccRCCBCTVC1yF1XiZL2y0zrP8nL8uyzAxxQRpgj1IvTIMwOL375L5uoLEo/tb4kzchtOEc0Lj
5VrcHZCstugny92l3kG1hLnMRQFWZM1DFpOxevDb2t4HOGb7KzBTzTfzVG3lvgKNhK2yyPrYqv4a
iSBKi/AT30Z7syzsvCKUh+4mRW8R7P7/fBT6Y97nHgQ7Fdm8zixOBhvmP/TUQNB3X9HYI6dCjemZ
ZCQ/VQGW9pRKKiDArA75QMn6pqVpJG7ouJtpRrx91B8WIT+K0bnPMx5AaPX3uww9MesM0GCb2uWr
jc98AdfJhJXk34yIkDEcjXlAUuyzF5WGLdfHnyWddqr6Gbm0WKJ0H/aoiqF3eaMcNR3PM8FoPChi
U32eu+MZFv+J5g0zUHFqEaDFrgkjIz5XRYap9en6+QTVw7l8tX1gUfCxb1o8yGtYPsGvMrRmcepb
r/K+LgkgyZjq4/tI3BbG/vS7JmroRKUN0VfDWc6dTMuqVqH3wZfW6qnlVIadmKMRkbGuT/SupwTY
zyU1AvUOhkJp+GSybdjOB5ZXnDyullCzlPaELMKDuflceyMliGDQSxqhDvPVoG9GW3+Pv5LgVwUv
9CoRDYwRsa74/PdzIU/kQ3oyHk9gf4RclXsJgRrpCGupXxkHRBIiAXWTJklQumWx2yMMA5Y0920K
crEKC6v4bDmvs0TTY/mzuJjGhfBmiMdVttyUsoMAVJCkD9citM45H8nHtycTs6bAr+KK+hArbyNi
AhiuDX5IG+/lRKvUUjsHEIEVuM3ay1fF3HWCxlTC8MlRRdDnZ+w9Ue1zkhG8WuzXg9fBgeVTOpaO
FIvtQUpQF7B/KAWgJlZUyeZdkOCT479Dlxduqf36uyQedB+vA/02ZXexiodem/8B3dzlORsgFYZZ
Zf08Ib751wxYvFRad9yhm62lW7YQDn4QHX4noKfVY6JFaGLZHHnuNH7AzaypXIxVS2gGs6vIOWVE
V0MtleHPlTEioVrazKNb3AeYbMKLWBxpFIg+RPOZ9VF5mWAbOq9ondJA9A8eBMRo7N849Snzx4Qm
ezkf9uUMaF5gTGr9Y5aBXh94E8zrZNiGLZ2mKR5ubwLzAuhgSY+B4r0Y5vJgT5WtnFIsoxYR7JWr
VsnEJkS3oyocNkPQ6af4DUFbAqtbLENMsE3agDKVR8ZK4UEUYz0vdvIKOUVfAym1EoB53jxiuiUE
1XVhLFyojvJ9V23vyFLpgJePhxivGU1z68l4gELtODKaKNm/MXRFEP2bVjaoyti46fP3V4/yXQPv
4FisAxVaW/NNXTuSOtXRXEQ+/PnL+KfZvaEGQ+/blsRBXGqWSNEecGNeu2GsN+JnXF9ixfwRJZ81
mKdu+6Rz8W8svKX/aqU8+1njFKjijTabe2Vyz0hUePVvmlbYmTwbNc1TCxYuimuKavDTlZl9wCF/
10Cv73zqwrQSgMqT8W+vh8vk6vTqvaxEbLGmlyQ3ThzOnQTEWjjbYCtrhXpttgektBxOd3Uu8Tiv
PsLSA1YwF2tsAjLdRRF047CVEAWFkMei5KhsZ0y2di+qOR3RdzdV3P78K08PpztkI59jk5JmQQXM
hBQ/1CstIdypK2meNPxpPHp/GkQvlBhC7rs/YPsNk7H/i1ezS1hMYplf8RRSBBURVzbmVAelXvFy
OhPIIcdxKhjGHrBsPaz9J7a6CXwd8OS86ucIEMq/cRH2jPgMv5bT8R62NBp7p2+xNb9u/LGcc2LI
XuvXiwwaL6fpjy0ab2DThsRUWtYjSO8Pe5B8Ofzp1hhfofz8lP3qr3T/oNE+7WIhvUe7UOmFzRC9
wnmbbPPszQps2NkH+UqQo8kuk4Z2cmGt8b0CVcs4TvO9qMoxBahWaD0MMCaV9mVs1hhsFr3SpBFS
j4tCCZl9b6m5SJNNBHrMo1PVHVOrvYh6bm04jC0i26VvK8yM2WaQBOMQ7w3w9aFeGIC35d68E8DJ
qCQqHoXNEY/L963tgTCV2Jp2X3u3KTgWDezMQhVYb/TBE1Izp9BQGtN87AIRKT8fMqvSmqWH0R3l
igidKONkpF4uvoFCvgKFmMLvgZnOnmnmi9E0TyO+55482rsSUlqpllkWkDl6aZ/jDK2vGCSsNDe1
83NHNaE07WbABOo08w3h5x+nTJ1o0QJT4Z0lNPxuwodpfSryox+UGGCu7Lxj+6AaaVY7g81lgBqP
lpVQcrUCn+yEsth5PBLFh9Ce55WzNGWYzOPYHyRxgE9BpW42nj3VCQkN4WyxAacCc6J17zBT9L3u
yu3DpzGvyvsgX+La+iLXGzL0i0EiRc7/WuYt7sdn7JXG1QA8Jr5PoUk6FtI4oHSg4dRffNSo9FW+
buZaYRSmyBN89zq3kDkth+vpROx+s19VwuwRRt4CAVZE1yDE4WQDjUhUPHvucqr8D66kz2zqIOT4
uifR9iR3Bt7c01HhE0Md7/Jju+bhKbsmyuzeUsfDqQHqX99eRaenY7XKhGBwB3Iwxnk8Q1k/oe1K
L9xMZsqTFByf9W6OGlRN7YRbde35awtRELm6Hj9+DWLkwRadVN2DIaxOq0Fseosb23tKizSg4Y70
y7hbnfH7V8cbzXcQrWNlQgGzSrUGQSpRbGmjkZxNRiiu+PbTDKe9jObp88gZjH/n2JYrAMkqM9ka
SWvorDRCrnqcZqTNbLcXPMlcMYCpIS9r2gDF0fvDvE02yyag0HLXYapfdBwEQDByNCPUE2C6VqcN
rWPIf/el6G1lFnoOF/DmO2nOB7Gr0lZ79ccXqV4pIgvc4QiP43TLmAlfkvSrJ/w7NOhJyKi2Aiim
2iMVBMT7mg2+cL1tq1oxvKTa1MeS5qkosSWMf8vg8Ht0IUqQuRsd4pN01jaDa7ocdW695Nz+4XYX
2LBhz8JN8XEu8CQBIOCv8eDCnJvploFynRUGR9ERKUXKpDcrciw6SjgOvrPnTez6lrfzmHPreSmn
7hDBM6naVslu0sHrksaLbhL2QLhuQZistRs2HITTMSQzgL6PwzWox8Pc1RWmMd6FfpgW9hyAHP+q
zHf2R7XC+9zNZaZgBshXrKroN0ldgjAuYNAgv8g5q4J/513kM8og1PVc2+EyBXOnDWllSeQV26Y/
ZZBWqua4WvjMQ5mlq55uTJYUVkpMV34LVVBFrKbIVcl8jpbeHPWFXE/0CoqR3TURNLU0HNDcoPpJ
gUkjTbfVlnpUN42LyxaXDXEwnHr333D0bf5Pzzc5YmQh3QTjqqgwJ7fyIwjwsvTb9xhS0OYXoKDP
f7IX6RmCKRaGL07MoCvLJcQFiPFyf7rCMBIWKfzEAhxk3527p9o/FXn9sH8izLVYlABGsgIAN+9b
bv7CxhmPOM3i5bTzdYhpdrUzjxSHAyAQB8zHf8x1TuCa6ZpuhqUISHKkgWbas/bo0y64THN5sw8I
VWWDmXEzch6IJy1RbrfeHUtdewVOGpLk7CyeZdMEuapL/RC+zZhdbe5jOJmSGQ0a+2K/nWxbmdoF
UcNfkwOdJHC7aQ6AsvlLgm6J/IfUr9kwbfFofS7+KH//TDLeQ58o5BqW0yWC/excRAvBRw29XUxl
3QNPTF/rbUx+1FrUpe4WKVtHU3iEPZUmUEmUbW7AoBh/SqhpnD0ywysvRIbQZU23YSXa3Ujzi6Gs
WuTxQgWaowHQbogC37OwlCD1QcOR+DsQ2TEODvDPW7QjStQh+dI7Tk19EssE60rdvWeOjyqi7ziF
AXXUk1zSxjUeHtVqXOUDB1I6T/xsmUBEXf3TIBe/i3HcHM26v+b1+gilu5HtpjN2jb3DUoIHI0Rd
Z1auWjdbE5IpPwZqqnvlrwu9+Ino5ZsK3cyT0ymgTPN7t05dL/cGM854JAYUyK8Lb4w4HppwzTel
vsxmZAHNolORjalqvBZXlhwUkY4Y/PZ1e+kw8R8otUmraDQLPrgaxmOa7RYmkss5uD2TDLc2Zo8u
JCirH7TET0PaX+IQFD0YlurgJCUfRL9FUZNiibAuO5d2fX/LakXNC4xupQe5bKL7ttRcCcqD5YKr
vB8YmYbvMzyG8MH2x2N2odI1i4aLS9v1gPRupZVtXInPOmf4M2FJqph6sRDtYwmqWaD5B+s+22Pa
06r1b37dlaOXTdcGbTxfr1hxs3W7jP7lZJdCBgkRO6Y4swnuzUTPix9B/m4nYEyGqn9I1Q+0lEUP
AEOO+DJiZwxSytQOyC1g4wCS5F1aBSCfnG/Mj12BBsX3DV3paD8BKhKzyaJpYauC0oj8lt+NhQ8k
dwYJlTceGxpCPGkeENsxn8sJiJCnQvqvdsqUzLxj3zh1iMc8W9syOPd8gLrihRl//ZXw6iS1IWGF
bLtYhRdFbdg9d6+PiKJRMuR4E+Sz1m1OmF3GDqUu11roj4pbown2MKKGJoYiK4fvukcZGbc6f3Xi
NA5TeXE66XJSnJUcxDT0vDb1SQtzevry5uP7o5h3Vm/t0ao92zRpWCkhF7UlcPLCdb7D9mymuqxl
ygv2dwcgMJAPojyOoSdMHTGsIB6lDWW2JKPEetpgYYEk9j2najezVUxBN4ve61alPaojbrFKEi3V
hT7RnHvgTg3TO/z7StlDa5dzfUl3dFbcYtw0AehU8qk2GAQqkptEVA5qRWbfKL0C9CwxPqdPfHV6
k1WOHSQWL4JXZV0gDcsMmdHVECPTlebThyjZVZ3Iv1E7mBlEuZdEwy8LSAz7y6bFe7h+aIxh6V4P
SNIl8DPLYiLUpTU1kiWMtVfLRdJgKJGzGFYmEfdig4Zglp4E+L50JvyyZEjkOW7SojUNbJpV0UTK
z2OTLJhbt+AzZMxllHKLIag+ew48Jj2q4KS7FQqhny6PlEOI9VESvuGrfhUj0nngNx9W6t93nIMu
AdejM2md+KXgWLMgZb+Qk1a6glNDVm/+ajBFmXajfW85mMobRmpJeykxdribMXcOvpO0jSzSOO+D
FPCdVPCrgoqPnyDrpYhAWLMgNny9Yj8kA9l0gb8r47GKcibvVm7I4/kpdO3Dh3PKmmQ/GzFLe+zV
4e5WMnUMpsBnH7GiTM2+xrCmtnYQgYLWCUkocaYtQRzV8Bw+ovDJ3RbVJ89kG2L0RkXIWRHmpjaI
SDCgCOFkQUT4UoubLqI4NalDIbTxN+U32kMIDRBOtjrVU6y8tcR+W5xxyrhdPTpYrCqRUQUxyc8G
VnpgHxfu57tEvwrseRsKQtN4XJh3qiJDZrHwmEdfLU7dRlEnWSMGKCn3iawl75solDrEKU4e04T4
x7ZuwzX7jwNC1PorUeTg0VKvsbSjFIZsjHhkHc1upOX6sETLIJosTOjshy5vZrJnpAt+9s8VzLBI
tbdxqIZ0DdfQJKY+odtfFrUwHoshq6WMVUBpzto4TR6xmakoDjRX5hiJ+92nVRdufwFEBMLj4Rlw
7I+s2bJGqLttlu4SdlhsQN+pGkbUym16hByVxQpZtKPJ6v/UzX+EthQyc9TZRhlC/H0lqIuoRHUt
O7TVxb1TEOrOy0ZkTs0Ttz5E15tYpk8oR0OfnOH9/Z5YP2gVVXQ0RWW1w0alBS13CVc5qamS1u8f
AdBKIP4dBogozv/3FCgq818igQfsJk1mmOj0d+hIhdXVIQvYnJx6zKMW+5BxwgQdijwRL/mQQ/md
6pzRYKOm9k5s1esrkAjLQLcfTY9mzsfwU1UPdJJT1dcOkNYxqTJwwOkucbjT4mUL1DAJry6nVAEw
DIsuqL/T/E2AD47Alq9ndYtsQKmtYJ3zGhbwrKyfKuui9q7KNowiLt9P2SAfQmy90z06C7hjOHmq
f5kkJwWmBA143ppkj2+l0HnwBT1/QtMkimT2/NEPENCtwCkS+m034Q59yw3AZCnb0yBDcvCL1WiB
J3AFlVYKX+EiehJuHLcbHFm0oqHlqidFKgnhgA8E4XqjAAGbKaWVrVcMC0Pdj4i9NL8bA6EDKvcK
yNUIPFJgWaHRpMU4qhkrK/jQaEDrIW2VVnFGbT8N4vzvGcumFjpFs4spHny3K/52kEXRVX1yPYXG
38w+A2F3346T0rOuaW2Zf/ARTjiR0oqwCKmc6XxmdGFwtqRp9mc014Bg2Xwuupuqluxhd7KsTZuM
IAZMDs5lwo1X6WxFykAvmccvgcg1p4FCELuc5KxHWT2rH6tdU9WZ+4+5lMw8LHsJUpI2pk7LfbUE
//NBMW8jaw83bizYZIOHoT5c8QGZE+MJp9vnSbTcpmqVyI6DBxPji/z4la13XPhFej1U6DMBs4S+
yRSCcGBYMduu0fMtx9yPIScPHKM+57jHtGn+xN11adtABicl3xx7pKDtNQMrTBmmct0WzNMj8VO5
uQtOP4Bt7Rcsm505KN37t3kP4khwuoVvUQlKTETOi0bd38Z/HW7AerGwFNfKV57Rw9IEJXznMS/P
wo5hCoAuVoNakgFY8k24E9awZBHe5PZadecvoAApuGNKua5y7tGpB7Bgk9EFUtzwv3KnNjkltc+X
iyNpIaWQyzyV63AYGL0QTtMd+9fuNkDI1jy5Eu0/tMjm4i3WDxSX8ELNFd3jYSjk7eO3f1cLFI9S
vXdTorZJpJS4obw2GoFyMpUrrU/2l1dNZjyjvqPNveGSw8vtpgk6qjwAEPIbojbyqOXE06wwDhij
m+G3KyO5lhNSpgPQm5wNrB7L7UaOe4ZiF3JejqYvXfQ1pBBn5agIYIrC5HMuB9QqbcQjBEI76wAS
zUN70M2JTLwySF3ohP96Pb3WHteoYDKax/ezxljg1bmI5dr5CplRJ373I9NAhT9QFkU++J1vQU7V
XmNjHJCWbCAv9+Et9QEwfoBieOln87zXWCAbC9B3GSaIEADXKXgGi5/PcEMUyjHSh4rOMWik6SEA
JegCJmxirQ/lTJJiyzpjTRdQEIXgvjtI1NTKASgbjmd9RXJkb6RKbM1H/hF3yPOFqcms4TNUuyul
BjTK0ccFEfrvTwg0M0pnl0y4zG3wyM144L4ygzQWf/t2eL9FuZJM3mXtnmpwvo7Y4TYUT8mMrDt4
EhUXDfdnXrdEHsXFdhns7geg2BRmZzsJNEWsvDzRMIa8OxPUcOjzaVR2QG2aHWtyoNaMljPHpI5z
T8axrlPSKfvWEIGhzC2Jdo7JrSO4asxsmFaCTDUV4N+BaPKmpDnEwW+fiNdc2qoYT24Eh7pLJZAW
kPv36cw1whVJxT162/F9oUQ68ipxo0pbBR39s/A+eZtIL6wqX/4+eIVpvaQDfEgYDAX+4MBW2NUd
ic5bZUbmlfQdindp3qjfE7u8wMvjuCx0U6ZPumdozBqeGjtvMe3UQlvQD4dEurh26OzWA+G5yJzc
aH4UAeyRtre+d0hct8FTM/623Z8tClFf6ikAlO18TE0Jsojcx3o46YiVigKXFVaeU0x+2F1gIqnP
Bntu61nUUU0fcbfSAqfwB0qKZ6bVECj6wF5x44+VZShZM6XFjiB6snnHqN+uH366kk2ImoQs0OuB
AZH5i/adKWXNZrq1cPYJuxUxL6rzOUQ4fN9ggeXdBOtNde6eQ1Aq3V5jr+A1dnfvHJqxrI/OCYED
mRknwfeCDSvdWMAieNIGXOHWk6k2w+7PFIqVqduP8EiFUmwaruZep2grNyxXxqt/83pDIYzInvwf
U8PHGGaYsJSE9IZYK4czk4sMyIznz3MG7vIBiKi1VxwtFLk8XMvJf1UDl6NpPPd3Ev1Zfer1ytn6
4wo3euABWbiDgDRWD1nkD0fFjX2+f4RVfHmQwx3tX4cR7isu7HWjTYwqMqB+zEda7l2b3xRrqdVX
xsnl38nfj0m3ipVPuFzdcP6kfLoP8+WTeMM9aLWT1jt1I5QzBulpGYRwApSWQli1x6hTccOAbIVs
bZxtkEdiBg8C7gu5sm7arB6UhVqx1OUD/OTviGOmtQlQMpI/oK1Zelv+msZ82DnCDgfjkX16mXSA
Uhvod5bSug2Ou+8G5pY5T9VbK+kFfua9jM0Z+kWI+nokyHA8Ym7pu0R8lziTCJQFXQcHTYOlVCYv
hPeSxEffAlfLtSSb+Vp53RBpzSc86WUGfAbNtegQGcgMuSoBsiGUhDgSIlzid3aMlFg+2eoHSgB0
jAbDwkEcqj0/tK2rJjJBiICAHrPnFi3l/XYJuFq0SIMMk+VAZf/wMEQu7qjjhaKsMnh6pVkOicex
hyRhzdVDA8bpWgK5fLvqj1jiIgcF6gkYkxc0Xkv0UHIpCw1IFC8mX0dqU0deXfrmc1GBMC1O6CUZ
QeDBqxjPcbU5DzhWxyf1xEuqpbn6+Vzr+gmrZkJ6MXCNZlop23SSHfMR8hvQHFOnFVDK6Arh9ljw
6TDYOavyKDeBAGtoFMFYrH13jtnx/UqSvI8g1qQYszuoy5wJQKS2GjybNJKd0MMS+ATqHN6jJ+WE
jR4pPDS8JwD7aMVDxRyHH9WOw/Q02kCW7iWrC7hFyHZ8cRR70ynequMUokFoKszgvVQeBbgG0ybY
RnB6dI/1DBSwINRj9PpdEumO1awBVrAgwSBXti7R+IUjxWXs1xHkz5IFMdVS421+nQxKFEQtTQMB
1Joox7Yi5riFQY9RRu/v5sdu6ON6ZisKbDhDDW8pl7BN/Hh9AraZaNCfNyvNF5Sr/JErUiZ43U9O
OUSKnO5BNMBlmnFK5XobpUs2cqM3Do/eZH9g9aZePZqU0gSbrHhtNgdkk+5P9Im7G7gWsX3zLRw7
r2la2ZGHsDw66fw8hOuJefHw92xnQgAuTt9r8PkILpyxL5zocCOzVH+1CFRA6G6iyIbrIwmEBPjM
dIPaogqVluI7BNzdpaC3TgEaUfIbyrBV28qRnbisEj3ymXiYRY+0rjRqzVJ42X4gEXvyTAAjUwkj
EFeQKFj06cCIgekddTbKSjHAoSU+Sbd+KoixSan5v5F8bOknqzFGefPkRlL+RfLpf3ygO0uOQTMV
iJUynwIKT7/WlIAGyX997ZoaxDqzxF/+vZC1dtIRzsL05vx27rKD8PW1W8khns3VUOWIgkMLl1/s
xKGsQh+AnYgGG6sD7o7Hucj8XVeoaNVrH4oIEPAMHwybKuNSjzTxI74wP+yMKpU7cpzNQaso4gpD
y05Gk2SEJPV769fBof9yLR8LV/Sor028GYj7G0RLxcewk4E2ZS9Ty24GvvVyHw2m/iaJ/dkq/TCW
s5LARHQgFUTp3Erlyku+NSFQrm/HkslU7J/u7gOEQKml/951XYCqSdUAN4mDKw1Jnikh6nDTSavv
g53cdkmcjrPipF/rgXWvhl5dCDxxaisz1DR5KP/ybMurfBUITtm/jcKqLhcKyeAt/wNzvVekZ2ZQ
Q08cQwwpRCAbz/8ux8NLRG4KGcFJZv4YavOr5jzhBlv8afZqHvWmDH3AyqmTvcZZsSgvFxb7iPYy
smLnM2JLHmaw2Nr5yIWnDJPInc/P0gV5ygQnHHFV7d+f/qWlJ2NYXqloyR0ZJJ8iOJKUIGEcLBqJ
Aca791G4rvWviaFSQSE8IjSSa+zA0FeO1PkfUMzObNuZuK/3/SPHEF3v09GsnnFtGeHJ+ZzZN89J
bLJhrV1t/Nfj/HeZjtdB8MwT5ublaWSMmJV7nbR3tnv6ccIY9L/57mZ+tnxlrdynzoFEgJnYtSwm
7ndyQTDv5eTi05RYmf4LusPNBGXoQjNkumBlsoT0ydUh+xbEsgq3ISWKBwSrxohhqE5UsObJ8PCP
SkbBUSP/99WSsWoOoOpfWNxPv5/y13MJZjFm7OHDvu6TuxTRSWJwUddXO4GDWeJ5ykVpbUfXIBLp
uy377QII1Wc7a5IUjffQuj62TO3EXhAWLD/qw7sHEnluxLetpZYVng01JPP+YYpnYVMp18qQgps4
Vq2z/00otBbjLpaRoW5j8zWpXBjT7umalcrtlZI/++GQEPUSQ6WlQ5ZCGI2cqeXzyt/pspw0gauO
8B5epJWnhOyjuEnqq5vRnY9tGduG9qyVVrRQ4DqA2AYgzkvoW7iI1EZCxox1ahiDiVGzaj47Pqp+
/+D+MTbDCO19UgX2sOLtTgbyGnZE9y6lhghfhnMp/J4Ai4MwLujOFFAnuUjxWiXBnJhOkkD5IwUB
klHHJyH/0ewrdn9WU+dD3dpoOEviw8Z6O9wtg0EQArVVwdWYwW3H4EeB4YT1BlyMXrzR33jlS9P4
3E48SLk0mYtaJBWkroJ5OqpznXLaRFJ71xjocrfc6CIA9pUJ2cliqVIgLbmK9LsWcFGV4ZtfGzdB
rjfb7ptVZ1KnzpBtUz/lWg8LUP+jAAGJC0/3fvhBAMdPX3QXlOAltiJvY7/oNeL5ieX8e8gv+ILL
vX0CSq+CJZGomkn6Urxv4j1suCo1h4Uzlebl1txeG1qd8IFQhNuWzBjs47RXO4Izmo2GFsSdoKtO
jOrBw1d5J0otyjmNr4psbBYuomM6EG2rHTS0da6kl5RoQnPh5WKTHHKUg9P6DrfTcJ4y1AUNyoc8
Pc0kU8kKc9cY9NRun8O9U4etADO+RG7UW0iv3KFNq8E3QepLuV41V8F6Htfhfmeu+BYbohkiNZ+D
aVmF9Kdo5Rbb2BS8gp7LvaeH5lhTpKXh6SWO7pTig9QvavxMuD1JBuCoA+Zvyxn1ReMPb475/t3x
Y3exbIrNemSX7Uw8m72G8kw7C8L9X1nsCkVR2dSi9ZeOV56KsMCxhPyN7CME6EeJ0/tn0s6pAbfH
ylVzRL3UwYTf53bcL9JktvHN00CCipWTqilIRj8123XzG7YfFaPRGNhXwhv/yg6N1UiELBnSuwAC
tZYoKduTEYFmvrs4ulGjvHXTqZM3VjOTrUdJkHxDCLwb1gh5/sOKTwTWZ6+PyobltScDvRnHPYz4
gHy49W9n1oBWzDRVCxemBVM4HXXImXILtfiRH4+g/rfnArNLGmM1rTwUiAxKuB3HeW+oO6WrtZxP
xYunM3fnBQBDcvBn5Q9SpJsxss1yPypmp9TuNPRP+w2SsBo2/irrZt7idQrDBjhUZN08UGnvjrSh
TWuYz+WutXUVfcTNwnCPl2xU4qZfYXz6tJUuTQy4GR/EmXbW/q5huum9XdgLAfCDoQ1igS6pE2GO
DmRugOMShMkcRCY0HCSDlt8Im2KuyvXGPSSMVo2WR7rB5tY9rEYrJ2y2B7EVKk9H4oDSWpqH3the
OyRWhaLCr6YcncGZLFQgKFhzPnn1NIvXiuQWTxUCnJ9d174NPkC4l2WCdEOEn4zdpGW8v9fMsXo6
NFzRI7BSViv8Qued5YOpxZ8K0OQIBSEHcDakL6uWDXL6nAAhBfoBmTO1m+Vx5FsBzz2xNbh+o2aw
rvA2m5dy5tfMs+c3bGKz9MaWtlOXjCs6+UNfnxfHSbML9E2AqQfz5Jt4Z8wg18u3enkVlKdTSHOc
nBtwQLgNxQeYKNVdiHQkKHmUA+TEIUo1zs+QP39blTk+T1tRZCZUlACnJjAFQkDrSESJqvV++QST
4JdQvvdXD17sbmC3a+SIBunHTOy8SyG+6Qq5OHQECF4k2LSZy71SkXnks2ve4GJjJKhHPfKX63al
oFfTK+oUsEzNDIFNsLK1FV2gqHbpfHfmnVxg2LflLRyKkOFq1Q8eW6yPcW47NZvUDo/pWrCEkUel
NGevaDksRxilkLxjig0lM7tdpsnJISWXrQqUbYTD1ExqBcNaR76+AT5edO3YREIQjYVOSxLaYVAs
05SEmtnIBf2URjKJpRpNzcNGd93IVM5m6VE7Sy/fqSBEDstMWMJc58CacTHzQedsYCRreG2b4IPV
7jFk8Rz8o3b0u1tFJ9Hpn7Lz1NzfpeKeQzreVpwTQ4BOa/ykMX4eJmAxs/foeuB0rBWBnFxI3n0r
ye/LEL7rhJ8KxhqLEih2r6hoGvrUZv4Ls4at7hk1IoTQSEiwpoHTHfsewTgG2MvaVeD+lKG5dHk+
825q4PjbHvwEeUi7h3l9hYsS7/Sbgwy7Vy6HY7pt2uilxb+n6CE+hpenaG9PZzixgeJfnGpsK1DV
azooCyj33Yx1zWGduD/oEmJ4/xOq2x+e+yfMKivzAeAvWcH4G3qYzDv3q0NzRCW1CzbCQOwTa1JC
H2DgwI6HUIYpEbcol/Cct8RNk4olzF5SK+bhkWASPyqB5pj/PRRH6aUj325Kw1Zp3RS/lZVUpI+z
FbS+hI97xmMXdkikEEeILlu/t5N/femO5eVkwALelWbwcyEpTZplJx45vj8KymIikbBVEytlkTGp
YSvGAlPIozZfqRaFot1ffRMY3YOli11ziahyRoQtLWRHbscUKUluE6n2Es8s1oXzk288OFt3pLHB
dlnWoeQJjAxZ+vh+4fbBkAkbOGFdyqLa/GTTizXDGPkNGMHRGXKr4pz5A86hPHfu7yh276jUK6Uc
aX72h981dVd5b7HN1h6orEVYAUW2cRA4QelOc/xqdYYFUzAdOkYv+eg6nGAIK5zSxLFJ7PQESto6
1uuszrxCiMmuSBiTOdRltepIpxzIIFRufvZTmBsklry35laeDg2AfaUgfNJKxPrY5EKkPeH3vAqU
hEywZVWjMKXjxgogFwKz+5JOQHgVLnlhoNCxkWALfKGSJUw8wsdGI8cad8fkfwm5Z2DqnIdn4SQF
BkSxiL4jn7XrgNCjPVH8YryokMtt1N4tpO9oBtpJaHj8fnQ3ybcHzwVGjk9fF6QfuYh6uv6oN+Qr
m8BTOkJdR0CkgApMbA0hdfXmP/RNzUcKDiMAUlNnezMPm7PL8KqV09kOBzkzo8LAjLhc2XcKgIa8
wAAGq8ngw5Lbv0CO04kPHTYgkgFf7xdQIkS0zOJTtHbBpncUQ1uH38GPxZGNzSnrpZLO/m86S4/x
EzzD+zTBoDP0B9oiYVB80JQhYuqosW8wBF7By4uxqB6qlDSTyO4DjK9MpmXsdflNE9MZHk0geUHY
Qa+AWfinPY1EGiKMnlmNPKLdOFXuY2cQnf8RQpG4x62bxtONSMZAlCK/BS8ojC1KWVHsn4DKr9hk
5M+EDqdNK8lKpZ3oeNqlweVwmubhsy5mv+76hpiosYkkPBWCB1zdQ4RzBTfzWn84t2+RM6Dq1sTQ
P+ogsRTZguKEjj1ML66c4uhwsmhFg7LNdZ++aVUPPQhP+LaRt/pPKELAMd3xrKIvoitdwQ9Cfgah
draGixGfVBvev+W9lA5ZNCeRNlszWv28urb7vZ0aBXI2VTQjCzGQevJJTphhtpBZnxZIHhkCKK/z
jwqQR6qz+n+XY0yDgATiLONrfXeE3tN+l5BIj8tm3Mv+MsfU7ZljC3YAZYezWuS/KY0dmji2b3PF
2Z5b88DbbRv3cGCO5vIu7HjjOqv97QICGFVntgaLFa+PilgmXG4OgSSWK2u8R1ebqPewD0J+s3Hv
Ph8XLI6OyjD0IQxdkeR+DtT6hJfsxHurAXc332dD8nI7VXneUlVWpLZkA+riDkFLsrz/C/Ug1DVC
zyJmc6a84YsS7JINGCYWZkA90luQTAwvYnXuBQmI9OO9RAglhCfyXfgl9f+c8QQ98CeUq1Bzxa2E
ZhosWfkAIEpNKERMTlxi+/Vxt3Q/I5e38MeR1RVjJUjz+b9RVBUT0UCnEeoMtqM9lMRWlJdWzpaj
J7LxHXkX4+Dht7Fj9nYHb1FOhVipVbmaT2upqQWPgxKPHPZ9hbjT+ioIwCQEDl9hhU6PMtuzAdLW
2uspk6+r3P5fWm2RimSBiCspGHbjR8E6gH59TZ/TwdeswmmmHZ8LuZPKg4aiIt+649iEVwS5axew
7RVer+ARIbpK+20R6Iac/wj5zTetFe06F9c4kYneC1N/P5sJvdqTLfexZlL56r/rSZTmUEdivrzq
MGwXBijCSUbSq3/nfnQX2IKf/vOV/4vTVJHTO90J4MdZQCxrzyrAUzxQISl2jsj3oh7R42o5oBSf
fwlHxEbITWCAKoYpcFILrRxJfrtor+YJTwhDVXiF9kZtktYrax3Sfe2r65uoVh79nfL3O0QjGIYP
0DrkXYS2TOkjXt1TGVTBlWE7lJUq0ww6mTqW9MU/2injua6Jk+ZszCxHCbAA9DvDWqs+s3VC5r79
BAphQoE1doAZKpOCr1VOoaIPAQHstkha1yDCHbyVsAzEUci/eX4GwBzsKr3WFUqo5oWSoD8Bfjq1
LM9GfFCrAuwH+6aDvpUwRZSjRveBBFcS7vIy/H6YXa61j7CpoiWxrHNIHbhEJqYiSSOUWdEu+yZE
uT7cqov55SFykFVWa98xrImIMbRRqWZqdGnV2hK8VZuB3UXLlFKYzZPA3CAlUhHOwHcZYb01FkK7
SW99MSyKiH6HottPRrmRFDz+UkEA1r2K3xz/2URAtMSwmTiepAVAUtmc3Syv1C4Yhbq9j5EY4cfX
kvVY+rkEnU4tTGXZbJR89dfAWyZew5u21GP/JvmUqfm1+1mrIUZXEyLXRoji8fHnFFhIeJ/YX3qK
8EIAnjQ5sryTZgvpeKcgkbaDk9EVhDxDHn5glUl0epda/VA5ktkGepBUFDSZYE2QBsgNxtc781nI
xwp0jj7AjlrkRZPMRf9SgE0hMSJ5AxLkr1Khl9ZXXTb6edGNYKNiY2vGxsTXuDOGsOfFSSeMkDTh
AWi6xY7nrWs/vpE3Ep7vB0N6/eWLb1wqq2qaEFSxy7OTEuNgcCc8UHvxl4LBtE1IfjtuAG+Lq2Da
U5CqxzoX0IUYEKe+rZKxTFUiC1EAKSTdAH9/3USXrDFU4M/MRtpJcgzs9KojQHSK9xjAc7X0CKoB
nEmJvN5RMN+DEGupsNFe2KSDAUzObkZV+ICjUFtacWoGcGu1HjnQtCxui5PNLSILb48IEE7SFq+A
YHSMouP57esmVXy+YyXzpgLS60f0XAT0nqk1GcOOjb4VkT1sFaL9tzYcC77+hyvx8+U298v2GOCq
lGbGzLu9IRCs5auvXlbvdb+1P2WZzy/SGaS/Kau6UqXbxuW3sQ76JpNvKy9eGWyGIsMoBouO3f9k
JnbNCSuum4khJZoWVmSQmcTsbhVLV1KINfJLGhHGnJs+dWcj62ReGdpdYoe72Se9ERFVX47iwC2U
hF4b92k2R7duxpL9cWYSvX1cCmmSnnfTa7TjLAJuO10lKsWRb3nxCYlb362LXYG1e6P9Nab7XDUL
40xMLMGrZoRKscZSbuUNNEP4PBTCQUKFnCiyCA8tsQz95oBcDXj7DwhtTY5Opiu9NiQ6+ZQB6zE6
M0NvAt+RL3a857kWGjxp56e20OXYGFeAHFxOG8KN0jq33duM5LSpZvI5wagObGHKQ3HKMxkwyfIP
NwobPwWEsNGzQWQbCWP7vGcqkVdlr1vV7VZ5TRfeH+maK1Ga3+hKdyJ0eIB1yasKqnERZ1iT7Zz1
uGWbP/yn+3tJavtlaDKlF+ARRJrlUY45LWvPv0FNDt0dwluCW+6b7bkFupgQOmBAtc3nM3SwK0TN
zym6S6cyODF5mHit+ecimQN8Boe0lq55w92epeaqOxKDcfnzxFZQTfAuo8KqyEoXgj8tO6gZJ4Nf
UFyCcYZp7GAdWezb7fd3YhrI6U45ZHSI8Fq4lmkNyQVTWsaqnxufETo83wqXnRNvoLMrUe8y43Yo
R1XIrfyev7QaKuzmjKnH+X8a2rrIzaehfOglsq1+WWoVuLUIuYTXTVyxlGsQpGVtVxdzF8ivMcaT
o8EqcQSq33Vvil2LcnQFcibIEflF836lqmZ0OXfCbRtajLiMfvShxQqoxUe0n2eABdSrK5eOB8+I
1ffzKcwqTmlQYHLRvSYadq3YTaOOeqV1mXMdleebeBQDXaRpqtr59I69saB6/aAgTr++DyS57JRN
/g40ZKQamDrZdc6KrxT0DZBJR2L14meIt51JVd6r7jtFO6LgwplXRK89SH3/SFoTw86gacNex89I
mM3MowazNPNXXoCziJKTgbjhla+RXp9JPQQqGdhpppc0OIAABtyVT3PtL3MaxkenhLxoaP41BiLi
T2icb3M+UNUocVmKt5bG+fy9eS//1UnAd37FkJflQUyANB7G4MbYYF1+FjqgliMFaCTU8s24/xNU
CSFNoLgdkAkDXk6BEqKD/5oCjKnhnqSXzvJUPVbpr3sahr9tCChDCpMYaKmO9us/or9dfbt3pFAQ
6d2qqvdlPLWN9YDzEZq6pgaBdw56pbtaiB1EG52prytXj4KdVMopnVTMJo+9XbQaFtVqzoP7/lMu
7f2PCn8764C8WXCv9RaQ2pBADnLRVqTxJE6Ya3GPImoIXu76KOPP6CouHPBTlHOkltx645zxQbV9
G1naU75zcLJ1y99xH/vMvch0DZTbK9DjFOFZ0+wn7ol7RrhVjSSID5MibEuu9zpCaa0bwyiuyg3A
1D8QTXQpOLxiKrmkEuGc4fBtGrEdQeqV9F8JkM0ix18Y/hA+wLWJIwdJYd4GTl2M6SDNjo2mx7Ya
V87Q0SEzzaYYDuCdM0TX6Zqsgm6CO1Gn8R68VMMnYUculrDDLmlkgczyUM3ZIdRfp2dYAUW6xyjC
HYEvAhprGKOugMfM6pfw50n1737K06UxtDpqj+sx/+f0cscdoh4CjGcO2ll8kAze4eo9RnUAnEgn
8a0PkY8vLthNRgRcSbdbcXMHiG1wDEIMX5Ynb82WrWGM5bgEbHw/VHxIU+f+C6s3ekylBxxp83ov
NLrHkWH7l80sNfyH/nclgodi08Kgsgac4ST7q7od+02FaZ5GoxgPNKzlSEKPleXC7gxHPb0h8uj7
JfaTNOrsxTTGZ805PzXQ3C/AiRiBSx5pHj5V04eBH6N7oJhYsx6Tlk5sM04SiYWaufE1cKhCJ8Da
mlIwBhQAiCQ5pHBwYRxGd9wWoF81ZHLhIgCKh85DHdNAIuPmaZBtpnlIS15bufgZya7hexG0ivj9
tmhLyuoOymDYp3UUouKcyE6n/jj2CmPpro5uF5pTV3gQMd/THikdYqaF3veFAQtHSuaD+8vIXFqe
d5XwYYWGR7cLckLehKsq39N0kxENDoOQ25uxcRE+t02UcTLgifKCa7UwX1UeVmyHccmx/RNCzcy2
M+8p+SkOJrP2G796+8C9Mpt9zdeCWU8fq17UVkORg3kniwPWsTThnHH+D+WauddQ42Cb5YZTrtw+
I6cJFK95ltXsg1BDQ9UncVR/lxbk7Q8FF1BFwy4i91tDzYlxiGk/AmZ806b/uTmu1OsiOrSV5w3L
uYAE5x+qc/qeWfdbrLA6XB/GO7YImYtNG3fdHejZzxY++KLStA5GT+VMc0czZGaBBzQszFvFeN2I
oyVUkEUjJ05Yw7IdJRAqfMx4jHR1+jiJ8wNrAN0H0Y+HeoP1NNarEFUf8RPM7n7tToV2eFc6Ly05
B24JxwwFI42ViE1prrSwD0eCsz2F1tfuq7CrhnW8OBdT1cYwLa+qeC7SyF7MBAXHGjDMD0S4zCIl
haxK+XEw2SMazVigujcSQ9NnCzPlJoiYO0GzbUhk1w8wkrLxJo2S0SBRd5j8rAhI8P3FBZxsHoHS
A753f/Y2QD+/JbwwGvQAF1N/X2rMv4CV3+MpwBFcYzHSqkTkyoFvZ+/8XPKSO/eI76fofqG+1/7E
FR42IhMdLBHjSnYM8NSHWHbQYxl7P0PKY1MwyV2cjRyXqAe/Og3ob98P5YFA49O/+IZWNuvqbIOh
WHztKWo8WfBAnBZbCS9KfaScreM4udNwD0cqst3O+LnXp1Z7vpf5DXgNYqZHghfvVgebe0LhDbCD
jmt+QoOvXJ7cVZSD9kuiAWciUg3mrTsfb6xZzHzT/kN2ZR+3F0YN66tXpb1NjF8mm0N+oWn4z9d8
YqRMZAM/MekblYNLaigcqzgtEPioSSv11lT/Su3z3wZ9VGn3R4uLnwDsrVdsq/RA8BmqMSguwmbN
ObcjHmv0pJqQypmbFCOsD43rOvhPrKPKgFYInCrFiYVsZuEjTPnIrpnvXKXIS9X/KI6Sohbgiyj0
G8h0mFTVGKYN34BbqUF4f+gXq4c6N/JZTyfNTGZeWfDC/CfOETVyK0G7rB7bCOikCi/jhqaxGJ5o
ru4GI9bl8Tj3k85HusUojNdA9erUGt0LlsqI2V650h1DnPX3zv4vpePwVPPQMpnVjbuMnvcFA7TH
0RsUPoauKt/yK/1MHKFhXuDZRrl2r60GjFt7ndUBrNV21l9H+/O+lExjhFsNFvB8yxdf0mWfYOps
3dpmjTIZjs9BPo+9PZDU6cXk8fhnH3yDvdOHBu1fO+ceJLY/xCAQjVSanYXIowDGGvA31q5aygE3
hZoKP4umbiXpVRVzfphRh0sme68KLgkSjW2BovMSkO5cf8fc9hbfXYZUINANg3s9yfBGYF6LTC6a
cp4T6oO7vW33aw4WElnAGsLd4wLwqtHttdO1E2qOwdloKtKPgEm6GAkbhvzY+qzqbA74ElFIj0Vw
MlRXRvFv9QcNlfnd5FlEq1xOz1hW/JxoLQMyuIIFVDYxr7eMk6D8YFAydmvd4Z9WTOCedMQqpolM
HkYxBst0gwlP/1K1dHiSs9KRFilwBI+ZJG2wE62Q1eIqra7hvveMOFVDji+QKAfs1o2wmp6bwQFT
4KnvnKxYw98GFckufULUXO8DAwaVL794BUaYGiE2Qh4ycs1xFGImLxF7KLqSEHcaHbwqMPu5+Loi
rTDfj+KImINipe9feYdZcR1VsvRvGmneWTypTMHMnJ8TfOtRXXhktN8ItjAQ7/uNEHoWoyYxWQ9y
g+/0wjSWnJDJ6N1aMENy82wrxVqEDZsJACzvrnuV4kfIVgaPSu3tEQQXZzSKFS88/K0Dr9hjmPvE
tp6l08ueWQ4ab+jgUBouNy8BpKn7rEbLmK7I6wLdcxssJoqrY7bvO3QSmajwHnqV5z8Fy8QVCy32
YalSHjv1eaARonlRZJSBNSTpcnd8vrA/MBTYgYsREENJF2R9fJxkez33pQDgC4BDKiK7l62ylnCi
h7c1OhG77A0Dmk2gzId/0jBu6gbREPPKzSWKjBbOwu7SvXdOEyBP2ckHoMuP174+QUQJkGWTmfMg
4NatMjoUFwLl62MhyCayug/QFGZKPVH2s+aPGywO0iUa/bO+Rf30mADLMV5fEtWGvp8Ix3DDrFiB
OvBcNMRh8oMLYbf92vJCnkQdH7N5ClEktJ5fqictdyhpPsNoze5r/uCCyJrE7iQ2DFtvTxD3cvvt
/DV2sipGO4/VmyzzTivKPXJMgYocYam0hNzeAAw6OQ2XhyClGh4NOm7B/GbFKKv0o8YFoVo9LgQP
jKHPpAXNQYjfJvYthANDfU+cjUlgDdFifYcd1S2Z5FahogLFvyt1SQ1aWmGHw5vljRMmEKMXMmOi
7Bn+h+41t7/zNsqhU8o6R7+mn5bWKqwxoO7dKVMrGaj6/ps1QYU9Ua0p/JjrRTErRwdR0G/ngWM1
O3h/1MgH/UrXxN54F3sUwaVOHemMZfc04FEtxu084KTFcre7quWsoEZuphjK+Iqxj8CpYyLDygSN
u0qV2Zxqv3xnYy2dJr8dc4NR7WbDuZPRztCr3ww1tthl6ybrP92tkUjxwzEhN4fX37puh8PsstIX
P9vi7siGxEIbt3g3n32RXBoIh2fGyzj6m6/pk257DBCEXVd5O1PKoIGnHSbKi9a7urMYhl5yYSYo
Eugnt6nMaeRqanRpLsTjV9AVnZZng2E21EVJQPHcUZg+Q2hYWgxt1h6DUENr70w++7TkTehU+UTE
jgaS4jRabyyAtoa+qLL2rl1JFFgh51OQ94Ix0HgATeqBUEXRho3t9t493M0oo7x2Wcvbl6FnujOg
M1ypOUOujP7t3JlkvO9/wDEdzx7zTKMnSSs5RsNCxDqmn846dp4GS4UXUCvQjNTLl1pF4JugAIh0
WspKMWoMGP1vpHkxTD/MWZZ4fPHZ14A+M53VR10d8/WdcGN90fZP3+WltJdp73iBdApf6V12mE5a
FeKUNj9apDoVOmgVsfB6zNttf1psOfRD+r+RBKyHiYxd9XfxxCJEC2Akg5teyMPWS8MeCBVnnD22
RuBQp8EFri56sKBAqAC3EQ2djjsqMY6ULiydJuv7L+5DVbWRD8SjBDyRqoIbWtGHrQ1rL0Ib0rgU
QJ5mU5dzdI3UnbCWZwDqZJXhS3rbbJYxTNMnhkpWXVj40NNVbPyL7t+qCwN78pppxYqiS7ig1ROD
T+sMM7cZFSqUyRBZWTHB46jFNVRm5E2qLLuqk+XpwybG/nJ+cS1Pt5XN+BElbCXS4Q7YNGAwTM6P
DF0vBo4Bjnc96kh3DN8UCS8gtDNDHf4OqfQmo24Jj8AUFwjt9WHHs+VmBp/VPe0p4CB6mVHkXnJk
E19TGGTy0yg7aFJ36eoNUDpioEdxV5C3NxpfhAcJYDSCy+9UbVmT6j24eaML4BppPxu1rm0oW5Rl
dW9mOWS5pLn2MeJU7aCGXjCbMlY78XXJ/HSf9JPbitOPXOuNv5GRHG0O6ddZl1T+ORVX2nKoT3gX
pH3/zwc5g7aacsoGx+RiBvXuNJyl3boQTDaeW2Iyz9IyGduog6VhjOF/ytaJMRAliwh2XIeJTS03
qJwZbDpx/OqaM4p/cosEzJTn/oiHB5T4TEbbvKhP40xFAjHrS4aZ3mdKXLrTDUXrbehyO46SmmdZ
wypysl6gJG9tctiiD52/goTPembNHREm1Shukohym4lGGRLBfcO3Tii+WRMEIsvpZ3D9GyrCXlws
ddOcG4jquUEo1bur4tkIQyS3DJFl6OjHqPb1ah8WW6vTdpbUkPfItOOY+xAMKge896Q7TQAOaGsM
US/JA7jt+iM15CvSWED4x7sD7fphNPd8Fji7Bc+i8mwOJIGYO8RACMjUM/RV9DKSmfLF0HyY0Qb6
1/mmoQX459IorSVp8T/GGQrxIJ0wWcUZw/vVuxuXLdG/5vFaLuu93wZbjrs98uen+VR0zckLc9OJ
bOxRlpAFf5zZzmS3Vs79wxpsR8sUU+ga810OPaXxmtr9Vz91eMUy0P4SK9EbTBHibSYCuU/YeP8Q
tE3i1HOpPMRn1WwBTpRfYcHxRXHCJZq0Q9BaizEZYsJ1RNphRkz+0a66UiL22s9dMQCyDGvvHeIL
ak3e3UIwroupBIiZ+Hpt3CJh1f6s2Cs/kWREIQiEfFIzhc1K6EVRPIFZNO2YrQeV/5DgS1fDVCj9
x4HbfJ0iP0byxsHdeuVcL2F7Qio6up9CWMnZnlptqWpFblHnx5OqbHg+dZ5LrI2sdCVkdE5RgkkN
6AJNJK3exFT0E0HMdZAt9riFEOH3RgAEbIz1GkQpF4VNN6xilKarMCtcBRMXrHmqlnuoW7iZoqhy
SEowGxi4BYdwZhKyLRY8WPaPTkYHRnhRlkfnuAizfIXkGy+dKRfyQBU4yaFl38jlIVQEg9++juER
ZzZZjPhuJPtiu6zcMV0DOXGPtoIDtX8P9FNuXwPUnZE6mBwUuZNa57GN7jFvaIem/qdcj9DfaJWF
gKl8z5EsOmpMkeygsRBqt/eARvPNVZ4G8MnWk2E1juq9Jn15U0X1cORwJSha2UQoTDc7/MNfukyn
NIqFJT7kDajbiHaKBfjLkvG4C7IVOd6LSmt8OkSqnFsd/Bu5l25JCPD9QK+O2rMNO63IUp1sYmZk
3ekW7IZYRyVxX/yrrPCqJ0SbVNFZXyV7xv+fSwoXYwRuw49/58WGU4E3BmQUyzVqZYTXVVDvG5xR
eHap/m+cEDBUlSXQI8e+Nbtlq6M0cCtb5kOUwrOw5PvSxSXptAxV9mWSRJBTrJ4Ifsxpq7nlQLXP
bWaldcNIIS2GMtYpd4+rOyb0WQ9IN21ZzYC+3zpE4t2AiRzAjW/AyANfb9nvaiU5bTuJTOE0A3Da
Y4mAvQGTrqCjebFGsTsWEO5VKpWvlF5g8L8benWz5aQ8A7MHyTNC0K6LRBkWhI8BITW/VES2zZ/e
ayhZCrjSMIeo2Fgs6Yeo8LZFWYh614WVK5dXqtbMhhlTl9toXy42KIZtBWzauQVi76vizsMDMbhi
3/HqA8uwTModsF0HRL4hjP4jJ9vXvghXZ72kvMqYWJGmRMUVAlwazBljhBcC5jhtU1Gchr0KKzcM
ALivAOs2t8FScmhlwZP8W6NbUt4n5OnjEQsfKmZUK7UbIdUDob0uNbDuwiyxLBQm3tqSIik+Ly8q
HUYMWA8wEPGtIvsyrisuKhXW5XGUwtnaG+lIxFa0Toc6pkuQBl+ase0/aLvl7hNwMtwnBC/tKcPo
enoC5LtkpoKZ9mXhW0fmOsMaQYsKzyLjWiZPo4JgfDbJ5WlBCJuJ6ElcOHU+Kl4USPpnqLWu1rJg
pQudW/RmKza4S9nr/Mx03N+3LKSFi7OCsywlEBhevuBAfCIFneQHJgXxVUU+CF6kBXHYJgH0kf1q
ZmQhvU0zqf+7TxgRgkEhzPCcigwVM8H7bzO3Ks7BVLOXpLlszeN7yfpnqmpVPZhZHgGP3oZI5HJ5
pz5onc603cdgGfF+rBThG4ZVoEWDvtIXH6YlP0DtFKJTovRJcW9sYC2hNC74l/cmBZ2wNbhHM9ST
IJSsKevzNJBvvyOxxIoQlkXWsIfW4+6o2j8JyEsNsgHxoK8KDd83zPeCG2BY12MBeh2o7S7QKIwB
pWHsTljF+yZV9X+i/5kBA2+0A50qYBMLcurN2YDfuZwvTiSt+KZ7QJ7Zx4ibkpkKmtsYHDaZb0tV
UIfC0xKnSYV+w1009kARxc2yQuhHk7k2caX7cI7A/SDHm0nJ/Nc4SC86WPkijBmdzYxRoNBY77x4
eiYgExbtMGbk6jeeWGNza596lU5fpy0D4/MFY7tt4T1Az2Y0lsXrnrdZPiVFCtUD6Esm9zGic5j/
pszsJ0clRXJS+HfUEOmBDfhg5hqVcitVM05okxf0+WV6U2MZP2/Vff78iwBMxAVOIMUnmI7+y0Kg
tkx3AYnJcKSZBjOwMVK1Mbs9iM+9hEumxHobhTy3EKjIwLka8CwUKrUEhRmurrXKPlP8f78vLrae
Rj4N3FZcmZhd+sKysHYLHehr15+FgF4eRhBZDZAtQgxcmpHcMbm5/MzLlc/Y93LDyOmztT0eAZc9
eEMmSjhn/WgyMuU5B75zaY9U5VuAVuwkgDD3Yh8w5+t11jkn/QljXaO12EwG8gdtELebqcIe3m+D
2CA0G5S+CayKhPCFZyaYEhxlSx8DxuxSYPwuXEqoids9aOQAUgyED7Xia9jDL+8LCnHHSfGX+AiD
/6jDEyNwBZyzVkFXaGAt/mTiBmrsnufEajsMkr0LSw1Pn3u/vlrvd5rwRDWAL59obRlLy1KqWC85
wwOeeehDZ8QKF7T292EasS13NK6obl7ev+OSdRbdC9JMAaqtmlCLOCfFrd1U2fCmXDebbe7kVBud
D/va7TCcgtKr5XYSxmU73qA7r1sRpDPerpchWExK8c/pCqcFaYAZESYKnWv2s2EqvdzLVXH25G5K
IRHdVfcio3BlF6E15rakxaIxheZWtx5G2RG4Meb0oIzJUA8aTPLpfsUaAhbsxICkXhBFInXru0Qk
173L6xuseHdXYhl5doIuYbipY50qVklb3rzrqy7egLfW5qgRNPU0iJLxv/qgPidmzU8fNjDAgpAN
N4j1Yi8JDunavpTPbGPxI20Rl/mYddQOTsGqQF5VooONj7ygI6utzOqkEsvNdUlWcCT0pNoGotvU
fCitovGZdUh/mriEIiPWVs6nKERFU/nte1WcQ+7SBQqZCXO8c1LI61y2x0pmFPTbf276yOefYehy
367vifFuuSFeHER9J7ZrQILiR5UATA8UAxIyezOcE/5grIwQLZju6FDuaVyV6GimAjuo4fhYI71p
iBQvPTrgqzCLSYLRqAFn7OLCOmxoAR2JQAOyrz3z5PCePN4ERDbyqanqEHOcc7CjGsQkXl+Lzp3+
7F25q1hFnFV7G+NIcOdyhKPpGtMcF5pJRBjdUnVdqfsYJ1XH+tdja4MNZoxCQMmMO36MS9Wvt8V6
wiwlPC3PGDzEFo0fLegrVhQKpSxyateIdUqviRsBO/f243gA7klVgfcX++9rBVLO3qv/ZDse4Y/y
PaRJicPNyyQOGfiSjmFUMsKv7mcZ7oXoPbMA07Gz7CvcpEkCjink7l02YZTU/gA2o38uYoAgu1lb
hdXTKTJJYEADhZ+5jG6epi0HBkMTAjnIEOx9i6G1k0e1p6lfJZJNv1M8XOXajMUtr9k7lDHGNw8c
hhRIIs7/H1h9f8HS2EhZ4ANj/w7/Qzi3P4GypHU6aJ43XZL+Fi0gIfPftn//05Yo8WFbMXWpB7kd
X5RotowfHkosv4Zn4zaSV9X6TDbd3obE6sQbAesedHR2AGJC+wL92SXJyBdAXGDBnVrs1+rp9Sjz
DBx7So7TfffHiZpSzUW3L4lhIuzDtWu60BDYM5AVk8Qpc/972L20eekO5FZsD+diZx8UM+TaBCfk
gEpYoqMbHv6W3Wc5mLYl0mlrQxi/ezPXxLLS5XI/fByz76j7IBjGpaijK1zPnv959rVhvj6vHpTK
U5Fs+cpnaeBlXzkk1eC5aj23TQAEszpBBmGxgrXLgmsIwsmrwfatvXMp72a5KTD09y4nO6i5na8N
cPzLAfGJHlkZCfwFF0xEIfxEIb1LlRoMHY2v2g5PfCcZZu9gV//WBJcuHCYW1HtiTIXEoehyVH7N
mVln6ARkKkDeJSUAQ5L1bS0JidEC40f298xiLbg2DI8jfOAhA/uoswM4XDy0DPOdjVQoLeAZ7KZO
ZTutx5mD9jY/roFuHVVVJLk9Tb3Zh1qMjCyrNRHBp6R6Bje+Smf1YAV2yhANzrxNkQhGgnoyNRof
6dLgUG9Lsz2UAk2xH6SP7PKu7oihq+AqxoU6obDosd3kvd7yUCCeqEZEvAGeX5AMXNSHyn0+0Z7S
ONZe9XWI+SbH+PmyxbDIaNxqsk+4nCsB9fr6PtL1xP7ejspucmJ3NrXTX95hnjE+GfT2nxtkJJUR
QPI6bNLmOeNqnLLHX7UTYhmrHxESeMZ89xMdNkpc5oK4/wNxcnKiYMBs4OyPvE9IMsoWqed5LW9T
uOnHZG8K42yMkRtf33I4S/gZv7rEqakjnG9yKJbdIAhZxf3kBK+yhqi4Dlm4Yq3/5QCBqTznQFjc
HJx2FWsyo4dYoLFWkQtlWk9ku3uR05tVnG1efyzm1Xw63AHnAb9qmmTL6xsPthaa1b6s5fi/MVdc
2F456tvIsUAir/RaYdmnPySyRnq5iDotYHjfL6npgVEQAeKL7W2pkff0oED0STSJplkDKhEQu4t4
V7oPPlGUkmUqdc7gDBuP30azC8yHw4bqQqz1dCJFfjQPu4wDwUWDk4eQ1MNZ3zkas/u/mvhlgH4G
Rqw7g4PjUQMOZcC2OITspurmekRBzF79tMMkFmvg40zXKYBFIl5Uzh7OjywqdGEJnzS0pm+HF9n+
i9lu80ftKrdbPLsc0FzDOjjuPWgPJYzOEVE6KB7rSmu4HLMK3fugy8pXZxQVbGyP9aixiBLf45iT
vIVWyOfXKw+5b0t16rJnNzbF/z0X+VlhWTQ3fB2ilcuB4Uglcozk8HWGA+Ze8oHvZ95qZWXX/siQ
atwAkp8YM1hHWBoJmRlO0ZlGhmzrNY5DORb6nqUrpxINM4IMEQkzU+4fU5X0yGPAzC1de2Szi/n5
F3FLeY5wjiQr7mZFusFvTnsAiZj3i1O/pNHIo62qgurkru6DNGxMeEXcfDMx611NJBgtPF2gD+fX
mKHnjHHKKZZrpawR0I0iLxSvMrLE2wCxZsLmhTfj+2mu7v+sOgtc5rYYqJZ45UQB99EgnUOdVjMh
0kj/2wy/W8aMTRUOMtV8gs5g2LaXxFji7hiQiWmJc6OZ0PDdLUnlxmubLIG2yx0ZvPdXQLa60tTx
1dShfc7A7RrKPRwU5keJ8YMNCcdBuW/SsGCd/dvCFp0eEcGIgrdFwbaDZCok8JEHWPgtVEJWXiAj
AhMqe2rdyjbxHktvaMu4QpLCDsQxqYr0L+cBif8OMUcEfjlolS6iA+98+B8SLg6oFteTgiPdpM/o
ZxJxq3CVk6dHlKnsyQXswuGc+Ltc6YwriTc1DYkogwG1Alc8lXSyeqnnJzr0xxj6NvyMYf9Fe4y7
aXNQQZ36L5WXzUqMfagj8STUlqRAO5LYDZvLQ4Jjhns2Mqpc7rF1vpA1vL8b6NWeM6yko36plkhQ
/wgfNfw2FnPLbpMcZQH4ARluEOw5vRcvOPOpld+eXrVtq/bGsyFex1T6sswpi98dnULuO6+A9lla
0Zho7AYAdKZJyGMp1My0TE+v0fooYCxM+B05MfYGRWyd8HUzAE6C41t7TPM+oWRBYxkI/+SF5u+G
v1vCCTUwwWqDgZi9tdNikA+/z2/LgIBPLI0tpaSLV9pFL66d/6MMnm5WB2yGgGNh6BJ+Lie06OmH
Y52D7KDerSnrRWlsl+9Aiy18pFt9DHvwDVo2XeE0rhuwAqWN/ZNEKk6ZVP9KIf+cQU7jbk2jScbX
QbyPlRCWJAaQcUK2eofCYf0csvvBB6DwJSj2LlOL7adgIhPEGkXNBAi9aPViPr4yjtVmm6xu1LZ3
j8dsCr2IemetCsDxwZ5DBKMJFJ91aqvIrPyeWQzu0i0crIe0HwiQEfnHamGe8kxyLqm5mlRv3HYQ
UyRO57FAFIn7CWut97qihR7XcLw0pBwJKgfAqljAcx9+eqyJyHunvi8gZL3DJV4OsLW+tHSVYfoC
dTd0ZfTddlufkZn6Kaxyyj/yFqlQqjl+qBbLkaE6o91TjQb+Im9A+CJ+Lxh8U33vS7JrQ+nkD/7c
cxiX+DNUdKfMI6OWYSPyqYnnaLtODMYnvnT9nmUZPJ3PceKs5gRal/9MlIh3J3/bv3PyarSk8hCw
nnpjc0Yq2SjtD/oJC5LNPNAGt1OEPyN3g0cvwtK8Kd8W7P1vBHPedB19DsZshdq4yceC0ops14lu
IEz3WPeVKhDITTiGbx5xBUHykk9pdls7QiAoguJw6gmhg2tTG5jyVk7feTrkIIvPH+TsDTh2cB0y
Xehl6dhQpYmBOqEcZqamXYEpQeB16FngHQuuy6AZ0xR2cMnshoHEsSwOr5roISPGrsv583FmgNe/
VHcN6iroXBKjngdiz5cI+XJVHqvWoLZwvpgbToT8PFsocx2VT8TmNO2096VSapkL6N4BBXD0CGiU
phfqA4Fsrlbio36dSPYHDWIJ2cYPS1ce6O+3QKQlmq6uoYhD6XMMr8VUsxIoM76nGmbJmqn3yZ63
v1bZfZb0CssuL/i+u2PRG0rGb1vgaaMZdV1xmbrTZt6dwJKyVC7Zptj7ZZXuYE/qcqjnqWlDaVg+
wOztMbH9ptztoe74ak7Ao+hvpdsBccdiBeDmFrbgpBA5wOXSlCV/CE4HmkYlk1MjGMSz1TRslrwE
2i7TMJqcBhB1F5we4X9OXTBMs7TvdxkMtWygO4ZXD+Vuh85V8iRPAaMS5csqOWjH7PU296xnBXJR
GtYtprWIu6L3x3mL95M/toFwIXxDl47R+C8B8FD5oA09RpBP4BG92akwfzWGa8pv1FubxEKin9eg
7OSu1QHC6ZiJmVIgeps1tLdPKVmF0jX5xC1JsG0VWDURw9qxkG+MEa88Wxj3N7GFQta5HERgAQZo
prqmdEZSTAirdQ/WJhbkBQ3Gi50F6Tnl8LhYfkSHOnOMYDfZDkJfhAwzpa9K/kMtmOdMqJCk/y/F
OSvqMobBOtpINcRyk4ZM633RprSfcoPtjvz7vEe6ZiJtHDwFbEWoQ8oSWjn4GRXp7pL1T41ZpNxM
bfA7AP2AvCV0HR0NZwTjdzKulOUsCPotLPssA7b4+zQqulT2s/muXADQzKI/BH8VdLNkqpyUB/WR
dpuinNSm0yYGE4w2V8YcpdiXuv/jdYIsAQ5B1Dm+kl/A32hy0KrBlWtvojyNkBAOBm0oNs91YX6q
MQjQBEb2HIRCvrmukdhXw3vAH54IacxyrYQUFp58kTknn2G2xzGI+JLlnGKIATEIPfigS/dD7IFs
qSNqeIIqPm2ZjAZ/cTjx2zVL3k01R7NasFVuSbkQdopjkdoXMOPZOJTD6tiXYoOItCGEZbmj3Ggg
2QYrOxExgMM1zYyitgJLmRTO2yrJKiPkoL1SvcCewZhDKDo9n8uUOKH7Vgv5YR0KrR7f+BSw+K1l
ObzEt6baPNyK79weZ783aish/xmRi4F3M3W8XbUIOU1H+oVSeeJjlzMA3q5Paf/dGu5e628Wfu80
gsGIAzN1sEPIykiGm0BMvSBVC1rqPPGbeM5B+F13G4Kj3NJfEI26Uos0TaR0hDu9eNrBeshCOjDE
hH1ZBnB+Fa3gM5ni3jQLJsmk3esB2TiY/JHDbQmk0wGNr0EesAi3hhIW5f1KN6MD5CQrhL1SWwYg
rmO96rPVDg7pru6cz+VTcTLmH04groFjjNVHkO9Eb9cZyQl5VUIHbKvvfy+9WRKTwFN2P4XGj5T2
/X7U8xPCWAkW6N3Wxupb/4RclyT+pVka9Cq0rvEpxbKr8Pu+5JbGzy37E+g7QysVN4EC31rpg8Ne
XUF7tHyTcPFds5BYUcHCZ++qrqcGMbJcQmf6ZsLMlskRUqf3Xfq2awuUV9eUzfzfA2ij5ljbrwYJ
7iOimwfYfuUoa6ecmmwn1L3aP5xjR3M7METoQzW84hyidAb9XtSx8omY7HeFxLkZSUdk2/AWemvk
DOUXxw9zDnkmp8KDRKq2DOOPUS+QbVCeCCnOXMtldkmxXOrYVn/57kqvTze0wKgvkDFqU1RrUL51
4EfoILSMy2JEgmHU4D5I9s0GmrJeRF6EHzU63zLufy+BHK+fjeb5iudC4xcLiw44YZFVf51S9LR1
np7JFFcZVKKxHRW2xULOqWwQYBncpETrd/KcW2rgkEs7O6TV/dA7jZJRU7ijGu37uSdVKK5GJOfR
3oRWSs8AKYkZCrvzCPx8yYWOCDwM04b8LgFjEGaJZgMaH9fjuKNtL66GpM5oKBr471iiH7Xur2Ev
Gr+002Xh5yU6SamGf9t3eDp+jhXh31sfZKi6dMhcMEGIzbj8Bz9PpJVcSpA2hw2RTjbMt11bLWo2
N0lP+77DiOXHVVF7djB1h8uMq8vv6MRaZCvjDHOqT4HD03VpXa0WCDO+i3RcRgIZ1C1iN2ow6iZq
welww7JLg0eMEZAO79RIt5kuOdXHrw3Ae28lj8J5XAv7ZrvHs1CEKzGuy1MVJ10Nvvx1Oy4xGKJZ
W9ohJnUZO5xmdfRVLbxvePpbtvDveWUIt6B8fhwBjm5T0ZyFt0zJ/4PTq6AVmFIMMz/FeccQ3oi2
M7eQwrQBCo44WCBcuP0eVlFnrpJ7QLaOLaLQk5q6C9THyU9XGK/MNfeZK8145lMZyoQngzATPHAs
+bA3r8z1bgH/juU4qhep5XZD0JyHlW4fJCCTrOusbRcn/eqF4LbYPMM/tqTdObgEyKfVbZ4pnmWn
rsez5uEs0Kg/0vjRlTNFeLFvce4T6lQwHoh1rSb0b2fvZROEYKVFbT1TCjP2WlCLwWBoPJrAFCil
Du6+/4upPyGeID6+xz5+e9jgHV6PosbPYOgqyY0rtTZB7vweNHp5fHKphqhVhZsESXwmi2v/4ubZ
DlPAC03ElOUdok+yc4OyibQaaARPcX82sKBsgXkK6WFOZAoYld7TihlNzLlHPYj6UEPX6pOw1whx
sRBXMsejh/mZrmalXtFn9jgj6SWE2S5ej09YIaau0KlSDzwGLRnc+uiyZIxE0DB+8w0nxFBgWbOG
t4oBuyrY8YHG94j0LWJfJcGrf8k/FO65jvmU4sHf0Nyxs7b4z48OlSrS82Dq26X2ZlcUPQXw/9PO
ktxR+8Y2ZQaDfWVwxVekOmkWe4mBISH1Ylrs4T6L7nCO7dHAKaCZTi5eg0pWSKRsWXNaRx2/+hBb
NgA0DrEDoKVdNZ1VZJZJhdSRr1HmWVRVnH9LgwcXNt2NlY+V4yqV4qo17zVmS5vzCC59DmvjrZQG
cbaVOxcMyNPoypWQ2h2IRryW0a+ghF672K7vQU+wxSqrraTSPe2JkM2Jy0/8rJBCQKFlPPazwH1b
XUiCa7mzFNixtlMIkoBKxcqmk5qplTN0W0OOIFl0WIqqVhyGTdbapA1maH7fkeaOMadoeFDOCO8o
PIFAPwJFbf/SjTIhQNHlaT928a0BYqDEV/jgxn47eWon/ofS6xkDbyNgZDYyWWRf67lF65AX5m5a
X2Ij3mRDe2+77Hf/l1w/e8IskApWtz60pJxpXDx1wBTTBAq9e4Q01xXD57nOPammNHh2wvKhNXn/
Qd2tPaSOW9IdH1qOPMJc4wzbzgiWrHJzwuz9apMNwS/XRPz7mjlKdfgnsu10XaPcoNZ9LtQ9iGIj
rXSmkJObmkym7RYIUyIb/mo8WZsPp3K0SibKEaXuRq31eeFRVtZcvC9vS808VAJdzpRpZMczPL2s
TfXAYy1yCor1PLl0ppjc3/P/P+LjXWPhJuCZDYGbH69JUpbyoBN1cODoxndtTM5m/mMGhkPdtB2h
jzP4VBahclUP41ikOSJnVI/50WRxuWJyB/031XJDcgIMCL//3GcGJZs1zKXK5yCa00OD5bzxc66q
ftcbOJBbPVgSHzFExG4ZMPmOuHy0tlBdxdxoxyls+MW1GHFO0kDPhXUyDXiAzeTS5Vvr0zg2NTuL
gYg4LzV1fniHtCJg+qHlX+tPWpq5vNl6G/Fw0jv6K1KAG/x+qd7jb2zYlrre72kUD4oE2aBKvrab
AiafjhAPOWw6vAFB9iT4Z5m1+pwdSYSRmJlpeUwcvLDtdZZri8rYiOi+xohV6Tp4u6RRE4RZM1MR
em6uYLtpUBO2TfFiMjKqTVSOm9exe4vYyEgJlzNRfK75kvMEWaBrBcaS9V7ua9bN8bPK6WFpVCWd
r3g5xYKcg/+8ost8RcLBr8dsEIlzUgkLkDyaAjkh0LtwtqzXy+uf4gdYhN4XjrUu7zxj6JZS3lzg
V2knUGOm7DQhMYI/ao4h07v7RcB9mrylPUjtQ6F0c1aGh4LRvM/vIWcFUDDnTQ6XyTjt7+DWC1Pq
y94YW7bStAui1NUkCYzVSEftkbMyc9JANAUJugP44l92YAU4DSWSsgrVh6TOQEX5z4JasJthxy/c
V7gbB7v3uSyfpbFbd3m/HobfCadiWHJsGPjV3h94j1YdWGp3pqWOkIIUFY34tNl9euq6/8fdhMoE
lSdtkxxWocWOXkopd66mlr9jOabsoGn+4IfRf7Ah5OnZdjF/mF2kVFgk45YCC+ohDMSOUoXNkL7m
TfaTWtW6RLqD/KW2VBMEgDId0FurB+PWtVWCQ8XtrNpDZCNRxKvTqjyOn5/9RoEHyay0aWeJo0FB
s2/dbcuH8z9AK+gX9Uea4pNGZZlYmwnW21Bsy455SMySH9kA0F1H9mTuhTE7Q2O0oUGu3K6a3ssG
+gTKzRFnWBL0wEKfA2bpDMVw0GCPR3J3XxWsLgc2Pq7L26jrINUXrYcVvw5o0uFywcFaGkd3SbOU
KWR7M4MN/Dcw2u1b+rR3WLnX2XXXjFjxskWBPhQ0vtOGKEZOstuIPNE/QZUrTCE1rnoe7x85GiI1
RYg02Y9DuhMwkcF9BTZN/vntJjc8yjAMg21qRnwKjlk1xGAZYER145HfUIXsHri/xC+HUEWbIrIQ
Oa/Ovlz0LwJeQjm9D6oDMuwILI8QDpJU10ky91rWafY7EMw+ceEMy1HvaJrw5spYSWteC3JkSDBm
xlkShrhDwzCE8axC0Fu3LAIojw3BNCZe7KSlEQdyIBBBJmrG5qK3IlEogeB3GRlt1Na9w+7Qj7R+
54mKp/WeHaz/m0q0BfrhhmfFoKgZTyXi24yZ+SLRe9mrCFWCfAR7+jhBve79ml9pkc92N9ijTt4E
vduVh9EyDsr1BQlgdTws9MIqUBZCwZ0ixu6eq1pt/PRbnJBgj/j/HboBAA7jByKERTMIoJGOd3+I
3An+21ySSE5sTdpGUfcFfF1FIueCApmzw5TgHU7cKb3il5zt6i23pgeVhKGnzYcgUItuX8x7Fxl7
Dcn5k/kmAScds8lHjA928VJYKQT2/Ie37LaWFiBbYVsAAscABAU6OyblexzfaeWlIucRaf5sk+dy
FZ9fbKN4kCH3U6fp3mgF36b4R3UNvProz3a1t2VVR4VwCmHR+/resPfTITj+LwRZYOmjrOh2X9c9
wjEIhP2vUmPqBtjaV05QbA1GjI7BERnHmjOls1d7jLNjU96EZfL4t/Vc8xHoFCuFYtzJxH5j3u84
88Uz/PLXGyGWpNid+XXHvXK5sl2VWuykQ7IyPduLMb6W19TJFqWdsZMnjPgkQa4sjDgFOSq5aJxQ
Hg6C045oQsWGcixVaR1HH3AwsuqZ+F9rjdB3zWIfXJ7FNNwwnx4Y7LH4/6GS3IecDLkWzmODQ5o+
D6HtMElddgu4LggPl7MW+d78QSoDw9x+QsRnPW37a5ST9ACANq3qqeLR7B1sxzZHh8tPQ2Qyd20y
VoJo9S3sp0g95kJLbn9MuUPcc0Cy1qzxZQmymCwm+vi0ZqSqpSWs0sRPTeOuTRuWtw0z994cYucK
/5luhZcM9+sAbdzLS/Tepgeplt7jCze+cwpvvDZQzs3RGxHof0XCOakilSnFRVJYjNV31BFJukjh
0M+kA4ZgxH1m8RO6hbwpLWqx4xc+0Z67PlYtJgB8jFv1G+snR23UKnpM1zngPxYKx4ouA9plRO4h
7Qd9l1De1SpG65+yVEO84uR/m4o9/plx1oYIlGUQfXlFamQ4Pm72S04Ia8quctuIjuOS5e+kepaP
xWmDPFPDJERHeTtMm3B2qovVZoTyIiPdzCQZl7eEM3SyhWB1LbG9ME5HOe/jinEzTtdzyoxqtSUp
0aEHAkAVCBN7nZMusDN9u8bjFumbsclGxTK52p75K/cK40wk3uCgHg1q5fyByhfXDhozyz3Xv4hB
g3Hn0VMMdf2N++wILwtAh2vpcOivCTGOAWViobFc1gpajyIYTWPBrCLkAs5Ax96gWwB6oOh/FULq
dpEYRX61Hit4TwROQeeiJcs+7t77NbE7rOQT/60CdNVBeL3mY5b4LwwUUMZI/MocHsoQsdn7IlsA
E+EFOvyIM4zA2/Mhh+wObqhsoHVhgFiV4Jat1GE2IFY2h/MR1FBQEMKclNgyoMwJC0pkPRLaFMT0
VSz8QhK5FKthzzGQJrj5HZ5xLVn4+6xHsMabbObCLvf2PZ9DJeMthaWFVAcMCLFmDBOxXRbH21sf
d2c7TOZdyes/bTFFPQFMTmcVUymU9HogdkvFM7k/ojYszU8ZCiLnGhxDF3XMlptDKWr5l9RCaa+K
lVoZWyqB2c7ORCgbKmw7NHy4fdCpAbUCE3GkYiXDfrAj4Iwk51zX5Y8zO4fsFt9QGHGBD7eWs21z
4KEl6s6QCfGgmgE7Ox9X8LwWl6ba+2P+FpsAMhc9joo2OWIK5/IlYeGJQ+7MljfhgjD+QuDr3U+E
4ZN0KVq3biypdPsbHxo2vcWMpOK2xhzrKrcXsrb7RmNtBaJBemp7Y6sZEt0IRE/MT6inPT7rOFTb
lTjebfatjfU/RQhyYrlKlzW3SC3AnosQKQKpFr+k0aCHJ4hBeCUcs+tDeW+5NXw3XzyugEktq6Uj
4czMb20RiG7uEhbORCjO6vVfJr7QIcgYrXOLS40nXdDdK1e/sOLmnombsS/o+IhZNgsBwNsdAe7O
k0KbqYGft/3oxTHk17F89WSnfLmCYvlj0rbjmfW4QkNAIAVAsfddb+oC4Hx5m4tzw6gQzn8OXas+
9Kt6cLgEYbGass4PzUIuK8Yf8dF93+rMXEsfCejGMOSKSfl6CK68rktWnaOt5FbWmudLAAbT21Qk
tQWxizH777NB0aP0PFx0zKS3Vp398Oo2y974pT3tODIeX2rxxK161BxM/rULbu+q3VP2Fn5/VC4W
4S8RW5wus/QgrIsw0s3iSZ0HGmP7OYU8PbNcpJJDVCnrs0PaqCKBDWmEjozFRSRlWxU9xoPcMry6
HOSNS/ueO8pyQOt4MDHJk3Ceg7AFMl5KHu5igy36WtylzOrbgJfFrnPod9B922UqXE8J43K0KcLA
/ZH1dKIMIUUn9m6rNjgAlLYBB9hemjcrEzRXx+KjGoy0NBvk4+cytw1lziydLmEIFzWaGn6L5IVA
mYEWVzFQP5+UDMbRcWWBaCRPwENiJMumQYMs+W3f8jD6sDqIs52FfohIM+QGQbtHmPO1CGLVya4J
+hGXJim16nu4+aYEAT8DczQiG/RBKQUugKabDseDXsXfmkb/wfwQDv1KCiE7IBKv+98R6euki64x
fs1W4IvUYm9Ms1wm+5d7ubfU1LvzcAZnXKzlZJG8SBpXf3F51S4gRzRpTijHZvMOeOR9/F2It2nT
DasGfbrzLTIkg+GfCD/J0fuyfqacIvXyKAmw05AWWBdgXSbCmxMO64EoAS+pYlzOjgOQMTV6947W
V9C4TLVkTnI8hmKoxO787GWL5+p6r7X9TVnVclkf6VtL2ZcorZ484i45bO4Mb2i7dmPYnW/IaiZO
GOh6lPsMd7jpipW5C/N182vbQaBlPW6LbV0xLpn5YbQ/qztrDWKZItuV9S+XSgs5VZW+kDuXGcTs
x/omr12Qm77Uq3G9XvkzQ1IQ5uZ5ni+rBbQN//i0s64kShBVWE0gLPJijly9IXr/dVP3bWb2V0dw
tHUoikxb5PFtMlinKn/BtHkhCvZdOObwDIkPrk44ctPcRPh8xOWOsB9okInrrfcu37Dyb+msCkOI
7s7+UQEumHgqc78mWaQwQ16a0PW7ZVSm4EvMwqSWzizrOMV7uZ5+ny7q35AsfNTLsnGnkPH3hPuC
iiKOQSEhZAPkp5WV9v6n6ls6g/nOxma3UWzY6BwdRsUIerzlHgKQWvIGLKTmwl+7NBw5RDAt8KL/
yWBUyvw/7Ue4Ul4i79tLb4ilcS/E6WOQuoRSUHj9oQoww5VXDqdy5D2wIQdX6oJlx/hiwLv9J6ZI
nJHC0SdIkuqw9llJsZs0m+YW4Wz1xRrSOvfkvLHAJ76sdB7hFiMWxK/KDS8ZfwnLPHieYMUXecol
2vtEATTZzHELgJ/kLEM0ZlIMQ1O4ocN2xhgEtSWoTU2JLClETqEWZHvJfPTkdSYxOCCHUXQuFuGT
KJ5NhDbx++NaUv7ga0bJmgy5C1C4liilCozU5SMSyxa+1Min2Lbqr3A07pOBudVNmqLDD38F9Lxj
g/nxRvwRrjhUF77MD8NKg8Gduo0DXicvBRvpc7BI+fMwNuDApX8a2w26kAasALBAdZ3Me+1qW6QI
IpQjwCYEGLt2IoRQBhV9VNiC2MvQ4Ul1mpMkq8IMgg+r/k55/xkWq5R+I5Ujfv+beRe3gX76tfSs
/Xc9tWjyMlK9+SI/WtVbx66eVHm/+dZZ0w7B2LFbKmEnA7SokDYIZN3aA7wcjSfDOdYHcxPK4Pdh
f4MWh5VRDEul1fZnymC2ECHgz0VJ/Su2+zhmJQIuVlsiainvBO7q3O2AXGvld8hZfNoEYvr4HX7X
khdBXVwaIldAuoui+RMNOn+kFFrrsLjfpsuk0MO0Gt+P1Ar+86Kg34dxarhN+viFN7q5SNSdcr0N
UyawBdQzr4Q7GJltkCySajCR0NghAF4OTn/dWc+MyVC9HvlTOmR3sMZHwe9MWKHyBKPDp7NWc8Gl
/3TKCt8nOz/1McC9K7QeD14pJZshgtI0+ajZQb0jQYkr/DIpFAj9f3lNFs99o79FQGgb1Wa5I01F
VbljE6eCelbjyg0HVyDieWRkMJUxh+3wkXX7hM/vhDh4cMtAh53owoR8JR3LnnTFJGM7w2+J74Li
WALpzvwYRAtY3eGYB2GpySESNCIBeTknCWFFQxa3DOYQ51ZHdhsh3rfdHaxQiMIaVCynH/B2WsZb
IGH7Yo8Gazf70X4ZHA1Kyp7/6GxCnQ84a15U7ZqnYSkehYQCTRI214pMdzpnwTiRTiYLxNKPUn8X
08CfsGAW7Oqxu3xMrEYVnNX4hgrFVgR09V/aFi6T9dqpdOkhg6IvgmXpsApo4RjF1n1pn56Wx11S
gvl4wKaJRro8QbVm/6ORvTEg6rgFTviUJn6coRSp400KageczIWAbhIwJsQmGExVBrC5rbA+KfO8
JGr9IMtritWy5Rde0WsFt69mQYqnq4OAmOH+BAq4ThJAPkoKwAZ/0oiv4fXE3X0aX926vC7j/xOn
dC5IM8pnp9iy9eyG4lpyhseyJX60vXITc4oLOebzza+dj0b1B2+qTRKR0b6c0sbtdpthoaEFh+yF
WIJEsZqD9HenbOMGIaIfWY8UjN7OV/RFTE6bJFzEacbsbQwBCwLOi6wi19isCs+0yd0sfRu/dgOW
Ods19pv32GCiNj55tXhBDyIcVbLw7bMiucQKYBkqZF7QSBYYvUkz03tdmAa1BgPQIl+2xa5zYdIg
vKr+sJ4b2YwQ8Ghicz0EEoUQPYabAOwvcTrWVXV2+d2EzzHH5x3D+iuXktHXSfJ3IXB7LXytHhsu
K7mj+oU1vbFa2KrluVWUSTnCTlDdLQ7yCb3jfvcUbHEL7AY2zdFN0EvhyxsmisRzppELobD8FsxW
ptxuvlKImTAwn/FHa7Wz5d00D48qL0KwUtqLLoN5s6/k2IsIIx7y3qwEUrcAgBRYV0Tyb608Xgci
bBrSNPk4wSR+DIVNlmd8GxepyiuDGGxfMpm4uFIrGPu0fy+mULKvv7TGzq2DlKdi8qP20vQz4IZt
yZlR8Ra6DILxSOjWDviPPLaBHRYJuvqRMY9iDjBCTKb6M+jEkZsg/qlfekpV86qdyDEDR47bTDle
N4QnqnvRu/rcV4CAarsJjDWpSEY0XMavuCM6tC+i9Mdr/ntiJOgNX7D7YspGpY63l1ieu+dAl+ie
qTrgnUe/0cqBbwFv0qFFsBqIym5hBNHlHjsL9OuJX1fMAGl7xDHurfVKRzEH0XqeT+kbtTXRM3Ge
PpfRO07H1tIfmwXvERqQYENuROOZrf7fHCBrqH2YQdxnXBcVeM4c7mUkVOSVtqLno4r8t4jhACwu
fn0oqIEuRofjEuiTi83qkNbBDP4hK1ZHR7+ViJOt7qbvMROWenjW9AjP4XOsb9uhFlae79kRGugi
gWYzcjpoX+yjvBRHixx+tYFAlYf8Gk5ZktBo9foy9FWmjmPB3j+x+ckdbY6dE50xESt8E+P4O1LH
ZbIIh1LPGQr3Ln+cqQ5Q6OYBlGX8XSxNAgDe+cvrbW7L3gxEY5SiSm9Jo6R7hzEUcbbTMnaqipS4
z+qxIozHtice8o6ETusLmktb4MWaY9TpWZU0e6wRNygkx1d+1EMb0fzZnEFd/k2h/7QjSwTVuUo0
6FJ7ZYMNd4cW4fAdbXbyyTKnLfhQaALdGRmxtYspmLBY+MUoEqZevIv1DbptliLblQdMYCa9bj05
EiKwHyJp848xjFaMF3x2TXGHjohfOSH7CKCavcHJnRUmT8dCsRwcF8Q421xFe5rGcoF9dwabTc0n
o5pRBpxtzKzRki+v8OCjgI51b2dOa+now8pT3GSSvraHkiAuMlmakZ65HvOmKndY2EYWMI0kfzs5
pBXVC2cjWunVgr2+s6X3dsVGAbPD+a0LmpVqLvIT9A8MHpPcgYLsOzDZAfePh9//gTDyoLA3C6zT
RdWEWRzHNSbWWQglg1xP5AqR/64IQsXf+lEF49I2gAjYw5eJKvDO4ZIYaZkskH8HQXzUK3db3E5i
/VIrnJLm6gtYUVHGOeSmUh0QHVv1gXQe9kiAzPweB6pqv1aJ/3/yGitKWvTmLp2iTu9u+prLI8yL
mFbz8GDcsFe4sCzAXy/7XCGKbuHWwPK2sWVPwE12levXuHcMAYWWJZBnoI56ljPIAdovtQmLDxFN
oXH5vj+H1DZGsWe6MD/QX52ZEGLsbIShdvWEDs2AG09bOHBWFfdcAK+XPqqg9fiBf+2zsLpmbjiJ
Ly09YdPNhvFxq/0Z9FZHgMtbcl40UbvxPTqM+NS+RFWM8LhAa1TQooTaltFlJGBAtCXESdjKjG4q
oYtiGLFE9PcJ6ZMAmmuYz1iLO6ujFjJXKkEpxY5slmGiDXifO4rUW0YMMwgz0Mm/ifAW9Tz3UeQQ
9NVxNJ/M59XCTZkkyA9zvyyck+EFcbXoawKpOU69REjTud8Nd90NjsVU9o6qetgj4FMR/+UeuShw
oZbk0/yPFIYFrbDYiLdIT8WvQjdkJigPzuq0ihRkOWNcdOJ+mHjWD9nPrKVd6+XCinqBHeQzCh9u
JdCh1druAjpj0Z8uyFMht6oTJo2XfcWpeXy8dmexy5kEX+nPHrz4td75Nbx8pak80LIzg8swtIvX
uzJDIi1dLwapVZrRw0/4qBvk4TAYIOSl36dZ0kB91hAENHNcXtQkFpjkl8OEg7fxt6G6rcqKVSsP
zkXKCo0DMH5th2rysVbR0XPJhB8S9lTunQbvqZycVucN7sRvK855+ycmyJM72AHAoX5urknCGMVz
CVdGAY5qPhkz8bYqHi2Ejc7kpQxtQytiK2v/mHHo7bcNpBk8TmkE+b74kCzm6wmlTQzumM8oK4x0
ySm6p2aseQk9SRlsPRHcqOfD1zqrN9jveQEsjPa/cz9zJFW3UoLiBHtm6IFjToPiBzFZ9dLm6LeB
DblKAYm90mhdizpEmbrNO8IyWPUJH0imC3Mm8jd15XxMRDzKVsLW1NtWUEc1rhKMkRqSDOZS2FXQ
9qySiFOUWn4vu+eWFvfWmUJ3XUPzNT+U71u59Kz0Nql2TpptqVTehkpJDlgUPCcMg4cT6GJVLKIq
z2Ux+rxri6PbhJL7oUFuOoZ0Oih+5Ov71dgH/cLkldTecooObSrJi4+pH98Qw1HBFDBU/ie4tuQ5
nDiZPr8KCxjK0OhEXp/TxEqj3eJCXBgw+JHY9jj2zb6KNWBfkDimci/eAlE+GZGkqKgGR6EKS5eq
9Pf6GHfpG/ffdDRHfdoZOwpcc8lMip6Vc+24sVx0h64ZshtA76mhI8VdtLeOiKNH5gO+NNbqDsdt
Oe+W3aFjXmBi2fHGkk8zL5d59HRVHn0iv8U3JUbbKDGNrSMgClcGxsjDjWb42uyhFt7AMkQgQsQu
voqsMJHq7nyAFoy+3ma4AHaNw+pU0JtPOrOLro1thLy9BUvE3272JzOHhEeGtaMP14BzFqNxsPvV
45/Ampf1iAAP+WlyBvrrDfCUPO86LAQprP62G8KpGH+bqPE1CvHzhoKzGlwMkZLC8J44dgAUAUMT
NC/x/4VAXVD0BB8JDbaLgAbJ1CCONvVJUZ61evgSLSqZE15+NxJoBKAxjMtOW8N3+FYmEmD+F6uk
UmqePedOqvN17x0VRx8MuaqMwc7N9m3U75vInKHfoT16yZJIXw7IViTVcQRYRJBtXOmCe5aiHydD
rBWaaXtRFMXU01lAMxwWFBYDLBPo9RiMro0XFENU0QhkpTsUHwrbvKoMPlv6Ju6aZGoo26FiQ8Np
S0fP7+FyopR58uJuzj3w2i3+4Uvzamvhi2lmKQXvk6sYnLC1qA5ZeMemLPbBDqVz3inmkTJZXQWs
oribZZY0s30mnb8YbyV3gEzsrs21yGlTvauVnxZP87tutxIBINWdo+lF0Cd47OT1JQY+ZJRjqSUk
8jeAj/3axaE4qeHepvlWdxEKdIRZUVbRR2QBeKMFQ3yETCj4lAybP0vX2aG6dvq++2F7+nBiompz
JdHHeSsbzS2AOhZXMoWV34ImCRHEb/WBi4JEBGmD3+09iX9sJFBnGMWrscWXQxjMN86FuSxUTsVI
XMcuFWWdlc0dkolI/MJsOacOYqMvdQr6sUd752SDH9COHo30EsQn/uuZfQ7FBS8eyo5h9ee+Lv9K
zxWkaTWqCdKFnK80+di9qUKONEwechzvKtU7WSKIhYczUjt+Se0XCGNK3gQ9RrsZ8+o+0FNQYfYf
0FuVATHZZr+L5SXIc9Zitz9iMezyhkU0LYyXD7JavMWAt0VEY9iJb9tT/4bH3Juhw7QORyovbz8n
pUbKcHWL4ULR14+XMTXY5V7M4ErGBq38wB4FGwq6+V8FyF0lCpmJheaRVKsSXVFZAdhNe+cFovPw
zV2zXOHQZtzMzfQTz4n+NoKnFWErLy5AaXKWbORS2VYm3TLL934bwgWipa07Xe+A4ZemVaIexPdD
AVgux59bx+/eHU5eR3sWPUZ+s6N/v198DHCF75r2dz0AzrxWodMvzd3Uwgh7LDBXtkQCxYVeIGZg
1bD2TEJeY7uy4V+xYZenHCtKnCI7rSHdp8UfvsFtthk2yUW0yGoD40bq1iCqG9vbLe3DqpSRW72m
5uG9S5iefbqIGhowKfVVQpQYpnraXEYosODa6dM9ipK+ENCgVjpAJBHf4R8pGyotkPT15DxT5J9V
dH3oaIT+uHpIzbKyT/KVdi2EBsGtgk5Qy3EYdAUicxUnklICp+TWaL7b9Qcf2BnUtev0sEGixALy
MHFwjhY3EtjlEGaxb9K0ENwZh9y29A1GDZqQxYnapklKbUTK0pkKsWwAPbl7TLVFmuym856BEotE
JvOMbiHsxamqKLbXlBDhSv464jpsV0Gkr239nARhSMCSCbPlx7X+glsIeGs6R1FZRRfOgVfre2u6
Ac1kq7DCBOz/+a28zWNjeoeVH2jkjThGPyWfu5Fld2oxgx9RNHqkT7BPyZtfChi2x6MOQG+4qBnu
TX2dcpvSi2eY6nKqQ5oo3JRpeogbiibG4HnB4oIrqwHyHDjWB+7SWYGUOCQkVWxoUiDECkE1YVic
vUgX4v4lUkjphkJBL3TL6YBHGaLiZdvpca9ujR1EnCpSETArtBxmouBRLx1P5o76YRvnGdIpRK9n
MeR1HW/kv1NdHLHRFa24JV8p16eF2GVNI465FpE4+aumMPgoqZvHpu6oBngQcWCY2jAp5fOMa/2p
6Lytinp0IH/n+i0KXONqePwjm0S24Jrd3vmrARuIw4FXl95pBkcISukkEojFmoB5fOpH3er1WuTd
ncPeE+ud2021SymDpyw/49L/NF5roq0uzZM6iFASnWXTMXlZJHYKp8qCcY40kClroXTU69Vj6/5t
auWEGZjWxqrpF7Ke7yijDnJAUbT/bUTAuntfR4UbbMZ8cXOfaB9rcrckzCQpwhPc0tlRj1YaXHQD
9uOpEQ+yuVliAX11OXdFWm3etV58g+Xg3XOfsEBGiLf7L+8rakTqDYTRt1ooAOw5GK6OgmT7DKgi
d/7ftOF+8uuP5QmCOnT9zZFULA1G5N5fbXZK+19q7OTCVeXtoytZHNbV1olkX4utXfDtzWEUt7A0
xmHO8ougiiu9FCtwabU6rbfPaifhFO25m5cEWq07I8szqn06PRF+2o/yXOTC4Sk5AALQh5VDH56h
HUslVYCUEk44hUQ1q7BXN27PDvlY4lxYpHl3hrc1O+ELNyOqvexu1H40GU7vMjSeGielITSJT7nt
+0Dw7dKksI9xf4SgQ+iFcMW9zK7iGMnfi7rtsmnwvkHAm1EcR6wTgvty5A/6BX6V7/ep8+gqwzjl
19etTJkd4iOKAQavP3jBwwH5KR34actMwZcXthqm42jcfHxA6Hv8Y1X8lpshLHY0bN6/Oc2bG+tl
g09fzkCMcSmFInuCtAQ1hH25wOCu3VsaBf6b7ITJS/aY9csBHNSf7N6r0LuOCrL2rLPh+TMXiLvr
dmOGYQ/LWICUfjixbT83bk3mAN1Sp8USlzcPksnDn1J+3wBsgvUzE1ClZpu/Pr2lowKcF/wcGIf7
nY9x+rHPWJ/03vxFb4R+HNMsmsS1WswavwCw42vTahHkkKBdWLgXL27BzcCglqJSw9rwU4AGEnes
nxh57NywTgsiEVN1lfjrx5gsaltGUP9//gpO9ZpqlbUFX6VbTsxm8ti+oX5dVRT6z1Mu6ZMtswzw
8cJSSyCZmoHrIsT+8OiaHEMEYCFpGXqD7r+6R0vvh0KI/Pm8m6xLUL3RjWT3pRtX2zRq2w7LbmdQ
HG1OfzEKJnQJXpwa5muFcQbA44GoJdLLbVkgrX4dvcWIvKO6KyHcdgdW7XuPjyfjuz0fx4D0fw7t
odLzOVFz8q8ALAaniZBLdKxOpT+CqQ/2veG6ko6XhQ/vJ/55/gG01i75C0YmDhwfftw+7aEh3Mb0
AydKOZd2MdUqKJ6L1b8HI2rzqUHrv91iv1yWksTBpTJ6CXCaQJqSxLhSfrurpM2DHXeOFVdLn4VU
SJi4DSudbfCMNG+OohfHU+wWigCNwnLHfmkveAN0BbBU3aVxvyI/d5cefWP/yLKLAMv+CmaxnA6c
CZQVQCM8W80unIFMLH7Pg1QG/laKGwmQ0lKwj1qMMK8c6foKUXIybru83EK7rSTejK/rUKG9FXnW
xah55wml+z5jFnMn7mEzLb2MZAL95ns4WmV2z8uIp8nYMrpBMw+q9zLCzt5uxpsgV5o3dgbKCspa
IQ9uBSB/0NECzVQSm2Y8JQJefJ76f6UzifMFGfoMAGLwS5Q4/r+x6FyQDZrYcGHmIiVvtFVoFixW
Tv2qnaHElMVuBldYM+0+4qmF9eXg8LQFHaWzYJibwkmCNjh0RIAM8swUOV8olFmS/Dj+/5yKDuIT
kKdPqO21XRn/iVZSE55LNd3KWCfKB0NfLjCSIWOsjNqQUUD724/kWjoRRQbcCpKE7/OKuz2wgAPs
AjUfCHW7m8fKvzdA0Rvpth67k6SeX7EBMvSrbHxRP/OEDqdWgtipw5PShYuRs4ca1k6wBtKC8Ip+
5soITUFBEo19zJu/m69rBU9/gaRBrYmdkSQMg0VnES9a00tUZDHuICGAT/y6S7fIyuGE7IVVYMBY
Y4/ndCGYztJ1Iv47JXnWAppLVWb5EfiauvxHo8dzFjRQtNWcpuH+f6urzLzIDx//lRBUm/gDp4wx
oXUHaq66ohnv7joHcljmmj6/Y7fSxZBemHgO2ew4fS3DzQ0+rB1TIvTnClHD6ONgM6gulKWwhWTB
LQtqEpRZ12U0XzApuPgQ9yL1DzPPXt/tHJrEJi22lLlz/JwwPR4OIE3u73z7oirx4WxBJitA6+YB
0QuYtrPXitOf9+8UjW2+eN4mfmJKmqdGbVOUcb18IIO67oHwvqzFeIOWQXFi/u0N8G3WOUS235jM
0/QjQWZtnESQie5tXvBt6p3SzDV8h34L+c7a8SFCAiCZ6lsd5DL9jK4vHlWTjEgKfY5Cvt6A/6kj
0zlYR7795/LQf7uh718nH6De0Sxs8AyTqeke4g2i6bRCsgPtm46O3I6JC2W4/WCdohikizIbrLSj
Wqr/TkHrgpqx3o7Qpv8ywqcLSYGsqYcb2ouf1E5KFruPythMOqU1/COnOz2m4EHHglY6Opb9/FvD
AFCApR7Fx69SBb+GN+wfX6R/9KgkcI1j+R6iz3RrlrNBQpVZ5pe491973BOTMK4OOlHLduvDT2TL
vlpau7LjfrWj/FRry0V0lQ9Tpfq9myigR+ktrc2lgaFi++aMcc7FwV+xIFP4l1VSzGjE6khBignm
yIGmJtce80CYdq78jwUAku06Cr+UA47wqh3Jxr915lxvecgtPOR5ojh6B5opix7hqp/DcmK8Hni+
e6sf/cWNGjRAFk8WOGVHbmh1OUZBJ7JmT7E9ffsi0MN73a0VLEU10PRredd1kBnC7EvXHfGzKBam
NFXJwnPRId/QiFIze7tisKW9xRMmrDax9nk35G0R8KsrpZBC9sLrd7ShoqWi42xM8/JUG6ZpVf7b
5RvB31vJIy12jtkEf/gkhv+xwrhH5rUFZHcZsWmBdrjtyfap9CsHhv+whYXqWLDPVxPxjDQiKlAV
Vg981F/vBvo2bIpPrtXPpuAcybjC2MNCN9WEwh8rln8HdzD00ZtPmFZVsPK0Nri+2Inp02n/hL/k
hDQMzUu7iI33HDVIrJ2L6KaoZshG8/9jvA3vDkSD/+uU25HuXrxCOaRq8iyG9kR9Uizu5oFoZinl
KOUvn/kb0xMRbJe1dk3WcwHI2z9rXY81Bzv7RCPlCnqEm91dXekprUyOFteSaBm57DaTbhHMZR5C
s+uJvRNYcbGQQQH9MDsUSHTtmehOknmRDwDLh8w2Uyxyabvwq6O4LTNm5uQhXKHhv2RXo/QiYXcN
1GUsmcdKYzY5G91bdJAKoXpreozaEXwi/qEntac8JybwuGXYgUU3wf/ttjHQRpHiQjP2dBpFExou
GjAemAmD3BDgnzTLq5CDG1u7+Qf9YI5T4A9Om7de1crbbJycnJKpF4xRPiTmI2kGgDhxuehL6Z5u
9+qqPnKZIzzCRgfR4ENNVY8bW485OZNPf5P/Ikq1GYXC+C1RJ2rZ4m1KRBjzCLzLClh3pd+QQ4F3
2IMORKGh3mQP/zaauy4Y/t5bEeoJ/h0U4ANrnlOwgRUb5kKUuciH48wV9F22W58DuwYZIVOEMCrL
kFm10sp7rngGimbd3mDMoYVxgnYhR18Zyo6t+AoUUjq4pOSlSZtI0jFxrMu37Gg/RXTEmnF0ozrS
1XeKoTQ/PWYX2XkJBEmvNhEXhPL2JaZiynhCqsLw5XY2ZGeJFRdtgzp0AvmivT+ANy9rCL0Y/9ce
iXDx4+suV2SlqhmDemH5A3McMYzRUt72TSDeVJIpg+9kvl6s9hx5dbLF7XvRPaT0iaH3HggNF1p5
TJRG6ZM1mc7rzlc7CWAfXoYeDhxXwb5EJ6TT1tFHp/Gwu2KITiuqgT6JqLHY8M+1XZx2O1vFoajc
WOSy8gEC1kbyhD86pvYvHgZWmRoKiRnUs2VOhdyWSbEvQ/6+nJpzqbiy7uYx/WN2Xs9Tz08e/9uE
AUVTOub2h1DWRJCQjFVaOq9bazTkgnbHrnY4gB09d65GZj4u/mJJ5OzVoRyVZZQ4CKBAz5g4i8Lr
rbYkVrf3cv0zKWKbb7vHLAd6P6EKgaJcFdK9bZfqd446fdZSVlFGjX1s920MFnGE3noYLCkQNXJ2
k/qk3PybAJ4kNl4Fo9bHzDZUUblKqYApAsDFtz8IqufvDJKZ2Kbdw6L21HsmWTJhnoKtzpA+2jOA
osyESuPWdh/nWUcZoy0TmTYyzNKEIYvDNapZ9PLt5Jl/DcysyLUgL1uJl1fZfHdXQJNNDPejgERQ
lEUvIbHdJ4Q768o3gDGrDq1xdrZHR95te+1DQZParCcKSn66Y3AG+hCiAzjaErD+uw48Pqtkblwn
1OxR+YAMSo/umTsnp6ZMAu34Pv0Pk9Kao+J89Ur3vGeW2z/nmA58KSbc03kgMoRF4xovy2qd+UkJ
ulh4F1d4/DG2cu7eDiViI6YbyN1MLxioKx+aP+eLNiGotvaMklAqucpznwSOWN94ewuBMQBFfyO9
o9z4YLVAa1rz+ZahNnbpDd754BLGTXoEE6rAefdLo3Va7MKRTAngu89iWJpAD7zE7cYLPFYq4F0q
WLbo5jrj821lN+RLiZH/WMhy7Ld5XwvG+49j+rNDwGXtf5AVFIgtmBDREjTmufIMJImrcINtEaCd
OhvXjQ9yDqxTSDDZzMGqInSa+ysUh6uirs6KOQ6iKkr2frEuH+dHCBfQWoRafBCmQMywFf8gmH44
xzN3czlsGKuB0ObkECRsQahv5BkyCisFwr8F+vJSCmi3uK6y1TotZw5A2cg86HyMxvoiQys7o5lj
r8fdHfMJ05/dmrgtxVDZVnsocJAiLdxmlVlvAaHxvFiWBgdgdYu5JNQOWhHujAZAl7vIwTyEJBGB
dTlyZXuKr29oWllpIBqVv2oCm3UTArJgKyvS1Rm4ShZk6QDUa9eUDcX9jvcxT/QCjvtawz9SSyAa
TiNogRyGUL4NZzzeuJKEGlWodDnHC+0hKfvvcNfuTg1b8IAxq0I5P7nNkyf+1aCHGcBc5by2dcNY
QPuVksA/bG8GMkYI2XAALbct1HYQx5F+q3AmStEk+3+S0/E3fp9++a767zUYVyACOwunnjGr3VlU
yuWQlioYvKcFMAKg8hoEqCql+7YT8hqSB0cESILBmHB4IILMqwjdq2lsi1sws79iS7CbOX+0PZL9
ktGF1sG5TL37dgfLNU+K98zVjucjZVG3evGU58liIF4pf4xucAAezbqLyKCpFqoXp0e4SIXLxxJ5
I755NlmOkEkPt0aueVsP0oumxUS3KaN4g4jt5oRllgE30CXpBFbtykRheFMDt//98ZNGlgk7eJWZ
D7slOPCYdELuM36rN6aeyXOwo+phIKz7d4XCFZuPxgPus9jVdF1vKnCLtXOIdra07Mz1vnCOWN2S
RTfgt563/XrHlhmhO2qkZLTgkH2cnehIqYltZtEAlKOiEKTM84E3yYWNSx2pk7r8sSdfuOVzemXX
aY3qvApGVEgaDHXBzQDamt2B2XzZutCJdyr17JZhL9X4WfG7Z7PXKp6x+7oIXs0xAF2VvmOuN+u0
sAzqdGgjlpbmyHPBV4wSGB5MpZsuG+NoCPff4ijysgLsKakaNymGUkqeDv2bIgHIXxmhuz8gzzrT
cxsx5ZeJE3qBOYi9+QWCR+PAEQjBzsDOy8DqBYqIkmxWuh+Q4Tfe2/qcrrBbRueZNILlSJ9dx6tY
iVYgSbn6HJa/x0B66lZUkMXlMQ5SHmdDHxoWHj0NcgrLnfPEynhmAEo4ctnC72A1lpknvzxfp4Gr
Had9IRbYgDysKlyFFVOpMTIXNoZs0pmlpI/xMzQ66wcKa+blBPR68wSZNHiQElpw1WaTXowzqku+
PkREPtBagg0D/QM/h3YloN6co/kgVnolAaa2j1Gb2mr8m2ZAp5ZV3b6zsFM+ZeGQH9UFNcnjJXYN
m6bgcTrhx2eKkfq6MBSU88IMwKHb9D97gE4Q70zGKk8iP+kbs7TZO5f/6SOWeLjzPDG5/lvniPnJ
hPkm8rVtCHhzO8Su+aemG+g0nKX2CF1saG56XWF4H5gwkR7l0a70wd/0glH+HkJ9nRDKt+qrg59C
KvrkJZ5F4dUrnmZ2uD7vyYsLjZ1D6D3tuNyL2UdBDGXmI7vdoWo/asv+s38wJ9TOq34opX5Dlklq
I0ya67RIzvH/mIB4MEDcxE9g86kFgRBvrwzr+fchpiG1/D+iHjI8Xt4LtwlP3P4MlBjA5U1rMut1
KSio7xAIKEIP0DnhgVEb85JAbpFh30SLv8ZNgfPunEFPpjob6Z+TZSRghsd9iXcPSAKU+g1indS2
N571d8bR7/35ooxYF/t8ffRXCFQMeowiSP076BXZ+xnyhCq+XzMjsDHGhVTSWHoTrJZ1jIgyi8yU
A3dQ8rnqTm/cG4SxCgsfOykZ+tFNZhHFDdK0rirSeowH7PiKDoBRKYPY0gigNtG7x9pB+OXsgxfm
LyXaPWfJxGf2fHBdd1lgVOpPvKnC1rNftnURANkha5Fhm2s5jQN86drzH+lrzvS4pUF3Y5LnSmc4
/loVgQCyQ6iAMH6nMUJhA0FqgNm8uFpctX6uXfLJSdfi4Q0j7PiiDIa346DzsHxxGRh7qD2+Vl6c
PCpy62yu/8N8f08dsD1+Ck9rbowzBWGM+mOqGl/LymPuJZKD0ELCpEAeXnK6IhnrzHoOlQceYxWx
6Gqpcbi1o/0QAG3DwjMZUQCYCTXOl4dxvDkiLeqRbMMrB7jKM6ex6GvGsMocCFjQsTFdUnCkNKpE
SLd17ZpvStPg+fxftg+0035y4l3HdXZW4WCK2ajnpS0lcQ7sv5ePrlTcGs4fnjS/rP32z3FYZ0Pq
I7D3OrQ5qWdP9/3QMdIsuFDcG46DPiXf2TH/gf/Ngctl/APAcBuEv+k+Rd092ZX5ZcadtXG9xK2E
BQhKhHBITMiEt+zL1VGPyDH+QhRO1LJBtGTC1UFXhHH662sIcDFfeDkbCzCNySwcBS+wBbB/jsBJ
QbJ0QRmB49UzrHotu7yE3gQD+7nChlqRnz89Nb1buCmk/ILJ41yPeYiOcS6WbVE2HjhmnfKrbhKq
PDbwW1rLQqlU7cyCqewRd3bHw4pJJaOQkiYVKA/zmZVqZuGdwt37cDoS2WkuUXOQtCyY6jZ5Q3f2
vJk5yevefHCp8Okj4o9hd2ttJUo6GGqA5xpGJtFoQvidrzzrH/vcv6vswFx2fbFvZPWhksv1mJW6
lHv1rkK0wHToHW9l6wKR7hklh4sqV51vTPC3ArYCb9bf3RcgclTVkTj10RglIcBRSUffREnclpIl
AwOtuen9verG8UWHhWgiZCQHzsirVt1MFB1TikqdKZoRlwymNkcsLiWKIPP5uuihdqySyJRDL4t6
Dypyb45JlJKQNZYkAFP2r5Cbig3z+xcWv/KtdAKcPzYjaiFqGdQ+PBx1u4XK8PS5GOoAIwgDjJNR
pjX0FrXwtu4C5tqpG+VPq/dnH0G5WVTDM1yzU55ft3bgmkMl7xHFxkQg1S/oVrljsUvYQBjc2SFJ
bdVIdJ1v2GR2v102IXJbgpuKe1GXTfp0g60iiVbsc36Dj3rmTkaVCRkb/Yzg/khkNjjbrFQeH58z
++QbtvoffexbynBdqfZrE8kuijabEh/lzicy49UFwkUmQVIOU1ZB9nxcrXtAjjjnCgOiLVyxOW2b
LI9/kHveygpBdoO54GEz6mCbc7MLQgC2/VdECSONj096QJBASfRHaD0eR/QWrlgmcTRR1u77g5xJ
aHDIEiupZWPObFdRb/RUUnPIMxmcrZz1CStBODbDOi7VhuVPoy228OyiOwv4AV+CIqmqtZ4DzI6u
jFbU/SBkAjTjkPc1svdGzL/wTFZGoFYBI2Cu/05MTPInELGvWmztIg3eicmqVW+cyPKRwIYIZi09
mt1sPqvWkynsNbLyF7frtMlG5+rcWWVYk1EkgV/fu5dxk8Ebm1xtECI3fGBkMgSdWiV9DwgzUBzn
aYNNns53QqXq5XH6S6JxXI4P6GAdy0Pb4841oI3x9JYLq4tleSwF3Bh+aTFHcJvpVlt0U0wIbUjT
cHPQa3uIcAxYj0kYFesqEbZehyvBXO5L50dzRI3A5lntVMwizd8VnAJR31nhph5BjnEBlttQZfHJ
11t1kx3+0iFmk3J+6UJOrvlSDHgXxTyYqq1oatbRO46nEB240mWtiGxPARy5HNJUQt87/+hy14Af
fLP12Qn6n0rikqhjCNiKpgZR3FQ4lUqh0Z39ANbAWFRYkvg0Hp0Ee3fztiLf3CrX3w7OiDf7oMjD
OhP9kNX5ZQw6JqIDRlplHMr3PfkmZFExstbb4AC1qWW/WP8hlumLrQNYMTK0PiBEFv2QopellQ1C
jiHYCY1Mfa7yms1QFSqZSHO3pc/5/hav+K0ijG5370I7jLggjv108eu7I2Na1PqMBw3paKzsOyzk
GJRo024slsd5g/4Plxl3/an/e8jJCuTxoBwLbtqJQ5cWZT2yodOGUaTde/jqD9hntye7yGyGwA50
WnzXEfgxvJCj+3GA8kdYfnPb7JsCYLP8ySkAnZDtRdOS+2lOefunH/B7f+ihRvTe5PtpMMpTugZc
uyopldS0Af3tqHHE2bZvv2JDM5JgLOAi2g0zgo42bSFeZsw1GbZs5jtVL3SfM4xAnEpjl9VsgDIM
5R0/qOiqVV42+OVzulhbKsVdYkbKSzuWlHlLhTfgSNNRIcafrL0erOzD1z16Y17A0keRi9uAaXpz
F/sMHbULXN4E0mU3J76FcQdpPUuYNzWDc0B8yMlwUJ80/W5zR0fYLx2LxNTbetV3G1F06TwqqtUL
5F2xQ/QNuxkQZa7oqrfOBgAVFfIs1ZXVUUrMwH/dC6dAfFqa5VuocjzSO5B89J1BwDFl3TDELydc
l5wAuea+Dt+KO3oGAMfUIrzI3vYtB1wg9+s861fGz8HEp+ey6Wu3jAaehwdIt8PhlOxWZvb4BH2O
TUD0GW0F35TSEu6oL7xy+Ocn1Vd8ytjuVZvZFDDNslXT7KS5tl6EsWUB8FxhkULJdUWDZSNJEstk
n3UGfiFVEg5CnLpDTAXYchHDjN11AtO0iT+96Lt2JDmAX2kGCu888QVOnI5UcLzivnmc3E+wznxb
eyjmmZU9E64GAV8E4vT1GZlZVMHkD4CvvdOsVkK+yqq5bKVlkBrqaA5d8ng562DNEKiRe1/vufkT
H300J1eZwip2D7rNpBWqSbbXid5kmqeLgoJqBFxdp9hLhSs13lO2Ujlk0NvE8mEQT6ighed6b0Ku
2pc6pk4Y95axBi10C8kpvp4I1lqdmSoRDIzd3pMIFV42gkLnRVak4syQLo4WHv7ZYXRmu/VZu6LN
c5UKIKocZUbwjX6k3jrml4LhhOt0XKeYIZiHHBGzaXk0LrTPU+7PZ/c1AFlgpWYg4BA/MMTqTYFn
Bk7UB/CHZsLVnG6wrZQx3CbFveigcTrGpDqOlxEmJOfjr2VDHFdNlW6ii8bx0uSC+ese/lU6uDnN
COr916QAoaN/D1pTPQRTwGA8e+wEstdOrKRHMatQwsvv1bONbAwiCjPKA0x9SbIfL912moFuOg2T
Pa2/7pePIIQSxfIzf517QD8B8n4uIxoMxd5hU+BEaGMntI0mS/gT29/vxRbQTonq1uUm1HLWCd4B
WQS1nIWM/Qa/vElESIkgPkLUxDaEQlpLZF5sih44v//QWdd94MBdlkA5u+qdptv0b2z6UTzXV6z5
3c2P61dJxbAbxexZm7bWtnHuImls5B1y5+mSY2KyXpJTCZoBQfaFI236g33FaK1MtZCfzo2dCA4k
U3hf6e9k+sKJexGceW4zCZTDYHyhqLTmyP+/uxBt7jEG1EviT8dmZSpubKCxzXI21e/7Eao2Ganq
eOV+4abarpnpzoGK1HhaaO6jksuNh/nky8aHA8QnJSKr2zpDX4uNbvkjPNQPwiEiNocrFo/cMVFg
E+CtaKzOhFK+lxiVnaZtbEmg/x6Nv7fXQCW7n4rqC3jIQWP9ehUAh0MAsSSrSmVVnMOf8mCm6GK0
qDPbXVNwP0b15B6HV8VgH/9g4ne6ZJAhkXL/gP+XEuDH5lOwPGTLKVjYdK9W+vYg7wcS1XEmCvvy
nbwAF93ozNWmx9jkcNT0MMN++03BdzhWxqIzeDbysryB0TJqaZl4PI5Zxdr9/S/GMzuv+xSJwTvD
WQAImSPYGRVYSXK8ivdglhBteHBmV1Fc88LD0PYu592r6CGxwR5obD5h2+9GMMmmDSEg53f6wCD6
VN7LaNDcNc9Kf5Tbyax7GbXQuTUmVto8tav9sWQc0BUI5Ad0Ib9TpqZh5oYMKvhrBzKmO7u+hCp4
U+OEfsKAcKgRShYTgTUcK1gPucpdTnlzvm4vQhmLOdXkI96iF+CbDsCt72pO2ImSz03TC4ZXlmLR
lAjb0wI6q3y50hjzvQOMGQ1OhlV2QBdXv91uokTR9W6r47BPO8SmiPOumcy0Ka+Vp16rpgBzwuef
/v02+nCFG8X+8ISBMYD+d7hZSZa9zi/Q8rSV44gBt16uz/ryrNGu9SEM2cFo8ZaaXqnQuHukAYSO
8vmDS8jnumDlA+L42IkS4V7/Nx48k4W4bdl4OqLeEmg5kZoY4N0HT+YfRjVaquKWn50q98IYZTv7
Uo1PeptljbB+pBi1jiiWaG89R1NPIXl148jZECDmzXt1Pu0VNyTaFszFmjq4h0bQFDtgVTeKmTEU
idRWb7bN46mzehwUeY5AdPZJZFiK59HJOnYhX+vKkqLopSFP5HjG5c1CxJ9s2o8aKrjJ/qSFblBm
ElY5ZrE7uvk5UVsD6kOGK0akQg8wg9Y11Xk+F63DV8VNwokf0JqIljCn8VRivZSg0/d+PIZFjVfr
axqAoNaR1Drb9AUzft34tUbk96zb5nBeuHD6fdjmmBORe8nRCgiYDCk7xnjp2gFfC8cFF8NiFLl+
mGXEwj+1RFkDyLNaELVbJjEPQJZVXxzpLut+53UCPEVsG0e0QDlRKBiG398k9mL0eQvXHp2c3+KP
2iFKB37w/PFckSd2lVi1EfgCGBn4S8KktHRkfmd2yPsIDfx3u8BolvaMxDsU4kynUdBCeq7dnHyz
JwS5pQuI/vxoEOOs5Mc9O6SNQ0pvI/IWdK+J4CUB3rXOIWfujR3Xs97kMihR0vPaRT6oMYoVtgtE
XPnfgiMhXyJJb31l+KLovVHqWekpGoZLkwtVZ/AkoNeaA9sQKWRwQWMJudZOA2kkbBRYazSAOUjB
CqcsXKFSN2Cll/ADTL9bXooMVA18KePbn3mp111OVjqVRGdIJ78iZOYzwwRKZY3h9wBV7OjuGSPe
gwJhVLfRZ2zoTxr4x8zF8TE/x1ypHpKICKY1cEq+0vHZQNlTaU/aNanOt+K48L2QptVt1KMr0Ub+
GoY7pX5ThoDVaPx2/6Ii1PThg3ump9KgnJ3+7KQ8fmU5S1cqbvNTD/0IVmxm7jUNoH20G7BjjtLQ
K0R+YoSVfupLsj352e45XtbGjrQAY3PMq2pL4oXG5cDN0AKOCrpQYwfB0vM1Znb0uzJn3UYP8SLu
WDxabHRzXInjUErgDmcJiQbk9yc//F+pCWrursNY5yh1S35KgkMk8IYMCN42SgYESuZdV7BkcQ4n
y9JPS1J8q52S7gXDHAICKC3SX6H2i4JvdzRr8DldNCYxkCmdEQS34DDtt9HyXMCCdL23rUC+E96l
6l878Av1P2l5aAxAWEI24zrcvKwmuE7zlFxTr8uHudLDPQC+yG3MV2Q0edTR/yzIiysgGdF6yJij
ruo1hXcGMSttsW+aWkP/iw3X8x9MLIUkevb/myGCmsXdzZevScmByiiCEJ29qgzwfe90eaqH6CNF
8Afp09ZBz02FBvjPFOdCQCmt97X6oVjEB0eUtQPfkhk6Lt+EY8BzpYIkfgizH0BcN0pBrHpa5rCp
zLD9OwSPA29Jq/S1XvUPiXDSQCrMXDZFFJ7kLeGgfK9ebmZuE6BJ31NRSv/FoiyA+DNs0PQI/qjV
9iV/KXLnCOBus2KeHUxMA4RvyDXpJvN6eXsXETdQYwpKDccvi8ToZHmOf8UrhZ15PQ9QHYmet6wJ
swym4gTbdOdNY2oPzBubOA5PjWtLge7qZInMd1Ux4oaUqSoGQeCzyfE2jYi7Sjo5CREPvZeoDlbN
X1V7KjJpN3LKrhryGJvLVupXAC2+Z0igt+ms7Jqy0zibDIFJbQvtNtIGdFJQeq2OqJcbuIfA7Ea5
EgPBBp90zHPmtI0kzudBc81NWizNwWScdHhHBHf9iNwTGSjqJ8wT4k93V6d6RF16pcSHvB7koTzB
D0NktjIi/1f2+UeGEY4/OftAIJOxuOFeUSz3wWTYsaVVDiigHSmQrCiKarE0rWtkjIGLAvwEnN2Y
rQJaMpdJHNTzXm0QC/6Iq75Txin7EYdNN+KoeS4qmvaQ
`protect end_protected
