-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
k7bc7mMSrQrE9Gl6ISTjh+0wn+tbVlv/ZTncyw+85ZhPSc0SnN8DF2+9ckYAGA3vR14vy2IWtENi
Erz/GnptyEaCxBiziNaUckI0/MqtWbI96YfDTT7XVC80V/FFtO8b4hPrMO2NLC8fOhEEKaO2c88i
QXFspkedaJgGV78Sv22N+xdzf8kQQ/9nglE93qSLsxImjiHglPa+0WdB3lyBx169FoePu6iNTbqU
y9s3gOpkhyC2fgg+RHL+a2MMyf72BIspHvnxT8H0Ll33gDsZm/VBAthC+HskEMYqWV0ngatReH0w
d8n05idRZj12TRBrtSMOs4Us8BIP66UUYq5quA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35744)
`protect data_block
5So2SjWXQLlkF8NGDJb8X75yayBB2fQ7HFEpxa0sfJpmDoz2/uHMQqM63RMMmHtqofTzOqzYQx1R
/nqQYI8vDUlQc2RDkPZj6b36eMbLp8jUz5MKI+99iUuZM6Bc6KvzrphjSDFost2aC0ZKiOYll29S
ryZkVBQ98zoU9hCqxRgRPecmyazow7KXJKsAz/uDjzGkNgUZd46C7PS6jmm5G+35p3ad/GoD0I7y
Z9eC18CoC9WF5+T3OvAiyqi0ferVUpRk/cZYGlXJn7PURwxIjAlMj3mglgoGnE7/HfRHOB10B4Pe
kVQTBSTxhBngbFelkMjXwFzOnUH5BBiimzkS6GTGlbbstb8jJhvFaDOiFIhcCb5RmjHPDiLBwIZm
6b7zCLW2EAgEgv+MlkLp8XQgdcG8SeFknXwoH0hkKWZRXJE3SwjKznHQ0BqEuXADFplFchJJj5As
NYjeO7cWN9VhnZk+4/CDc4z/HqJTR4sQRyBHo+xfhwsnZnCWDqjSjrMXenNRAmJVxfbQgo2OS8II
7xPRxEbimjoZciT41J2iM3q6mirhkDASifw85SIR4wfY/OvbGThnp51bZ18LDJcZzEnuyzhqKTmu
IWLZEdP4MbVtS8yJhYMMW1M5zH4OdlESUH5uOOXB+39P07iYWbVd5cmxwFGg8hVyjEZsogVb1/7N
2XopTFLv4YBw1m8auwdB3kbxi9sb3R3CFIk5uDyV8fhKC0OFeobls1XvTzcFGV0PhQ6kxFd6sf4G
YqYWKssLity2vh8yOQKZ1fO3G/7NTkzrTVD0QL6CobIJbe6LrRULkWty9ZaJ/dbybMauk2lYsuCz
YvUC73cD2ujiEHVYglOIe/WbRdVL4iQ0MAfSyl3HA3uMuyeLuomW0F1iFeHTjS39rAU8EhVgI1h2
8iRua6ZgyXp0qa4K71FhbOT7LLUQvJtcNXQ3gExBF+HS5Tvycc/zeeN1qIhNjRGBlrnnBptskp3q
FdbuZYr2kTFjHpO7J6uTx0rbsJTO6nVDfiZI4vdvPswvU+uhD8eh9qp+AJpZEb2jCJlPtagqaWZg
IWMurRllGSGuBLJWI7qweikAnSatC6qhWlOY2cQWgCenuQQSG2zvfEHYPx0ObMC5X6qMlRk8uEU2
1Y05VqVCMdpjRWHmuLpJPYnivO4g4/LTzFUaS45s1N39noXwFHMZ0dIkClmiPQmnYzxTBsRyue6P
afEbrTpFXGII/Frab/Rc8i7esjCtZFfaOYrNBgXraFc9XOJiRxiG7PS9yzDhKO4P8QE15EHgU1sW
I8IYOKR67PtyjC2OLWnsAbFi89RD38BBq2fNQvDTfJRM8N6PLbbSqVEa8sCdjB+GdQlX2eysgPH5
HPx1VhRWLlqJa1OfvR1KF8Rte8qo8W8hHD1TZgXgjlABNzNZLe6n1rlAafgvczVTdsypZaYn1Q2r
yVeQlUE4aWf12u6CDg5DJ0S6m1QJJeYc1P4p6BcahYRszplsxubjOSegL78rGgT6b9jsv0HNShU8
NL/u/GNByHOthT0VPDC0L6fkP0U6a1FqplOV/w2gorgGz9pjYJTrOdkaolLCQkt1kb9GZO89ryjI
kGGmG9alAmZ9goeWdsvX2GfpQ28tMyMR+sourFyOQDLCQ9A92N+dFhjqGmjZ1kQBY/oNRbVtH7yI
3t6CjIq1m9yAs52sIOMPvSwFz5LpnDCrZ1FP3uXaNlIHLILasO+krcQG+PXdhzV6chLebgpAAmPT
3XRdD5ghwBC71TxVEFRwNLMJ5lRVdbf0GtSqeF9dFouH8wJj/WIvRdrzREfhB4efhCBnq4vqZXPz
u+U0789nboNYMkZO/4dpkWnsjH95+f/idQKyZ1YqWQ0lLXkzE130eAO/xIDoEGK+juv8Pide/bCE
LxWOBOZrc2/+UAU44SDQ49s97yCfT5uKJGgBG/6feL5O++goBx8vIAvkxLdalwYtDELv7kelTY9X
I21OYgPJfa5Anjnlvs8MXY6PYlby/hOCaMVvtW3dRboBLugnpLvrvDU9PdPXhkv9AxwVHaWHthz3
QcQpIdL5OLQyJMEXd/t8rjViedjQGgHfuqOlIQa3bxxOvaeV0qPs7hsWxGDOUKjuv5LHhcDnzBQb
RG7n7sezmKOHukZauiqfWRx6LJo3BEvKQgjtpZM1D/GwXI8mYFjXLVUJ1k9rvkQqgnQFtXvSzkm3
29OgJlVOJNhND3x+zdWCuHO39cysCkvsHF28VsAPjmFSZfiPTt9ci9W9a4fv3/wxxXolzXs7Wc25
xskF4ID+0HvZ9eCxvFrWrEiuJOrb8gGnllDVHfxCfqnkRyMI3hFYmm6GSmcejQRnb3mTK+KYpSUC
aaJicHFnSduyO5j+aPVLQ36gRgcxMVUXaXdK0tYKT4LqnuI4oKMDc99v9jaUA9FmjGNh1riTa/3y
i+gxqfQXbf0gs4SZzKd7bO/qDS6812geh1QQvkJ8eKhuEvrVRuy3iIaCszA/a2f0SufrEutlD4DO
noLfqvkMg62Fr2qZYAlOzVn6QuVRQnuN/bXyxwEV8/kHltvdkqZqKSSBHkngOwrC5BddkXLJ9fq0
kAukj77yQ8gt+ruzH++Yfw6e6lmc503MQAEgVtPJ9+yeKzRWzXT8IM3vxRWEPZxX0h1kHVhvkYuH
P9N8HIGuzPUoom7RirFHfaT5pUQILSR93d4Z+P6D7Ayl4w421a3lU/DKol6Ct1DKeTqJOeF31Z6E
MIlgyDpc+0X6JQcan3KSLeTJCmejixPW69LPAKkL6F5Z73SAxeGENyErLeF7VA1BVQGDNVYAnKbC
wq9JK4X3GaROYI/qaeaq/czS3yzMl9yb9eLdY/an8D3fX0F+6dllTCJa8FE7jHZITujQhhSmu1u0
pl5GuThGxWZbL8ybDXoBLz///vSNQhFWsMT9Iv1UNbmaWR4V7YB5yqF2e1gEFDnEvZ03U1IMp4tg
6npee9fFi92IAZ+cw+rtueboOU3/sNqA2GTmYjnfgSgwFGMWGax2bB9EGj3TrUs74i2Sbmpn2QMA
g/L0KWNa2ge+6BQZ9EcYZnwYWD2MMkj+PuY2uf/BHv/8AUpmRq8utGiNUSKavWbtLcUieOGL1PMJ
ZWKcjBvLFnBPg0+kpcvNKlxssn8f6+Z9B59NMbAhv0GvHdFic6DW012ROBfYF2AIP4SpgOxn5Uwm
VFOKc08u1cgvnYZYk77K/BL9L7N16TwXzD8EtA5xxOKEYKQwAiV9uwR3p0s1LkmfMk+1HqqM36aw
kZFwyNwQBd//aK5J/zYV6iG9OlW/Nu3AB49x3XJDxhnHnhCYlNYncA5/1ZzrRUNioQ9lsZEcxxcJ
mAOVrjqaV2pk4uqGtMd8YgIhIS1H0G2KVNm13F7YITkMfh4cdhEwD4hR1uUAMebP5DHkvnjtf0Uw
pX7+VPoHMsRJ9fqJvrvIOgatnenS3YF5+gjWJwDAlg9GFpuE4pjVg9FjMvBW4fFTDe1DcupSobef
xDVTHGd8ryujEOZvZ2sbx1r2zLYcup3YtyPklDO20/JGn/iAZt/hMv930mO8qQMC3w3leldkzMQw
X752hvm+uykqz0/IC0qQOeAfOKQv2f63QvGEXR9ad9TVWm4PzuMLb3TE9y6INiuTh4+wCbwHk3HA
HpdF/jw9nGyvTGNxNEVyGLPaZH69eMq6dPoB2sImIscMUcoDDBwUKymN31BNewkF7LOV6cuKxaph
+D/qnbgG/ULQ8GcHkEbIH7f7EK2mweYqR/krANvRIMaVzs2sPXAS9Pnt/Ht6vEAZrhkR4U6fXEZ4
JFt5QwDX7v7+HcmQJCnwtMFYFVkDlQSxbuqfsFmvTElNc28IxxM83wwdEGyaFOeQySbadh8S6917
/Pp7HAh2f1N4V+30TtRkjFxGvDL/fZOxRqXZl3GgIu2EkoPN6XYAGGTHDNuM9TmM0sACi0vs2kJA
455ElOAw+eZJn/mNhPqHkwjI8CmQlbAnj7MuOGBFRkz/IR+cMsziNFadtSI4fbnqDeHCuRkXcwnO
5Un0fLZZEuyxWFpLSPbLnzTa1ZiG6dvmspyNQ49dDt5gDLyluY5OQefYmS8xYBUD0/0s97FDpTJa
O+rAh+Vr5vQ6xWjmBV0faUq3P+iQj0Bjoem+OpbQ2vCejZtVCjLj87x/VrmYnpJluYtOaePon7hW
Lqx6xPgtKjyPiLLPSxK0tNd1B2hvzUlBhOj0q9S+n/qTaZJZv5JLxuPo37qJ3eEIwu5gc8egQX9v
DoECJ+SEBw0sTzXx9cyng1yjBSJ7cvEDDbNV/likd8tvpn6GkGnYC1jgSsvUBFs3hfolAEfRL5Uc
MLf0e3NmbrjUwJIFa9vVDn4a1F0f/wn2fdMFeF3CBrk0QDQAI5gdgHLkwF/9jpMnYVXglXGbYCtY
RypfsMGUstk29nNMiYtED/zQ3pbwFV/2QPxhiuZcF+ToIOCI2saLXLR1WwJghi0L9Jh2atVf/pCc
In7U+Zqe4Iv7A7/6UUxuY1+/9SeaziUy1eu2BPSMpkGjgHox+ZsH3tgAiJXY07MrZgeTJJ5zjqV7
ZanKjcUag/YFnT+lyiOyISAcwvc2W24dv8/QN4tQQENO+eMCeSG9BDZUKHb82pLva8bO0NQUikQl
54r3rlUbmIKzp8T4+QzLMd87z/qsASZR+3+Vb6mJNUxBMXTgv9/nJRWYVE1L4LoG6+hv0IcDuP84
a4GeVF8FuUcPQzEQycAkYCTwawLsv+yD5ylxXPwVjY5o9VLyOD0Ub12/vlM4TKXFbDzm/cw6dDaU
5jwYyhGFKoW7GySwVzVLa2mleYd/UzIpQMcltr0HmeSVGFOmquxyOStRm2nZjvIx4TghSkmGdUMN
optgSYPLNQc3AEe9vQxxljVFTXeT7vrt57R/c8CceBcJzzGcjgpnaGyXRq1AErIVduWWzurs1HDA
HCDV01+lWjQq8NSXuQfXMuxmVvLVfcyRxeTPHMCMCM7fACbIJKIM2X34UU4JhEMFvemsJuqg+iqD
AEVBbZwuOggNuBBaTEHHOta/ABYFh9i1HB2hpCNAmkDO9Cic7igARdWhsJ8lPT5+TvRG+ctsdRCP
2VIUJ2KhkAn0zd+wQJYj9KKHkJ64pD3ipPquteL/N/UZt3u5jvVA9dJDFTo/xHNCVDL0phPxa1eX
ymwoK5nR+ljBTjEJ0/lheLTME1Tt5Jyzpg8+gmUQabPD0yomU+Etfc+lwlbHwjikIYSq0JL0qWRN
2aOsxngi/bOH2TCUFnplCBFJxWQ/pQpyBqs2VWOWYe4+Z+6uSBvt2Cjs7KGWZFTsPVDrMqN1WI24
o2qa+lSHUgVazyNiN39h9+5mmOTDg2IOUcxA8WioxSqJop3SAn0ZnVOnc3cFRy4uZdlTlJX/pv3P
pCvSWEdR4MJYp8yK3rNzxizPjprwxuUEnlRwbC0VGZWP9ovYDl/DOGNynzvFpPso5Gx+DmFTEwAA
XPKW0K7K/+7YnikwK85khmFR9BIt6Ehjn4OLhOAAUXqeA80qBZBsf5UVuuG7AUw4Oc7PGBfu1M2W
UNmTdST00ddoQjH3PgABFKxWOWkxs2mLUmqv/pFerP4zuoFbGr0y18rU2u5FyuPa0DRqEvATCTA/
uv3WPLm5qFCZZHeLlk/EC01ZqDIbhtF+5MlGxr9EiOnJfbmo2VjeL04EN5lrAjsruxlEtCnYnmvc
UibM3Fy7by4UkEo9TTVckG7DaU/y8ZKZiCwrZev4lf2zsfuFOgMc+udteVxitHqvpCeyNf5FZrmE
7d7r2BlOAtcvHZp9PllYhIV4wAQY/52KvVg93LheI3KMOFKc2LrmCNe0WKbrIfYS5j91M2gqZAqw
Cja2K9nEIDjduuLv9GpHMyySdqQfyGyxFyYlZL+zk2m/FXGO/iubeZ2W4vO1cxWKVv9Ts30sBk75
VXjqIIA5rZgyBpHH3Pn8yxgzJ4iRXZ7kOTDrCUoyGwiLQko/bf1MaKFlc5LhId4aWlN+eL3kRwg7
bBNndY0dU5sDtf+fe9K4idfP173wd4McbCZz27D6uzEATMmvT9ecJldcONL2McMdsUHh7899ka5f
KaDwBZwzeXp0RwmnFB26CMdHwwkpB9g8ZHCUezhOM2gLm5hO5sK59UFSgPvsLKLl17v4u7eVSdQc
/3NaO7XB5H4tymhxZzb+kXK+mAHqhsvbqhvKJAS4iAJQHzwbpIt/+zcfyeVHQG5rIu6WA06EGj6u
Mu8tOjW8gFnDAcrznXE6XJjPCByyQ9pmIRdfUsase7UM/bl63YbgZLjmfi3Y7xBVIAzUMVzYVrnt
+AL0QkhxIC1M3t4msjFTpBJt9zUTCpw3K+UqVien4L2UvT+TiiG/5BFqrh4rgHzqEleO9Dds7qCT
8iSskdv/S83T4NzxRTKv9QeeP87/s7nLKpqf7AbvJHWun26DBh9x395YRAPVpUMORDZwYdXpt6OP
iLmKIUO9iMJEtgdIFYD0Z+ew5Fqwq/r0XuTd5lbSEhl+JkgCzJBgrx5Rpq2LykEBCBavqCkKhkQ6
H1RtlIlXlPvexW7Rpwa6nOCCQuMAUN0pX4ZjSNsZ9q2vN1odho+P8P4h5bBBT1UVNsA41ySbTXXQ
uYiU07pyQhqMGoDLJREluvIYrxwZTY0uf6A3eSo13VHsO4RDukbPQL2Z47tzHDHMig/FG9M+vYDG
UqmgjlVbEyZa0VDTFtlU67IVospzChlCSe5e6CqhHv0z/Dv4UlaQQ/c8pxqPFTXXvQnh90zwuNFD
Ma+1sU2xg1Sk7qlnrHh3mWFbaW5onsTDEgPzk7g54rxiMyt8eoFgSEYTYQ10NhHHY0j5yVZ6UIxq
RitpgvCxfHHkKmsg0Z9DTMUegBJL9AVwJNhpW7CD9L6J4cmLusFMFKgb5KXT+SW4s+shlRniQl2W
lkWr4XkXwS0h4iRREjWXJh1ugUsmv2fgkTTxG3jyiQvVTQ3MzZ2qOzi/0gqCvQFNPsSgMc0ijPKJ
vDJGsVFJTGlVV+BjIXrosAUvmDTlYe1V1yMH2j7w6jVA7qPFz7CfWTtmhTCsxPFtNr//eqeI39we
pzlSjN8rwcBMRoYtfWUy3PIZrHGldFb39KBY/Yn093kaS0aIJQA1Hy0lMvIu7O6kjKuxVbbLLO8R
ZGIUMyaUeBt0ro9UICjgilsouJpblWJyyHBDkUxBxjxssFGpMNoEuDRPbkYj8EzbCSrAgYZqLxpW
4iqZzJ/UGurv9/T0Z8bn/V/G623lE4R+9uwj0rYszf5KnGvK9Zs5q7wMubToBYrqc3EtNVVwLXKW
/CRbKChaUYamhCuXsfkTrp3RHny7UjnF4HB7JiaxNt/QyAJ/uwjS7kWTKJFu7whVJfgv7c7wHPTJ
dazt5oyC8ON6pBiLK5UWUffOox7ry3A5YxauhbjVAjZiSY9cZ9D6XnvqYO0UMOnMoRFEjced1YxV
A5m4L5TQzKkgYZ4ApzSx4Zc9dt/m7lbTjAYrSSGKQuIUFxntn96Xuy1mcQQt9yjAW0PfL1RaeGch
2mwPMoXcT6cqOaXiJ4eexRF78pZXKkCaSEuJfCpDfr2eJqvbaDKMsJcblfb5zmowppmYplmnMtYz
Z83MD6VsgAIVByyfuRpEomTlAKZ1XsFu00nNayT5vEmbO7+fAg3feLYbY8inG8Dwhow9CbxiIiVm
Tb4ws3lEV4p7NNRUsUTJXJKSVGTTGnED8Yi7Ez5f5jbPOBYz+Z9/HbNUWSxsBBG9FUh+gLKnTKx8
19DKTSnsesGU04nHfIEYVd1C2MYJRv/67aMoiri4pvB4IH1rn+nmZhF52OCHLnAb8appRomxV1XQ
jLruiMCbIkSrMGcyhx3A66f04d/WgD8gkFIJLflbL3pTRUdLuRE0w5YTqlyZsv40rMRWjE0yJpBp
RiUwHIP2ZpJYy/Jz2RxEWk/T+eT4KfQNjgDmq5pf5oUHsgmIXRKIhJ9ePqm4C8AP92s7/GigNr3H
CM+mDlID2Y4bnbSA39/oGCWwhTesugEsLFb7GXsCFTHSufGXnP7G9GbcLZtKr6cuHoTTNsnoZ0cM
VUn5yvXlPQFpJUKjh5LdP8V36tRuBjuMrMge+mSFgqDlOHxebjvQFxPSm+6RMxwqGTxlbLF1wcIA
R3wLf5LewVTH2aMiFpSGg/6wl5z2HaUjA1Fa6/0il9R7/OiA84gL/bHI3YWH34OcTf0/Iwo+LvtG
qXjRoG3aJ11kTpq4OawMOqGc+md4dNsWgZWKDbqCx49uEybpoBJp1WLMZAwxvx96A40X9JYllLko
22AbOZUZdLdnAOEnajIKmhVAorEoNr/lM4QS6SIGg+TDq3mbd6PG3y/JzDYpmcsIiMdqKRdmwVFg
PVvSxorL+IkTP5Jd0FSdO++t4o6h0xVe3xyv6FtsEGkpl/PyqLPoVJ90gQu5u1R5lsYtI3ODk97H
N9uZbTtvn4FeMqnzcYvEsFo5oi5okR5AXiyFcKlw7cSvr+BJ6Q8niE8vmLJg4hYI1O97ha4Q+M3f
+TF6h02l/5uQFe+GqSkCmafqC42UEjZHyJtsz2my9wapeuYtm8gtkr/QXdyZ3J6B1T1B6fietdD3
nVDR4KVHs5h9bkuFW6PkNFM7ac9zJ02s6UtBPLK6ncDLoIv+GD+G/Y3BuydRCYEBp0zn7Oi+jRMV
nSFLtba0AmXvzpkuLxtHRYhvMIF85ZUFBTufNee3ANp5peM2NVuStQJ3DfYBFn9+OaoeU9+xfAg6
DjAoM4U44TqNacDVO4zhJhQvxHfKOIEESvNjQZdna2kU/Z2NXDMckAthjI+T7/oGDBTrM2CzK+R9
waCBwgvLv349xVuZZcItmZoneKL/OpOv4dqG6p/JF3smiLe6RVJC/gqs+9eUwacY5c7LREV5c6oh
If+CN7l2nvBaBXjeDKbQ1ZG0z1T1XmTViBXFHWr9rmqJKXkoWhQm72vZyyOvwZc4k3+Prhb5PjGV
WNtBSUhMhEOvOYUpnolm1f3wR3w8eb/fHojsmINKq5vy3XXNphHH8dWqpuKP0oD4Z25HCNO8M9jC
lT/8yhRwBUMw2m3i5Ifb+wRR4HB2oUkiEf1yFMfyuzxfrtMGItytuNnl0D+6FgKdkQcXkBgwR/Gj
HfTToUnIAo8PO9oj5esvCbuJgowbklcxOIW+rHp1g0qFa74fBQp73ANzNCYTvEIvYcy82NVQrSkH
sOih62rLelDh+Mk9nqp9BIettdcYeyqoC9lSgBhxSckIq066MyRuCN5vSNXsuljKphtovpZQ1224
bUdQhOx06bfJhRNNYc8O0LZJbR+OL+ijqgqlnvvFV3hyTmqZaYX3APRRYNCCJw2GJ3CcsMSXOf4z
fGLY4JDL/tu7A1loP7UZ1Yh7BQjSsEM8lBr4AMrrD7LH/95nblzoJxIfbgszU8BYMCHaiRNPgcl/
HxGMGcdUuX+B0vh2pYV/yvfiCm95PnJgRKXeN5wVzHiuo+Lop5LY00kSRXgvBzZHpC5jaMIoppcV
Our/nbg9dGE45D2T/rN+uFOly97xWDSE5sOySZZpx/TYcRYntE7H1z5P6kgi6J/Vf3MCiJq+ET03
Ghv+oMfvPQbYaGuakWJyAVwaawpv8+KCQJGwc+CIdQX3xkRF8EZvzYlvpSmx7nRGqF+JDJDllAwt
qcn64lgVrwSaRi0bjY9Fjg2m+teQtLnryqoa6B/K0n3iJH1w6/3Zd+Ic2+OIXPZsBhzZe8EPSHoP
E7g/6FTv7gRdSvt+rFdkuZrArmME9mclaoZs3oRTYm6d1x/ZHbwuksUwF/9elntfSOkBeGtZranu
MX8l3i+4LBwTa3xmXULlVglmtXHfrC0sVTTQxkJ+xLDwZ08vmDEcyrjfKYuH/wL7XW0vqYlku3NW
elAwvrWJXqbPIdAr1wGa7DLfhRap4KxUEZdQOygYGU555awEYOgKwv13l9t06mYZstzIqpQLDa90
hudY7g2iTUtEtrhvR2BMxF0EHz3ZZ0i9d8z0dg1ve8XgMzwO8GvyRfWZzSc5Jy3Xgfw89lyPkTbJ
Pi93j69/Trg+2uTvDa8JH6o1JQXbz1XbAoQhGWHJi+LQkh7HgXLqn9URCR39sG3vgEZePyXMXhsD
ucHjGzORyR3DxWzWhtxz5ipadqJvevXihPFqO6YrTm/AWIAMBnc2mCZqk23DoMapJ6hwCcjSOhOK
8GxIqMXTJEc8QR5TCRoU9qorMFEzclg8KfqhvLrPIkdRQjD8uPy7ba5iVqW7Co3RYqF/tvwsVMU5
v1Qc7svf5k2F935sVVOMS24jS/QGrr5j1sNpTf7qsugaWTe2VzYen4ami7BOUFZ4EAbbxBe3Eayg
abN1tRvhCjcqH960rrV6y6fq64aK2sk2RE0O/GTawNaJQnHzkWqig8ylPnRlroJ3LuuY2TKOfk9a
4xyKgwQt+qRZnl7+ju0S5mOj1yNHw7qbGArqdW9IXfJ6vhftPoEdyWUBrCuhEegeBtSiXCEOx8zw
hkg6nMGT4G6FrxRakE/8s52iIVLBG2aCacd6GSFIZt47cq+MFNiz27gjqZbwDtrC4d77L68kuYas
mJLWC+dVDoyogtNgyz5+F7+T/khEE+aXG+MGn/uHVbXb5zHuCtOujalGHmXmsmpgL0CTDInShv78
yglYdqYaWZL6tLiC5aZtFvm4tVAgAXrsjJpYZSPHSWChNy74TgPhwhax61cjDVH4RTABBhrqxYCb
MRMyBGxjSmeAndHUQ8tdvJ7AeBWXe8MSsBllwXATAkPTif+pjvJx4LRnAQm85EDGdtPKRJbj5IDU
8VKDZMONVCkVmnpEhbLLLAIrxxhUgKa5ljuVTAaY/8A8pY8xtZlC1m15NM0rTEu+odRHFnAMTczW
yehi1btFISMsqlwNdDg6g7TiriDNMchg90RYVsW9hCgAAMCyIk2y9E5w63OeFmF3l5iCKWrIjMUG
xJvBkEDKHNigaV+HbRZvnApTOELaukMr7+NOWELV8Unpuu4fJLoJgQpjn7KTWCEUwa3tjcmLQC35
5ttOm/3DZTB2yMwikgJPdxRPcGD7CPhnWjff9GJwV4l7IA6C/gewxq1QuUG73zAC6M1lkg3XCHc2
T4CoqAfPCOvIIpqvz/7266NYxa5epwEbn2EghPhp2QCo8iFLdxUDB/pPOS0lPMED17DXmfrisWiU
h+XXV9fL+FUFOkTuxj1Dhjb+XCenyIh2jzdRRywxNdxqXcNxrWccnO3L6V/TB99tlIurhW3Uvy2D
N8oFz4KsWNfjLm4dR1oSidDx9bcr4WC0JfSvv55r6SUzbw+3hYePMVg8VKpi7/TfT3d+HK4HBg+n
5NTFQG+4DkG+ygA/u0lcr1a6QIquOAiWjw/gRfGb+KbGJ/gbFKtMgEDczUh2iCK9MSm07zRXMfMz
kDDgWpQ8mVLyluL+M2HpBxlk+hJmR6FfzzAKQOrAoH5JK1wwHi4Wdz6aV6k591pcIFp2VYXTACdy
l/vXPk2RXE9BA25MsXczao9HJsJ7hWrBFVlSTldZDgbbjhzrImEQfOdOosJb1kjXjfdAGnJGuvt1
K5GMrJQ7O9zUQS/1mFRYdbbrZTx6dNOyWxF6SxUeGSfjM0rf472XTKnJvHM3kVpNFg6f8rwzomSR
lOLQ1PYbgf1JO8CJFdnLXU1w66WoDbhw1N61jUsXbd+06Af3d/WJa6zHjkwtsHklsdwHIdFjsqaD
Sh7LcusQtM036ck4rOJ/ew9jeWpJVOWmB7AhZUC0UG0Dq3Jvhqkq79seHHHkYT0tpfnUtnMJmUgT
/mZCDO1pLevw5aoQYqaIuQcmqWYkv07QtVDubJ45vTOB7s5TxciSB3IGi8zjW/OJKdzxt1+m95G5
j75wNd0r64CNry9zzWE4APtnx8FSlruCTh93Mlp2ghO3QfVBTQvddU709PEUsTTaUnE+in2OGAWj
+gnmtsMOJHgnFD1oYyAaX9hgbEXDREt3VWi8tbpLvqzSbXfCuHA6mOb0h6UbzpcyLAmgVRde4klr
wwM3bqyO6IoSjbeKkQB0kGMaj5HijSjQlLv0Xw0pwWKLFw+s0Njf3oEh6M/23JCnnNn3modhC8HP
+rA7sxqKE6JvZ7FfpqNEISZTaJt05pAK64lEyWhC+7CqzFcLnebhTQwsqSB1QmoBoVCK3j+vMVIb
YsYYXa/iVUTrObDGNHasGuTeqfQm3gB+QuWd9zhb4XrQFwc9nS0qrru+SeEGPWYa1JdtdYgyTxhE
2r92xb/o85bMOT+DzEFWEmVCzK0wRiRwPJkCx31+vI4OVXyXHfxdS0x6asg3mh6M7MLKnzFm/Ied
D5pte48DNJqQc5p4iW7OTRFy38Y8B7m3UaaRWRv4QBeQQunWm4gqjgk9cyg/zbRRI9Z2usPH54bV
0LNqb/IHugxzsmWsptfte+0teJcD9twG1CDphZ2r+oAt3RIUQsJp20L9yiYa1K1j1sPprtQXPdkg
N4Zir0YSKYyPL+XVgsOTraR8UyxVb7FouGqvBVQHoXeJurd2WEnahmUeaMOiH9mdCI2/MxMNw1Je
aFWA6sx6o50Oc0CjV570UPYqa7yAyiEiu8ND7IKekk0dxOjH/GjXCUIklErqC2Nt8Pkrj9zTt793
d+94OIxKlDQ8ZKP6FFNbckS+4aqc24eA1IyEDhgu2GN+CSvPCeaDva6aoQ32VvfG8+LMzyW0u+Ez
oFn3IpOO6CPVJJxXKJuMhWX3YvyFbTxWZpsuvm9lRVEpe+ha4ExhonbRj+Vb5NRXNtnA0F+5EnKN
Epi3s/ZivRwdiDhub6h7+NYyOZik8a0Xa5ScsSeZruojgxFGzzfGB/IhG+g7X3Canjn6GScbSAsL
+C1Mh+yOUcORNHQHLvG4Q+W6WJoLLEsFswQoMftQIzPQ9AsFMUwmD1h7m7A9uChB1hvfOAN/0AMw
cVIo5zqi7eBQWIRhWkYMN7n7kfvnsKkGXsndDyuPvC48qDeShUuqBsbgraEYuldDxrtI00Gc8HUB
cxFFLxOyScJ6K21ecM4m+HP7HQNjsaHlIqgDOguFPq8Zz4vZyMkqLpFqOh+lHE+H30PfcGz4FyqF
bypuQv3smQ9+HjRCC/wytd0dXPsFlaY7BxQCvUWWlQzytgysJa6f9HURjPHvUzutRv9l5o4TIZwd
JwHVkMEzTSTgceuMzw1tsvghfeF2Okw6Yae0MH52AvOkz09X0lNEJ/EijBHM/457cGehUOnHCjqO
pIPAUHr5WPGvMquY8mEraANDt6IC0tOmLt3+CrlSUn2kXvALU1kPlIF4YJP9OeYEB3HWZ+4epr33
dXNd6E2nQBDJXOw7SFAzRqqsRBaLMBULELz5qzPJyDCl14H+LtZNRraRTLC07+DvfHVUEEVKsviM
8eyc8ybdhYeORVrEjonra79V7iQLXZ7X2v7phQq4QKHIYTYbtSINLe4LlABfA2t20jE4+fCAoTfw
iWi5Bc2q19PfP5BPzSwuIxI9MiQ2quPlKGBLonjVHXhisR9MfgEO/xLLFyXN364Fk5nK1iNb09T0
nPq8Pnfya8ziLKaaLE3UklUlT7B5asMTFbhZxXVruBjqVIm5BNxOSVkaqCEdFp4Oy9zLdpp60Izl
//Ja82wAZfiM8R7DpMNayEo+GYMfVlk+qZF0dDcDHQljtvYEu9tzToE2ZYj9G2wK7Dhm4ChUzlpK
m3yzlkc8qUHVqcc4isyYfAk3/MSYEzkRaOpClE9Z4CkANa/YtMoixXzzgpLSgUVAukKCoAe2vclV
S9JG3AMKWpxX6RrxJSu9JKdNzb++p4FlJSfCsjb3eUnyPApU1U4wrATcJjye3aMEKy3qOJrp/wGK
596ZO6mL73VHD5pF9mg7OZpnqS6SMOn1LwuNwnkQKCIr8WgPxvRJYggwvTDLwuPy6Vn3hGHmVtJB
ftItsoREzwMjt57beqZLGBx82UbZ0YdM6V+kahXdnLK+9B6XLjNbQMLjSX9GCYRjJJ3xdxP1SbDG
e302QzbQNMqKJqojQ3MKP5w9BFv9W4pUPh/7n/Dzqrp/XVl3IZM07f/mJNTAcGUMJGLC4MQF5XEo
VEbpEdKvnZUq0Sm75IHlgXYKSrwsF0amOc6QazOH4D2uP2jt9HG+7O0Exv4vsXnoeulZjZpUL8kD
Qm+NtejKGC5av8gjDDVSzPttUrvhodzA/yVdSxLD49GwwKU1WiUMVwsCfspfdDM5uLdnfSRM4OHN
ERVKaKihJ6eMnvF6UXctfeUAyRe1KdmkvBgy6neKnFc7hMMhb/TGJD88VLmtwgCAJxrrHsDoYJm2
h7j/GDseDlbueW4lcZSKUDa4hO/VOuHThaE1liS5LPIj+0LENETBGMUK9wuC8CnpLOCNk+JGJyqg
B189C/0RJiqx+P1lQkjtssk8ERRyQt5UCDsQKuvboocW23tmSEyUnlRx0ZSX4vvyFKjsBkwrYZwj
TUlQmUq/HuyLSHYmxCyxSz7Cg8s+G7q9UUv4RBj6u7K/HxOuoZvJFNsEsNiYE4Hn3hi9JBNbLqxH
q7M/bDez/YoSm7tKCuPMBOCy+v9jh1oa2gVtQzRwQvusKt3yUWz2IRsUSbtFyHTUiuRl01jm41hD
Rv/LcLfawcI6uV28eT7K599eYU29qWsxsfa0TKkx81ySU0JXE1nQwiPP9hqO/kZBYA4gxbKdi879
6a0vj6d30z4FYoLH+v/xDCuJ1JTN17pHz0CCxGDH2LOZ2yQuFB7nvYJZm8W8E/QCqvZbtG/dGHwC
zvw4SD+xEiO+CMJ49IoBQudmvCuOXQxRy40+g+6JS+5plemyL5LmZWVo4tTapCaFz9+bc53BJAOz
Sb1KuO+YYd2ArCSD2hsLQoVJ6FzpqooRGI+C2Zk4zd5b/NmR+zOAirvxvKaR6n1NGHxQw392JZ0J
XtE52zCj0xeagtT49IYQ62plLqWZdTF1a2mtpS4Pyz7TayEE86Yynil2tMZG14mWfmIJpmU1DGgN
JBWi/rfO8uFAWAmDDuB1PtSPn4h9p4nNORCFzFbBGnLTgBETrbrFd/QigPyjvXvH/yLfUE08FFVH
yTTezIXDHsL42dr3rB48gSo27rUlnLqv5UretkgvbxVt8xey6J5rHvv6vPsLyM/nxl4h2yyYlgE2
XOmb+KQVO28e1FqOxVSwsBZZ456phYSdEFyI6oibTp7A3c1n+NO7h8XCbgMoxhkRNj4KqzR8OFVN
c9wo//u3pw4iNUTzOGLc4Qr2w5dkPOqWlVCsc6spX+0fO/roY9/y5hcGVPeBS0z5bXYVzb/Jyhcw
s3q6qVD0nx5s+LNT9I3sdqlntgWFsFqQ8GqnR42BW2WaIrjUPjgto/bruRr34Ys93Ry2OmnW1yHC
8WHJBLi9U26pqSn8X7de5rTkRR+4feBu2l1yGSNTXzKMuFZrGYDFAMnwv/QmBsynSdN3rKyEQy4H
fIPwviIVjTVmS3eY4XCZ1WfP17PkVtpjlTBqyxAXp+Ud94WBX1XojIHxM2/aOdOOyrLEbab2ckDX
FARIIIYyM6JqD+GSE1ZqiuYNHEP6pQNhotHcqx5j2TwbhCrrOKKalBJbdqWapbPFOCI4Mji56nsE
+jWpVMMazj6tjdP9AA7g9Ld+QVr4nRjMAFR3fB8H0gdjjDLuYJ3sFhZfOft8bCZ/gVd3zaW6bw58
yDuDCVDEAyAEDRWcaYfLm119tZEBpGuuOK2SsNgVxGqxm116SgWE2bXs/tO/UjrWEJkt89euw+bZ
HGE1CiC00GTx+Msp9BqlM1ThERkFw7YNgKGgx0XxcpJCQ30jkUo6yYGJAnmTE8s70Qsjw2FtAK7t
A36o57kIYB+773UAPuSfU0ByQezrelzlk9BI7dKohb5DMiFfFhceg7Wpzcs3VG5kq16JIXyhwHs8
izrSWsVxOJohs4y29ARSvVCyAXLcZ09hf2AKXdi9dBEWSF7Wfa8s+lzZF5asBt0fwEt1fTyVEe7l
k5CMjlg/qo9KztVz458CRVkT9qMVDI4Kx4xQDRHgt43EQCz084PLdH1/hpjCy7qmR9Dg8g7Wkjps
0ZBbwVpdT2XvSUbpD2CMGzMgyPgwDGnvQkBj3sHIj3VNsnQQRRZAXRhsSkEzOeGeeVDaiNfKMZsM
K7ThQxYywESEfyMdgFDHvMLs2pK4Da0vHL5rbV7euC1v0ShzIaJ91+KF+2yUPeVozlNcuamDACS7
CVKefU3F1fwQ/HveGhcLM1XxZiF7NB+3DdLdD+VqvexJ34hgRni7vdEmEMahHHs6wOz42fXDNFnd
pjBV4M9MHTdg+nzLiEGBzgq437a1+K9yo9CfwdGIu9XVklHvCU28Pcyiyrh6ynfITvt1zHwmFFA7
JO0dOWOydmP5YfRnaBMg9+w+azeKoMUtxrh9MHHtpFMt9r2j+usheKdWW6Exp3+X1WP6UaG8C8bm
bcTyy1hM4AtcS9HJlWnIFqwJtZKMC29okxeqpmzvdEfb2maS7LglBrLmXgYooWRYIZA3dbptdK/4
zhy9/O+F3Da/k1oMpKjMKuTtPMNmFoIuzDyckRg3Zh/j/PZ6DD3vI15/UTLuVcHZq90AjDsBgA7V
j7wYMsdtvofPCjlbbMcqPOmePI2UwivvJ7UgbVV+GlQjEa/2ZHKOV9ZL3YH4p0CRqWim8/sNng4F
LSJb6lSAICIF+Ijt6shho33UqUm2/XYd+uLy5nXaYLSyHtCwnEClFRWNB7RzQZSWL0nQhA3j0Wbk
Rr57klbm3v9CiD+JkXN27e1DZncnInzEM8rbv1srhOpXTd1gbUT2k5ayRV8bBDbGAczaVma17yDT
FaANXEFxFK/lUCGohE+S0cdfqf0epQpTvm6noPJVMcOv7KoiwZSwQONlQQ1rqfa36t8SFbVpX9fe
EjapS9L8OKukAbPxBF0y2qcCa+jtVy4aS1dI20b7/Npoaz3fA08XGp3wPs/eR6DooFjatuAh9L5w
rvWSo8vUy6SpErJPISgKxQ86mq+4QZeRcgZDD3Q7JV4xRjKvNV/CBfWszzfMc4AaQQRDVfk7NdI9
Xmj66z0NicKJljgVM7FFUAFGHmy7PlqYcoyEauIhvyBv8WvRItHZvaUbKCIkPSmoP4w1RIOFgGPz
JIG1u8dzdqvjO8P6s7AECgPFAA9JYxsizptM938qplBcPFv1yLuclBELDai2ACruawS/TvgOGlXh
IP++gJfwp/hr9k0lVvswrBTCeLco7dcD6PZ5tLwkmnAx5jPZiW1ZQIqdL5sUH3ql8gogbTeZCzHq
ICpf52bTokZEPDcEq6r1TWD53qFShPtSFzRI4BzKjWzmcGdouFYvdoVOSzydUK55dXdHZ5dgy33R
dPR7gzJ4fbsV8Q6ZaHeCwW2JRh0sRURi/x9GNGLRTCtiAjQzgtsE+Lcj9UcK9sEYTg4/ckH/0TvR
PtHMHq1tm+qFXsjemOSHlXkpkWZ3H18BM1uwX2X67eZxHNsoRcxxNfKJKw9UgvPuPaNjcMrrgfHQ
NpN2UqPdftsHrGwdmEaSN5SXGYJpzEq6z/kWrphM6Brd57zwrkJIhnetNHbtaijjMz/xHjLR0xrI
G6rccSZoirtds3pJ7dWkXD+H30IsHzR3JMSye71AHP9ZZxyLg6vkqsX6+uMFNfHVo62qpbYfAnwI
U3xcHlKrDf5fEkvlR8SUhoMxlUw/01aHCd5ZSl/OMUYM6ccwJc7n6IYA0I1c3knWU6IChgHu6Pce
pxh3hYJjrZ+FapsSFKfc7ikHTg06VWSbxOqzKkr4zCI8CWsY99BtvVGz4KwxKNlpsX3MeBFkD1tn
beL5ucAhwUTWrSGO2OOBZCVrSUa9i2VZN5dRU368MK1EbLn2XlXqOvVmaB2X95yBzvOp2w3hT+z5
OkEk2WyU9Ge5PDjyE/AhmlYq3rvcQSUCYMMzsBkFVr5NK+PSR6QVmJi4KTmueCDS+3pLYBp1vI/5
qwz2QT9OWZl+jmhL2pBmPi4AjkBGRkmkWm8f1k3ttJ88lckkcz5bcSp2RL/4rgU1gxk7Q4IfALPV
q0pBKkG7D9UsWoC1gJF722+B3P3/XIP0eoqtsPCTvCkqML3PYffUUt7kl246a07mAsFDMxwa1iwr
tSQd2tGfn93/6q5dHqdZ1+JxbDIVZFvXKgT5NDYdWDjxDSojonD4kiSJ3JpQ/nDkFZ9t5bKbf81j
rV16MTCggQuQFWBpI2/Q1sAn+OgS8QiWoJp8SmVswguVQpvmB3zuL+AGapKFdWGyhNg3A77ab42u
NxgnfBHsyH5rYVsygtwnY5m/OcJUuEcUME5Gh+MfGNGNHTvR0Ad/5eOJicVWSuzloPq3Xw0vAzcL
n9K73w6he+pGmAtUJtFR2vOiUQhh1sdf+pnBAakJrnKYrJGni+oKqK8nlD4dgY7kpvKcoKWpCorb
sFjnIIev6OWNTLGuDREJqFTpLxIWyEH5k1cW3AHFrEMFW2+FIb9PNprk9XQoZQMqHadjlMk6dPXq
D8lpQzgMa+Z9civBi9iy04zxT/uqnNIjkH4dqRobiiEor/hm+iRPbEy7nL3XcSePzMKS3ggNwy/s
81SVzbnFyZ96eX30TtpSi8YZ1iLCWphcIhN4NWqi5z77tdyDv2FTIHJcSz+DXVE1Y/Wpkm5KJ//5
dn7wq1QYvvYjxRIbbvsuy7tN4zjdgpRU8Xh5xiBebhLkiahDLh+6AEPgM6jW7N89tkoukJsUxg2R
rpAvA5dSql/bwJ2I4hQMOQFgMN+Xpn8tOXvDRCFJxtUqtRWahntnrrkQJpcYUrFxzmAbiY7NyNwB
Pv5+aXik9G0gbkpg4izivjKOUwNG9qfhC8ZdjA5yRb1r9RCJVR5Y2QX8pXgEmiW82TCQdXG6eEyD
zj/8R6bcWGDWWo0RImizsQ5iWm8w24RMJzvl9O4JfKRR8vhOqgyUhKRngkJifJmrIA9Wo+9fhQck
oF3NeDOuAnPCCzv/dOJ4+WD/w//Er/wNCGNy1g5/+fLJckeC1KnOH+9ftineBNGwVz00nGs48w5A
oKWwQpCL3GhewLRL1ZZEUADsf1QjZOrHJePuLNzx5BSZJkEL7rYBJhRFuEJQUJ8gdOUjfE9TdloW
ATTA5xF4gvCP48iixOfNtxGvv9OA/wpo3N2QO0fIR5NzHeRCcvc9wQBGp5WEsEXz/XnSi3UjxbFl
cyhlO9xDmWo9yj7pGPn+//6tbzD6ZyldnFICjZCpDyPV2jlpjpBdbdiqVypPgPw1AfOfzdJgn0eS
sPU63W/xDwKBg4aCi5EuiIiaamsvd3TUaI85gk6nGYZG/p+P+0tPGcYHftGf8imL10Qe9CHksfW6
S+1sctkjeGmjtxnT7lPKTrD7E+vF4mjriL3NSJ3LqRxkzU6yiE9SwgFZ5E7h5TLos+vHzxrOO++o
qwfuzt+Rz5Y+K6bq7C9IGEzY1qKItU56AXxFQ0Mt2RJlKuIRua/NK6GGVZVhtsG7tRcI3U+D4m5g
aShPw5HJ0h3SrEzqFQwRRmU1SILkknvuiT5zwKSfAi3tMttv8owo+ubkeiRc8NHFQPO87CFxNWIC
AjPhUUyPY6VX6DlXommLufc82m8YxunF23q+hfpF55urkhCjyt5fH72fyoVv3LM13tOo4/B2n5SZ
ios54iflu1MWc2A4sueIW7bLCOW5wIie57KOCIwQdIBx5qaPWKIY8Wu6Hml3m5ZkMD10kre1AZiT
IpNeIlBsahBJ7E0n2rZiaoPD8kxG4Dw4A69PteLd6++XzrawBU6FwHmwRbN2lscIgp8eIAY02BeT
2dkuAyQXlB7yS4AS0XUr0p2MOczdifJau+EeWgTY8aJvNNbNvWwV/Z82sECa1jMhJVyomqMEpSXH
1T3Clm6ZXUf7giwsANoV7dkqDZZEEi9V8kdY9UO82ljFawxv85nTFQZfXLTbK/+CPvTy6u9KwWZM
FDfloBvWe3iNb4BEVJLEkTI4TVjmXV+VYd3fooBJ/OgRDZRswgo4q3J3+hmzFtxzKLywJ4bbczLh
9isfV/t/DoEEWPu4YBfpgamIEcqJ8I5aD9fApU8gyxu7d2rRlyu1s9DdTjDTRehFs4jYO4t0gRnI
/R66P4ac5V0QpeCApr271vQ5YHnyPiO8RVLREEJGDndClI4FVnW0rUIwMVXxUSerzzdMTJojQ0R+
TxdJeSmmmBOh34HaouqndroqaVl0vIEJ8im09O+gJGFpF4ZMoBma2iRqdQn1Rn8zQEaTamq1zH5F
Lh0WsKSN/XvoEdrbC+7vVexsDHc9yeN2hSbxXOFOhuOAjRP4ViUJ7Q+riWhtpxGakQt5sA6oC9zq
zahwAAqrMA1PdFriOPHaORQN32duQ8GcN+c20pDhCRFsdBTVLa89WazsK7+71AcgS+pMRnZ33m+1
wWrjxPau3ns7GgcbHfsOMJe4BVkl4Dbo45RvOJWWKgZfPGQgxaRDo+3/ln0+M8LP7IgEZKWh0Yck
Qk8HJCRVhLY6qXM9KSux67WiJG2d0O4KfSxWCFwwBBJLGFXmr+rcqgYO+wwZ5cTWHUJ44l0jEWxx
na/faBI5965IFRTRaOTK4c+4OvBPjycVc1AGmenJt2L9OrTa23q9dmbjgRBXa4MtYm/rot07XJZN
6MhTgarJzLH6pO20B/KiClfVhf56ITdfNr+c4K1q28QfFHwlz17mNPQuwB2tUVegNG6nCetDo8vk
PfyiWiaCtyiBe9v2YKlVralZw3PSfCIKwBDNxCI8h0DegkSLmHQQC/QINSLdsOI8Cp63Hg1Jv2e2
yco02suwm/tm7DZaAsgwDUmGnj7wtod7/w8fR3tb84qXwbdUumjuTpXx1KOZkLd6z8rj1lfBdBsx
Qf7TPExDoUSz0BUwLIbQUksQg7kIA+gl0d5C77s6PQLEMg0bc2ubMKMi4aq8bS2CMAtN0krnDZPq
34C6+74lWYT7GzTmHszxjLn7srLOIVlhhbXUE/RUcWeS5mGn/7JSEx9UX6hXtjpj0ArD3hrIm1KN
R4MGyXgBsh6xNcc2K2kbOGFT/i4zarJRWZYGB+fh2JsSarqTrskDtA6KmpVCJq8Wj8raFuYUyLiV
9ylyzOIiUiXXtTPAQOWoA5FPqQf/MhXebiwwwAJb+AeyK5p5Vjxkzvi1B3qOjGEvlKW3I8CPOvf/
T2zyiQKDtcMEQ3xcBtyuwn994gbjuuNXZDpRqWSE2JqSYWzsm+ST8vjb+T4xFJBSHpGIMa3TNUro
VvYvlHxD6xPyZYSRVDdyTPf1nxlSl0s3nfpUy+RI3AqxEsXZUYQNgiTk0bZCHvsGQ9qLl5IBeJ80
8BARBi3jPYQ22jY994bXFmyPZKCDdwzIqgUNTn8Ap9oeqMORI3yUzZweQW+ZA4XCZJw0KIkwhdw7
txKuih/jSIjvRb5MPC7iLtnisDnfZR05H2vOdB9LDqx3McmD11C/5aJ0Q67IfOjHO02Lqt6KzpyI
l4nrjEfO3pSRdsfRK4EyIIhzwBaGgmmFdJud4hxzzqaZxrjx5hcGI9auQrRxghV/R9SrFHEm/JFX
g0epKC2ghhDDrWV0PNxJuv7G5xOeGmuRH+40DSii72xpnUjCAl0ig8rwHdH4fUSJWlYjy/tIE1ck
Ba+ST6Tv5b7LkjwleDxGbsDxS44fFa0OPiHZ/V7IfKkryFnccrD1QWkwUA+lUV83xmoUf9yvngBC
Jirr/BvZ3RwPNifiSYo37XXD1k/kAlme2j+svgrET8hWu3Y6dZODHXPhOhpKIZzWhDfIsNm4+W7s
mEaIX1FyTFyhmaYPxWEaXIpO8MqzP2e/hfLk3ethTuj3iIyYmDWDzVabdIwvexP3yNr835lF9CEz
rzb0wIZ1eDY2/XFKz22sGxiGD06K1COGKd1avHThsbdZTYX4HnkgN2DUK65YoKim/WNYKgKeqKw7
qFhjogCY+u6ZF0nRW+L9OocHxwEHO7cfXTy+nBjMFRSuYGQHYXUISl07hZw1P3WHChocIXO0DoZd
roQSC8zj7rhkvpCjWA3dLQPoCpkAijkQFz8kg5mdtm9xy8I0RwfgEqdIdCkNiRsJRCjQAnIhWMiP
CSxYoqsYXPTRncVVwOBhWkrJj+2r8ryrV50rU3pOhApa437WSBBB9gtqVQ2THaij4uD16KIizfl6
FIgNH2VMxbEPAWexvGK45AQHGEOi1pO6BwjNbopYrfuZ3wJvUKXr48Bc7UX7Z8gfIhus0b3ZRIhI
2M9aT5/w2drrWt7CmeLZ2CTzV7tDzUOU8w/BVcbm8QRguT5Z+XLyymRfp/SGMbh09tYpW6fZFaen
C2oQq5gC0c8G5QfKV8xK8PC2tKq8mIQ6nVthW5tXCpVMl3VX+PdnZxHRQooVltqoUhGXwHejkmp6
8KJWmumVY3zC17ExfmFwEDPBdN7iJ0BHfDa9Ho2lpMz9g0HqOZbnvB9s2qkzofOFL4aoQEmY/ARK
7S1DoeILiItT53D+86xG7MR4YzKSTISfIeWu0dyLMpagegp5vZpOPDVLRR99/eBozH9bHMtZZOAT
9qilmq1gMYIBPEd1G9k/ixzCoczdizcZsJc5b/F0z75ABe0e3C6pjWc8qFMSo3KWK4W9T979+8rJ
M3CkiagjOpgq5DObgK2fzkPVWWiLX4qoESl8Hmxc808icfjOCj50X/Rbs1vPi410tQ33bvzFEcb+
zF672NmS8q/WKIc49XY91k2NzFFO3K+MDRDz96RrSr/gRU8FKRDKwWJZJNq7T0CGzOzfBbEBuP7R
IEa91ZUcqxcHTJahS8P4eMGEVC/d0RzC0ddgd30S5yXu5DyWx+Tx76ADVvKuXJxWsid8x3kNSSh5
LtBVmtuc127kq1suDerIUJS+b8iwHc4Nub92p4Tr+/NJD9IKbgF88C8woCLII+5LfUDnEUWr8R66
KQIikdzl/DWlYD9cyFmSo9W906J8x6xq105kGb45nZ/JJjB8nCKfyy1l6zYsAMezXht2r75FbrDg
s7aNX/PlrgaD15Ke5GngEqv9VI2/L32vKNzFp8pZH4oZMaDRHXQxSu1hgaahl+dxGtSqw2poMX4g
qhdRIILZpCCXl4LhxR+n/3FBpuLL5HwbPVlSsIO/DJjZkDuO38aoyaDaaEIVXPOc9eYAG8E+IJ70
df01nHP0P45uVjWx7H5zlXnY0CwV9xHK6qSsjx+t7GuMoAHjZwNQJaRNdZjoS1WeBSp9B3dI4kH1
cetbsYiCxuiGzq4Bre03+a8HkW66gbE+BxSIKjCN4ptjg1Gn14LiSmgH3D9wyFvFWuxVNIcXVTe5
u7jEjk7O0TXqypn1GBqAHLlE4ch/lLuR7uVnW1EZtjYbs25nL6j+3zjaVnUsXF958CEc9viz0q0g
FtCyGqeNu20cKljB8+WmmQIz05+qyoEDPcUu1DZlDsPABLFS1lgXZLPj0LoVJ3CfEsnI05cQNI6V
t/yc/wu028n0OTN/LoUa1fhbUGuVefCu0yGlabyR7sVvn1NIS9ZXr+MH4s6GrydBhL80EKSWtJs2
8Si77K4nb0A2rXeUIm30vZsbljuEwBaWfAU15v+gYql3klcP8OK4A9MMUOi6nT5ZMCBWo2j+9Y31
kZWqVI5T80FBFdX+AFgr2VIW/DajgfR1Sqxllp0DXZBFvN6QguSHJIgKelsgteIe6Agdzo4JrGvo
5d0GZ2AEFrlPafQuuoF477JM6WSvKJjXk6mG2aHIgsmw1I06m3OToEHi8IfnEvrckUFmpUNFdDAv
pW+U1uNBCkEG8CuLtjtgOhBFBrLk4VNNDvTnxdP8G0QtykjW06PeSFZiDLf5wsuhkQGbbZSSgH4F
oBVjNUHTMn9esnBShZkd3/lchwqJu5aJ3BpwWbVd2LK8z2K4gL8aFfSm3tZ3qkPMjT/dNNzMbRHK
02iuzp19y0xYkUbMC3rhtvYjKZHjtKiP+TeTkGVOZDOVLUaiPDEh/mfcAklvvh/21qPMnFUPRbGQ
5hJzGYRQWksCU3tkEMOQ5jL4gfaOIkOdbuc0GVFCPKBEPHKQxBdB4cWs9EzsDlnVq9LZ5IYrDfSF
w8MKKHAebTFLSltxMDEFB+N3YyTf7XXu4wUCSJfVOTaTvnPMBmYvBba+2Gj7kJuaEKjFRtNUs1HE
6VPz9UuKK5Bka41dPwRmfIY3rH5Lcacp4U7SdCy7IKo0K5qgDNr3z3deG2y82V3cDSxv3+7x/W5l
gdadak9l5E6ae6KH+Uboyd3tA7N6TKk7TK/Rw3YU9F5ANNA1LoZswyXkkQ5YirbBd2mWFxcJqOH7
O8p784Sag1y3aE5s8oGVhNlTGWPOOPoaqR7KVtXZ7/G865eXhxe0qk96vr5muOv84ekcfIZeHMKj
83Hc+msP0auV14sZ6IA3SyZrQRn4UnOB9GPKuivtfQdZuViCKzLM3z4KpqN+38WU3C1FInVKvQm4
pTeh28Uszhr95F0sTEBxPVLOhhxnVbwS6CWyX48by+S5Mef/uqkac90+k1o83ePtLusLjMyshOwm
g5HOdKA7dP2RfSbNdRMuXT/zM6Jzq34XCFwRzU9yvYmmNrxWfwbM4k2zJwBvy8h+TBGzayb+zyur
Ec4wAmWhVnf5mWNiyi+JMesMdOQFBXdFyFBRKF+X04sIiVgXTdqELa83EiXZ85EIjK7wYjCrpexa
eZ9w9i/qPA3tusRJdOOj+zMg+HhzZd2UONvtCD2CMxC669++q02H3vt5QqD7MYD+CXv5dCeBKpeZ
2q7tJcSWihdm1WIa/fmQOkfaOq/x2x7qn6FGvI7sMoH2YdTCGgFIyhbOUH30ga9Hf/V74tjTnwEc
MtwwT7c5TfX5wgPDohucXqkqbzxqxlyYrmGPcqe97xvZV9oLLXE1XMJ6ZRHyBP5ELBYeVB2Z/XTk
GJ+2dXv7GpW3GqewdxGER9K/8yQt27xLzh17VKvGk0Q1zXLjA/9q5kV2bYZeUaWf4LwQTDR5EVRj
Td8+LJkdyYy2ex0uL8EivZvXp0WnPV38LpAY4JrGapCpzgXbns2MUwiTo4pquEZ8DxbqJ1Y0YvW3
FVykKg3jYshmQdibsg/bUc6rk0I1Pui6jmryoQPWcYHWYo8xgZFwOoyh6XPpbCgnXCJbpf0BN0mP
srEU1T1VpKlbG5ROBZgreADYrCeEsKH5w1inClSJISJamUjr19lrj+n62IjCv59RzEJA84/WlW0H
FOuAdffPDFJhdeBmNzjQQIAc5mmXS9D7wMjOEI1Fex1yejV1GttyIZVJ2h+RtfhnqyPykyB6bjGn
hFMTXVZGcxtA/WgTHzY7YK4s4M0phPV3K1dRA6rB8+3sy4c2ff672D6DIMYpakuGz0duyGIF6b3I
WnniOO8DQHupDbXsFeCahKhqMfYMqQVqpub8U+nhVMtGaCUqRR9R7Ov17debku/7vNOVnG35S5XI
3O5KtjN4RrwMBr5Q+5ZN16V5EQj4ty+tZKz4q4muxG+qvscg9uHg/VzQbFxUGcgoxVvBr1gwkYhv
pZyFnLrBz2tEueCiNzDFfiBNwp8cLLftO1PcCRRKTm2raW+56i66bMaqYYhYXIFuUjNszVR/XmIA
qA4bM0FjLDW/qmw/zGWjB4t21vUA0kcX46Tbs/Q1mxdHcv5GolAhnmlOvLMQf6rBbzI5sCebICVY
tmiV7jKYiLCo3jGiiIB3K9FI965yGkWeqMjp+mKrEgG2e0jMUntpHUXHIXYfkhW5ZzKKo2SvzwBm
XBzlZtsctbboFsBR56L0D8NUG1zPe5tnzrAfA6q573rhPA3NGdb+C2QxjTzScMO49JhGXVSI5ggR
5BqllVs0TJl2JQbb28/xkIKJVxmPJOCLQDCsznSqaBuCQtkE+dJx97Dni9foj0FczupmA0ewk6Fq
PPCsqzdBUWELP2PQZ7K8JFjnlw7msJB4HcbxTFE0D5mtnPZ/vRBjMYw7h2zMAcI3IAY8fGgPmWDI
wU2LA5sxBGsCtIXFa0akKOZTeSFXRFf2Y6clpuCoGNLNrMSNITP5M5yKtNLCcLqX4FiPBDDcrIt+
wPioWrPxQ49NxKLVHCn9XqKAP3kG/TaySD+AkOcNKp3KEdRC0Pm9NtpJyx1lC4KNqyLbIGPTcTJR
fAgnfl9sUOtzaKzUUPees1cnxshu0T1YUJQdeOlve6QDOryJ6CgoJc1DxjL33RuVYXpI5LqWJ213
K9LSKgPzDWyRHXyJsDkz1SwOOvw546rp30++fZN0yp7tj0Bgnz1IJFhMNCoZ+xdT7HKxJWp15WWf
EDTatNwIMVlQfT030anHgNbaZLESHBtgUr+HaiEhpc0w+S+9kM2PO+S7Tg9woP6eBdbdAhjt5rmW
ozECucDQygeaNqS9eKyjrMSw4ZNGRtLit8wRrZAaHhhRwtBoHRdLtRSEJtL7XmPsV4WIaRur5C+y
NnmJ8cEl5AwDgLHBkjR1zQOUV1q+vLCM0KePYB3mVx9VEE/C/kQbA+FsC8538fVqRarH/pSzLYuY
0QqFiKT/x0AM/PXiodtGzAvu9JvF7JwymKIgUpIITiGJESR+nEcDTvZQWrPFjQB1F9MSQPH2JElV
Jx3cxyckjd41n8EOVsD7qPWu34dIq63PF4jEqfxahhXmblPY8s9zjYow2H+E/DKdjDIJ+pUt0pDC
fbUkaWe689dOLhx0KQRV/qzZ/PbPu189VgZkcwt5ap3oaXAMI0z1gofWqT4In3zv+SLG2k1cLWJm
tFy5aju4faKYj/P4xnBcfIAUN1kiZoBVTDj7Ssn+r7hi0rsjOEveWu7oU+lgRvtQJDcxLiuaQ4XU
mSgI3tsc90+C6GPFbpqQteFEWPiIYdGfSw0lRa0elKmD0ArZnIcFdrM7GkomyxGGQvW8s72w3BLK
NmgdZECRVkDmCz5eehqv6zEv/p8itVtt7LbV+2ROw1/BJoaIMsSDfJIbOjP1DYIGRfmp1VN8oMqP
nKQU8Z8km04ZCzCDYfTN75kpu463KRymEoxbf/2Z8bHQTd9nHg8s1bUGSfDBpS3W4qX9c3g/H1Pd
bXSAUKqe4IjZ0P0Vtcu0QzIOjadTsaR6vkGj6WviBX6v0ucp04lVkVbXXpIUfM4Oj5UK9yovZN8X
w7ok0z8RR/UtjML+wQkXudQ0EWXZ3ZCrTdWKPe+XMJeYI617HRdJOR/oOQc20W3iFjLYyjih5Km0
Uc8aWsJPgQj2/fiWmtLGJHr7AgaUAdkgqEvWo3FRquEbFc/Pqj//NG8GrG3rAwh1+qG8iJlEf811
N7bo1B9Dt1dvDIn18ti92VBu6Fx85pRYNPoQSlJkwjTJRgEpOpnMRDsr1ZTpDJna54RNZa6EIrtX
/ow/POaFt037mjObhiyW9Q3slc+zQWwPTCWJRzMC5+TOLoQ6j3WepN4n6EtES1sG1UHhYJ+pq51/
stekHFg40gA6bh+8mmDO/kQ7nQ5JLvPEw5BEha3u1rqZ+fldHltSb1m+jzMy8GJxQyf8+q27SV33
nvlOIhL9rGXUsh2vj4N+eWkZM7fu+YlJFv0ie6LWKvzr6hyTrTn3xShlxxVG3nj9bT3zHKUckKea
iRsaREG6wqXw4xCjqgkFV4FQLPWUxTkqFl+jjHUNPazu8hPuZEDw1TrcJhZEh/nISha2ltvxboyO
tppEmRpjljqj/vfJfqX3L5AHYppWGRFAEOHlagH7SAOW/okcGt9kkEngzhDRIVJazfVyvcuU3Xwo
mtIQa3RMKpWmsLRDGvRHABCkAOMsLRvvadYS7jsvl/k5U2/7XQlLabWWtLUOCkI7lSJ7eFeNxrnx
g+/gmaOEb5qgYktk9j7b0oOUPJdqy5cEzd9U/v1RT9z3LN7151yPDVRKpCz1rKJyjqGbGsLgKZMZ
wnRGa4wuxWjcYhuck3vW6KkW6KuW37ojwaafBs6hL4hUm30cHplou4aZKapRJz71BoPPB+LbDYs+
/dD+UACLzDPXjw75xPvXkKJjBUP8qYdcC0FP2hIiWmzO9x0IBEZ85B+zSTPuYrGsJgfXk3mNWk7s
YmZa2y4Xw0VmrpUtxwEqgJ5j48AeIYwT+kjh9u6bMzZsnMrQb5GPWh/TatZG0qDYtzBxUIDLJpt3
XeoJ2KNv9CIeB/J4qNwUZkSPiGAeZegYUi3nRq4q3hzb9aHGZWE2NG0p9zCFiuCyALJ54lDTfv9F
ooorwatDYLtTd++i/hZtdkS5RATI3198EI4eA69jIJfFkOuFQ9z6Z3WKA5r9RQ1cAXDSpDszEvz0
Gw8uNK8+CvPxrtMYje7PrmjC/EZGhxQmZqyEbkCxf7ykiuqHQ0OjqbNF6sODFCe7CqLAgmsjlr4/
iNKfkBje3vgRBap5EkjODIQ43lLW2w2dBhmcRWdKkEuE/yAw75N2iaeL+DHidvjqXE4H2MzAFaSV
+NVJq927X7fHgJM+h696/r5gMj4ItoUEADQ4xAFnEGIvvzRlVSNFWmS5RjqGLQ9Jbx7NeayDMGdJ
EFfGfCaeUcfLpSOvmY/4Re0oOd3OcF1lCtb3VLEuF1HHsdMVvuqOi/AA925sB9kfDfUaT80qeGNq
oaPe64HwWp2qze+jiA6UoRPs2H/A0eKy7YKZHr7sr1WQnemPpmjgywfc8oafvviD+o6upHYsuLf/
zdgasfVgwx2vYxvxD7PSG3f4f2LgRziqedIiRJSFF7xrkp+GKBiGNZ/4dcFso7iXs47p8+93Q1Ez
pmoSp/uBzGXUHTLaCdzINU8UzZxbM6OQdlU0foNC3l1EoG7vPiWW7jWwHkR8kQITqYw9g1tCB38z
v9ugMy1KH7PBxadtPciFAqlPFtY0pDIQbWaQ3KVA8c3EtqQEdqKyPQc6BTiQ8aPVTiwsd3V9LVXb
Cn4Xgaap9JJ7oCDrJPQlVCGzjbZbU3X39+Sx227dWKd0Nw6a0ucnF/tVknhvBRNmnDKhGHrn5b96
z+GkhrirqMylsQnU89lYJbJKfUSldabe5DP0RekKygNEdcPkZxMTrXOFsu/2Xbs8a7zf5DRPUnx9
guIQQhEPAD6/2FQqUXrqEiNS1awdtJ+Jh+vrESEtoOslZS6SI+DgvGgKy18AaEu1kmuyJPR5e3M3
TAQcr3iZpFlZ5y/T2qWl9gVid6/EPT5TSJvKqdnq6vQWqTSb0fsj+zdRJiAXspg5C9du6GmZ9Z7/
EmjaWryP5KtCnDW1KSNn/KhDj8LYznKbBVrRQaGVKX9fgzB77ptPxLP5HoCoA9q+poHXvUL762tt
dJS9fqujTPuFi/Yyb9yDjW4Vi2B4O4BHDdxQLWZuo5tcQVMO5p3oBH5usukUsN+HzwKMD97EJxnD
rq+TcgZb113+WxG67I1FVL1e68DxOSdg881tsVUaDwy6HNzneqYZdi6cQEmQAjXvJ06i08VV9FpC
yb3m2ThyvfWFVH+dS2NbXb6oOvwVjZWock4x65pH/k2+oSZ0DvLgQmSYE8oxkRksgM1h/o4z+L1k
sN6f4TXujdXwdaElapTBZGtkxj2PywhDOexfhV2toGJAv2fpemsHu4iS1MkSwja3M7jva+TDZIwS
85drgcoNV14CZoK/UYpyn9PeXo1WMpm5NilDKCFxycEmxGXywRjsI/8m4k5/+pz89OrTDORBjAe9
CGI1+HHXMyHenclcI40z4CMndK1+3RRMiGFOznttCrGd2tQQWmgO4hX7riWSrnDAOPJIDMl4wxhj
QJjqqxQ7gXHAGB6N49g/lnVUvqwzf1mScJnfnT8x5COQUmGCzZLsTSbUcmFafX0ZYjAbZjqH5DK+
16mjkSmuOvHgiW0P1E6HSXFIuA5gql96LHoUX7uEWeC1Le340DEHqRwRKhN0iNfPyITVorBugrCo
03tGOCeZJwIG7MAGMeHp7ABw83NVMTZN4IK3XMCcr3wzNuIkbVuHgneqInPwIB1HE4b2Dnn4Bo1I
u3AaFErAFR3tqpYTtGcLrNlI55yqvNKIL+H2VM8E9I8PqWpMzx+3uAmTvTQGwrXpN/pewN+v2ioA
pqV2JiuHzeAsuJ44gg9shjHGpg2CDZBmllDQc70zXbb98tF0jk6GIPwsnftDxf9N09RtIN9R2U3d
N6mLbBi9uO3H+AYcAhCAIjAw2dcMZkGBGSBcmIeovxzpRCQlLUSUYoXwmHEgPbOiTAqhyPOWDrWG
kTMTbGUcmMUXLSaxnrNe679cD5tLFMg4A4KTovU+oYhgl++JsKIXiSUY4yvz+gSlYors2bzgPeCT
3mlqYMHOTV1seKKIJA3HKCpobpNnjliVKH6Ofxps24pVDWN2t6tnhoTORrSS08CgTJ6vhzCb/EKk
3Sa7peD5FO81yXD8SLkoNBIQJtVyNMDwl5brcMKWuMTKlOtBVt7u/bfx7Ui+3KOWqtx1MPzuV+oC
09WoqFKDLCO96vbbI01zi0xwgcNNc7sP6dJ1moXGn17QEMrmm1oXrHHZNCXPALkQXpUND9lZaKsS
OElAZuBvFqvGxeGIMxotGGtDL5hd9yEIOeW3YBWmBW0c/jWhCqiOCi6cO1sqtVxDimosIrF8lNVl
kVF45+zW4QCNlYw8G4tougj1C8wX8R7FAxHsn5SY3t2WyHSX4t9PxAt8YaCM6EXNWjgv9OpYnT4Z
ONO1Wu0XVOQrYG4foIJiCejksopfC5+9KQGhtrAB89S6SYy0Gs8KLnRrn967KNB6ryLvwZDJTPyZ
6sQTGaF3qp/9Te8HabQVGzd/TjMXCOCDW24wRNr+6wqcX16XR7c4dcybNpCS22TyQ5KCFxl57DLD
WFjdYWYL0LWnUoDYhPjbQyeZrBhZn5DdaSIMnkRPiWwcho/+9szj5dCX0/GKQDi6BAyg6sf7DIOM
z4nyQW2ShYubleUfZBtpAk5ad/cZ7JXCoRhLkmpDYOZFZ+DwinDNDoxfZM+oM0Tzz7x0nTScCWi9
Pzn3LsY6M2QN7NffywHNpFRsDyARxwpRmpBKkCuSjU04E4QAWXBLtM/J1wXKDqU5ozZLhFBcMxG/
QcNfDltZoIZ8pUKvNEvD/HqoEtSYSZsHrOGBmNU0rtgxT/hjq3fD//IFJ+gr/zBYqwWTu6R0OXpt
ZsctyuLLGa7iVNY31hroKdXPECWB6kgMpjnab9HUDQ9GknLwhPrAAK9j9MlStEiawluPuWoeGYV/
xULHRsw9bJGnjgugDVY+j9HVhGshFPgUQyxBOtlUHl15G7g/ESbG9M990F5QYIN667AsJVKHufFO
nI2RFtX14hJNbI3afGVgpLsQ7gB6yuozLIAohPkXX87w2VO6oUzkXJtfVfhisB5dSzpZx72j1sth
nb+rYhQY06phRICy3q9Ae0QSYj/VI+J58ZzGn35NhKREzyK24Or//iT+qAFKMDzkbh9c2UsytHwC
K+mBCU1V3ypjD4t7+jctavrdPJk1piwatlbrDtJ/iGe9yLUr9RyQAivI9ewRfEEHTDyaM6vqRCiS
+kOh8RUzoXio0Jo3/rdIZ8tEGq5IpHPVFVSlhTLMWFsbTa/any6AnUmZgEG8g9wAt+3hYlVXS+Dc
8CFE2pcnT3DyQ0bZ3p13U1hMD5p8MyMk5goGix1nUv+j/cbJQ9+06RRFd0VYlMw2wTq6vzDA0C+7
nW1B/OsOIRynPAfSww9H/k4DZn2LF8+2zXtHK2DuZC9YLKiaVrQ+pCI2u/P3840OryckXDdoXQAG
hL4oWXbOv5uskzxzwq+uUCStH8mE1/lOFnIaOV9RlDsY8g6h/iHmGWz2oURe+UvauP+6izNAbdco
pVsA9Cze8Yw90/N5hEX9d5/W1PVy3Jn3qzy2R3aPU3tL4Lp2dihxQatbKBU99RjWHA12vS7Gsw0z
XxYcRiSxTCv4zfUehIFSGXIj+EiKxe75jYyIeVZe5dvlj476t1hf0ufugGy2+IePTsouGuTndWuq
hjUf0nrQvimY1NxuED2SLjZx0BGrla7JR258qYNmw3TCguQzVODH4jDX+UckpqoRq0pL75teoizW
PxSemeifq9BBPUbA3weUgYwO+iXZgLzoAo/PRG4urYdODSQ07/7NJSNGTHOnPNPyuPdw3Dulv/Ub
hProCwzXCiyoYoKCoqv3bninvbw9RyPsuBE31AYd7B13SHGyRi7GGhVAkBsEjEeHvZ97NdXBgR9U
nKr60JQDiYIhRHnvly5pt37olAba1bOYHmOvfEP7PIJTPFmOSNZK3CF/AEyfyOI5D1IKd7eryHPm
TZpZWl8q7S1yjOv1jYkvPN/DVR5u1JWNg28UvwGyAkm2d5mRQ+xuhCkBmfDCj6I/2r+RahbhLCqT
ZiomMOk0qoL9V9WB0otaTpRO7icPETuvNLojLKZi4p3MC1WhTaaMgSup7+j4HXmisxUZVB9+sGeu
tx7X7skC9L1aietsV6PYB08EUsPFEjk53nRfrieX5nBv6kFkVDtUAXRbpW5lNyLEITnAD3kKyD5T
dPzXNzpN73LtjKo0q5vXjyMclXQSUyqP0bDoyinRnwfOivZ6cVkup/LAU5S89C/Y4Lep2efs5NGS
FyKdcpJWXL55h7yKzYK40qcqM5birjFGtMMnBB1tdf/hLWUJtb/dAxCapF+dXi4SZHwm0rcFxvMH
Q0/Z6Ntq78E+YdMJUZYagn/0amPcO2za6doh+NKDdqw9EezTjuaV2N0nH5F9lp9pa17snONva/uJ
lhTiNpJ4phM9O3nuw+wHR8CpSOSodm2pN/AcNbLldCYY4qkiS5DRQL1mje3epylEGR8qi/lPUXPZ
0JYQFmG5U+3y0k5qjNEuWtwX1uJcoLnPMcGOwM0uoOf4gRpk6mAzFj0IRcwPAbNAicb5L/IlqSHw
95v82Fdk7ZbIXtnJizyR2XpnBMNPev9xgv5jrGe2vIsHJf/rUcgegBEU5r5LDtAeLY68tn6C5WIs
tTMRwt4QmVEywtReVxUNhBLAN8wKFj35rZRzJTJ459/PPY6fMu/h0xlt1a3m4kROKQaUcpYqAL9v
EghKN5t5PeXpC39WJ/njEvqbuYZLxqVp0/5IjzMOkN3lkKlftXSuYVsnaKjKC00J+hpi3feZH4YP
lTvp29EYd6ej/KQ0010xZSwAUuUVJqBqADbgq1wyY7j07Fb/un/GBentRYpc91yJRTNfk7mkVuN/
fOFk98LFly2knpfooxWPw5VqH2ZWkb2PDNifXeRfFvRPjdXTT6sOwM6i06+2fxfGT/Bvqet5ga4n
j3YEVAY8CNomSXMy4MLkfWLGEGTnDOcsSjtekWE2K+uw9SjgW2vsEkSZalmeG+BdxAu7jBWT+02L
lCE8DxKe3MzAORRk3h3KU0W25DmrBPrss+qvO+ClrGMB6vSQ76vjVelmVI9VM4FfUpYefgNhTiO2
9lRpmABl53U20PvzVuRKA+pVDU8kMZmrNXOZrCvdTCGDYOsYAhqOM6ewsTeN1aX6zprJB22GXRj8
7Z/r/7qlS6Sp2SYk6wIy+z4crsE0wRq+5A/Iox7A0YukqAS71aSe/C4uhY1UmvG796CpJvzAS56x
PneBAj84urKQSb0/ZE0lVekxpGB5xi7x/BYuwSBPHQijFAk5BlnE6j6nxd+RV3CzhQlTs5uscQgN
mAgz/h6SzOWXVlnz8G0h8eTwlhXfz4lWjJK9ugI4LBczCzQDlzoDUjb4WQs6yeaLu8HwqHzsuulD
ZzlZAZY6yE0c6ab0Nkp5r5MfhrbA/Z+LCKH0Upd74rCN4onxcYdps6RcG+uQaXRsT9i3F4Q1yPEs
p2+XwAzq55g8spNmnjLep09SMgsz1zyw7jBkgOGNuRXN4dUc6qRb2jt+4Go9VHcGNQdGECr0Fu8L
fqu5F8Bq0EixiUcRVBckoFgbiloaQgOjEc432utCPTLt9pm2YybCzaoJfY2t80A2fb5hkSO257tR
ORI9ri+N1RZaDYqsbN1vusLiwsGCZcQI5sbIEZKYmem1XXDF/J//nZsBZwqrpBYOmd3Ah9VITW/G
ysFiy3qCedtkngwlSZm89HLIQ1jwH7UTS87BkIY46lLaqF1qxvZosZT6OTV3YAUP9UqFDMHicvug
iC09cLOH8yerSc2p7uN4o5rYNYQzgOR5fxXGmOmWYuA92rtNhr5hqZ6KjwLsplHDaD3dXYBX8Vq8
ZBSWmWdtNLI+cW1bAD6noFAMR4wk2ZtRdnIcddawkjfwQq4wXsjQGvXTFYbUwSEAtr7N0TRwN1iT
jXsURAsfCh8ddEp4beH9A4w8ep7hBpzRL7Q4NCZuyzVI0c2mo1TJt89xcArxvHVvVnQ7NYVCe62L
IudNfzpnvqygbJrIZ8aRl7tfP9n4UFWUab6+Yi/Ja4TZDETkyKbYAV+YxjYIGeMwIddWWHmLOTdn
OYCfpeY1NVsAtMcgHkRxDIUfRR60wHPriKT5W+lTQh/Kigj4FMDM0NIaPFxPovJUaytNnRPwopme
B2wUOqn8E7fCCZsV6CUW2ojDF3At0Av+Wv6hAmGUOnXimzdBzQg4CiO3MGioLTcp1uFNbYdMx63H
PGQJSL/Cs53hgh3epgEPYVbawLgokj94+AJDdsq3uhM8csYxufwVMg01X0umCN2aSud7zGwMu9Av
PKv8uI+cpIj6Y/bk5YLUD/2knxmPOETqgX//ZHt2vYIk+bXLFXFjcRUMhR77ZSHfjF7yVwvIgpwg
3TZEvP7a5JggD16zsdrdA8nZFinlN1hh7KVEQKDGLmLK2rHVzHG5iQbNt51oU1AueL/3Ly5BSga3
Mevv4LDdvbwjlSfQnN9lXbvY3hKL1xamo7p/8ACATrrhKMhfeFusy6KSnjLLQ1AAyFpN8HtNCxkh
0ANZmgQMqIHT6WD3qDzjb/ptgij9rotAnH/ypctnlpzFZjDFYThO80xILAWaxLxWfcu4rumCBvjP
gGENJ51Tqyle0mUOPFWQKCCsEyrnuyEYWAkK+7NupVfFzRlKgGiOjR4zyKdnsKTi2KsWT3/2mfEr
c1p/iu3nuWCFWaEWCPGdQCo5Lm/gadwGEgxW5irHWT3VrnGxF7NSFmoPtgfZUEbXFzDZ1Wj1PLrI
FXjD4uOSOG09uZa0HoTQuT3l5er0/mwRhYs3OQfjvH0zteBWbTP7DVE3WkLmWLAHdFxsSklmUswD
DymicdilbFK2olTNlly1GY1EXXfzVxDT4zCzMhtSbnP67CPT/nM0GTVg2TLeGCQGqEw4ETMVrBt9
y8mLos/OKPCOdniNZB+JAujHjUSK9YX+bX99KoQgHIprdNqXGIaR0Xfatb0cIZZC0bDO3iJfOvuF
JmBEDU/7O43/HSGq3y09CoCIZcl1yiMiDLNYp3R52ZcFRz1hXz5EqogxGZ0cK+m6usffCim8UEu4
SmTiZZYebxFfE6tI6SxNm3yzC8mmK0bzf7o7QU6JvzGxGYPJu/LFcEAqYHlcbPmkx/EY82/Z9MCs
1jc6dB/lBk7CgEVUsE1pgpOqLo9Jw8DSam9vm9/+IJd3mdOjSxJwoh8wkDMcSpJ+ZwHF7H6psdJH
goRyx4Gx7m3IOu4XTLHQEAQvnsDGIO0vCzdu0stwMVCJgtd0JfWRh4AvTo/NnGuc1omjfjJOoGM+
1sDgKxxs5bzBYLzKMPNpelunJ84vGEk580hcLF8iNQB6fMmIuF9GpOqE/Hk94FLF80Vxv6ynYt/8
AwGns/NtpOnU6NN6pIr9/kqZOZ0gGdAV9kEucK+cVMAAdCAsq6RrUepwmONdjgIKYy9GNZhIVByt
kTDcqf3tM+I8cc1T+dXVuaZ5LHIx50mfZXNN6RYl4kiZkZZS1tMWj14YYC//fAEUn8dKavsgxLDD
3Xn4xx+I9XjTFScJGICdr8KE096gEqzqFYLC7kdH/lS/ltch210v+DxqrYaqigjJf00Z9/ruyaWl
RwzlIhIH2DSiGjJlGuq/ZBHNjL5QsRsevNoCQ9PZJ0XnRzKVnOmgN92PTrzzTN5vMoViKJ0gTGC3
hAz1DEWvei+hYbo9dzeBydq0iUDvzrbp1tQbfw5Sr8e2a3m6hrPunuAYE9oGNAxMEvrIV1ndmvbU
d5D2AWVoOILRHtQ2xURYBQG/RpDalNRnPb+pS82i2AokUhNo6Xk90htL3jCTUrZXKMsxDxaoqSni
Wc+xoDgv5x3ybUmSJAr51umH3gIhnu2QORvU3VB8PmReCMuJQgDqYiof9yZ8Zsu+9s7A0keuOCxj
udvnCYCwxCgp9G71BE62un/P2jw9eo/Ui6DkkPfQVqJuDdKPNbIrPO3jVcBACRZ/gpKDkNg/FEoC
Q55bUvJMQXh8trw8ascSf9hJxjtSl4WtwaZQMbEkjMHQaJFyFWoXf5110xRnyzkPl6tNuPpoDxUm
wquQKB7iBxRQGV1hZofTSeA19ard3YdMHYFTscNrz6RxhXb6FB8hWwkBoVvJwgAGuDl2D5reg583
0naXWciJK5J12SrRGJJ5kiRfJ+ZtcmfAL68WYELRTiH4JFBca0DtgrdtLBPkBwx0/7loljmhxmA2
EnRVJHDLCWDvVcvkc/ivVDEHjzXWXkY+wXhWtr5/Lp0HbXFIZDaSc2oDlkIStlA4oUekeLmhjqWe
kCcjwZUOS0LKifqcjiDUmMGny1WZ4LeR1gfe5ptge3wAi7O4I0ZDiDchQ6KedQtaY0+mugX3Qq4w
t6vzKxr1t9zvDBSsRJSYKc05EtReCTGc9At+QsLeMWc1yMSIc8R2mrsyZuXKYYzPHg7C1sSU13cp
xxi0fctfV/rQoQEayGnUDdNRlP+JiEXinuDL+qvKnvtlrppDzspQJIbjhK27ytRnJa21pAERFPrf
GiZRdL7M5EFVRA/jTIly1RmMZ/2deP4Ujnv5CsVo7U1JX8Yz6/MzAc46R0sZlegy67kvFwU7FVRC
rb1F7KkIhVK3Tm0vM+Ukij5WFWwwSaDA0dRoAa9+u+FPzhYhG5ZKuyhuPBeK7ZaDhTrfC45uMF4o
rrGu/CRNaUFew5JR92xqoynDMzn1zHQRNiWusv2R2eHCSgSW5C4Gto+9au2JvhIW3aE4Ulvx/0uE
NUQewuU5zDhiSWHqY+tUTMM1F5AhmVGZB9aNno7smL5Lm76aCaOkDawQbWJ6hgSxFOTzeevBE8Bx
w+1KuzDa//bbGGONz9VcnshrU0RThd6hXo8bqbPPHSTHsoY+92DiEcueYPORxkSxhKyp8407NxU7
ctlx5c8pdJfNWZPudqJsyKVTkd75OVl+9vWOn7PlFsHG+mNp7eVYfbSDiigafbKgxoVSycp5/NgA
raijA4d+EUw2Y9QCcsqGjV8kGuhYxNqJVihWkD8YtQIaySb6pa5w5RI66YuumwqrVNN1UreB/x4r
dTHvf5RtU+2vh+ly8lgWxyAv3xcquUtXeihjvzkVSFudsJ1d8C5iFctsVYOOf4Wist63G1wDI82D
TUftSytpD6rsJEB0Qwirhye2AIx2muIVgOZlAvX8hx6asJiwlrW9dEl1SXkhtXQCd8BKzIgIIUT+
A3TEuw7BRvttvewQhMBIlv3MtmWdWu5cfQczQ7WgfZtAb5jmoFGQc0MAjoLX6Nj7Wib+9a1UGkBH
biqjnr2/jPONivnXBsJM8yI9GwlD4k87PDp8X/yDmkj/Lr3GZe5NPnDkMBwMZm8vcdq8jilYzKo1
fBZkYcMCIGU87Ybr+Y/UH3d3k7IufxuQUd106SvXVbMmoYzm63GgSL8Ya2rrHgKACnBsl/uPBSzd
5qtcAhx8xf4EuM68ZBmkQ+bewBNF2CZWmE0ECtwGZyNqWe9fXKhanZucRfGJpHV6ZHwPIqShGr2W
1XApXVa7K4y9E6wXkqu1dUnefN5nM/EQI7Fsjap2G9PNXoJ1TUoZ6Kig2WGqW54obRkwY9bLF1OB
iUtAWKc4LtYdfaMVrX7X1kmG+E2Tm+C89RSNDbYKynML4jThHH8QShTpDV2h2j97H67dqVNC74HQ
aB78PBlnQPPmKxdu7dkfp4b3O9g+3yEFklc6YjK9Grs3+qO4j9RRkHXVXK+EiNfUAH7xnLju72qX
DANa67JAZZ3HmARB8IU/2oHYnlVEG6X53lksstRGmu5p6zF0uUMlEZbKeBmoYZNQxS9dVoDQ0kX/
NHnek53gXVdc8qT1reveddk+qGaTIrwwRorJ7nRwRTvVn100wNnlvI19NslZQgSmiF6lgD16CvHe
PWX9RicXmSpEcLNd8oowjXg6sU/wysjPSZx3CQGiUMhMQubRg3SiQgwQJu0sHLBHLI3/0wgc3xzi
nAJpAzihEUsA76uq8DyrlIa5csdZ5suBBCFjwUixG25d8uNTOMWCYHgjr/MnwZPiO0rvEcFjHPGe
zhFkE9PgZf57QJFqx2hoxFGj1COzCDbM1ZhOXpKepoml3qLAXqHwXlliX7qx6bI0RjHAhm1a27+d
wlLKGOtbMaZfbojjY8qf7B/iCsdg1NbPGDzKDl42kMm8VLv1RcP01pNiL82fYsdapueydluGwCzW
KdKippBVTLpyOQdaeZm2+CZzoKQJ3XuptbgzWfeOHIQI0K4yu7p0K2PhS/QRmhvZZBYJsJSxsbpj
zWautj7GgQ05QVKANtkURB/J11A+1+DSA/sdUUjLiO6AmJqdhHropbZOzdzd/oO+dQJT35fmqBFN
m9JHLz3L7EnQKCx1ENyzfLodZ82QVLOKaj94fEnuET6QwM8LDDYIyJUEA/Q2wUFf3s5+2HQ6Rl6u
vCDKI7V81xIRUIQeETnQaRZCscnaDdBSWXekbGoJ8CMJzhk0nhjKKQj4RlbvLA4/ptt60KOdbBMy
n1BQPu0Q9t7d2oT3+sC5/pFoUj9XDEI4x052Tbo25drf6WLeUR4iAPyTSl/sN78HnBcf3RbNs9m2
F6eNXmlRgukgjvwuHPEcESm6D31v595yf16ibGPysShxkw4TwrJI/RgiKmrxbi3lmpax9Q+X1DrM
NW/DaAHN2AD/lGSaeOgGwPXDIvI02PuGDlN9/hi1Fq2Ovm2WocsdbmqmJYzlPxS0SNXYSNlWL2RL
UoZHLj3aTb8aYnT6mFp+wlZ+4i8mP3Iv2XR2vwWYcLeubzTevcv8gWjomK/t8DdkYvuJX9qTUL8F
nJIc9z64tLrX9jR5+PW3P4y1VvqvIzZ9pdk1b/Viqwrt1MoeyFfJNDckGOVxrJkC80MnQr2BcVFY
PMQQUXOL7EsvyGtbyWmVjB+qLzGNS6dqsgKv2IfSX8vT9UxisWe9oEL2916HNtzV+zv19XjRkpyt
btE73hEyZbZrvIy26oR2KIFFTHb+GhRZuxGRODnXstkXrgOUcCnmsE86jSkm7xT5JZM5p/bwZLMz
hjOA11cwzvPhjVBhGiscPM7m9lfZtoOvZqDBqBUOAjUKFhmbmt3XXMCQk0thiqYmJp5OVMbCBVei
yNnMZ9hbW9orVQSObXcp4Gy6wmQ3l6x4JdDEs7aDlQXFtiNV9i8elxJaI6BtF8niB1zVAJqRTMIK
3O6f1VhSJUdp9eI8gYMaPOsuhryng9K0TX5i5MolOhkwHusJmmtBjyShwdKTXKGE4lPuAVFXHxKv
A9eQ8FFD4KpIhDDHXx+yHsuS5RLqRlbdlPcmCgLBDHeUYz1W6lGW+vn9tkd5OkbixxDjA5wPJxNR
Whv8zYWaKbquujkSOIASlu7N7xSuMOl80NiWZFK5V/JPo30wFlAvstrCTL0lUirUhw+MUtsHNkde
YCELomOXpil8vPxDFIphx3xEQrHwT/7zETgCouvVGH6Bf4hr7H3GJfa9POuqTH09jaLSrlU3BYXh
2Jv8OMyVgI6m9oRs3bFB8qrDfMwc3bO0WvHIdg1WRrx/u3k2bEqSUBYVZbN2zsUg3+xVopx8aF7X
Zt3SNImLNZ1kLBoJZaehL0Zga9HH7qlEEM3tXCOeKBJInbC3Nu1NiGpDpTItS+TgDHH7t/rSgPij
2BTYvsXH5BKrMlph0amD2ClU3cd/vGP9jAvHsRg+XCK3ZjIMeHAwNHmGGOI57uo08sB1nVoVlgpW
66j57hSlcoUsM/1U3PjhoLn8cedZ17ysoktbK9NCbQjbuucFc1iPXDzT9yYSsqw7B0A9Rcozo8h0
pGQVA00ANVXiq2CXwV0PCJKqMEgHg6qvWTgU1gKQBekUl9akWTqJ8/GGt9qqfDND9Sc7eLgjAm18
IFZFpnHi0KxYKdfzWwv/GQyJAgjcJNuuCrWz61t+nx/a6GStm06zcJn9ugmkwU4k1GZ3bBSAXDmo
q1rvlNxH6kApvN7aPiKy5xfEdNT57OsSOjMZkt/XJJan4JvW+Y4uzMnWhMkJb08T2rFrRNKB4ofw
B37hvDXd7FCcGLFeZRgnobbsVUu3e8bbapVYOse8GruTf2rCkfNRgQRhcqIDY8xskGtn2OtsXx6Z
41GhrARdfXUwePrDv8GG1Q/f5fwqB2Fuv7cv9IibrGmxRdgYk19I/gH4CRCWOQ5RW3RMb1k+lIWs
E6IyRW+gmoMmCU4FrhzriP52tWZ2+hq1Bib2kUPIS7n9qQxgU/GJQcwuGoGVW4N4AnnCrF1b/Txx
v7aD1Zs6p9snZlav4ybCy1iFJL8cj7JY7VvA6SJ+NEvGG2gwU/4vIc0KbwdmE0HfiSPAssVrFUCS
F7QEhsHzN9J5pn/Pnd9L+Q+WMYq6zmYeUYeXazYcGve6ZVpsCs2BnQUlIirPIwtSU6ohgoBSYxr0
DpbFQnNeRigcA8xb3NoskM+Acr7EpFlgkAnURUlKPC1SLiFpaSoyaUycIhFuvXD/rUEPuDMGO6qU
j4W46iTUS3aPHz2yHeXue6opjvL25uzHW0pcbClChDRomw7nVXBbbFFwWNR4O+n/Esjd14/Uf5Sp
cHbwAcaczv5+Iq53AkHTgNxiHCEUUveJXh2P4xxI4HFhzBZqnUogGMWeXNxrDyZ1ajYXmOCMuWBf
Y/Y4ELTe/r2KKL9EOOV1ednsnJf1LDb5THCS8jSWgWcPRRopLBnYR913XuN+YejvK0hOqasCfOKY
SrsiAny6U9PLdHQdOBKxVmzft22WULRm/igsLs96XQI0ID3aOpMVbrn9nc6vA4JAE9hlKP1QiB+Z
f3tZolOukZ8v/nz5ld+qTc5Jr4ndcW+PTOZXg+HB3S20z0v6lx3XT3viz+voy6TI4vxUg2eMLUTG
fty7BM4lYy3Jg00c1fDh/4MR6w+AAjTcULzL8TIszzEjBiAgHE3bw5tP4lihPbLn+N7ghUZnHSqW
iEQGKeYymtBjE6QgaX+FMPy+xH4esBCHW1bQvUXpPne47lpgGSD36S2l/FnWNrxYHwHI0eIglkyg
mPyD0ObrmajjBs6MO1Iy0Z/n+NX/vXGcg7wISr0eg7qKV0wbJi6SH1EGsJMGuRB6QwD1dGWelL2Z
sKM+kg6uU7j31kF5qSP8c8wPlDKr0/rgp8CYO+Rd2vY/RvblF+/4pO0wUWhJQiLdcLgLhHYOlWgw
S9PkybNbZeZFDTk3YUZOi87Di2kDw6NzLTQj2kxSip/o2cT701n8EdxrltmtZVDNV4HGTnKeqGxX
4L+xG3RQKzyxJD69tWBsVsvAfFCpPG3I3rVQ6cqezKXp+Av0fFkofAhJ7qhlq42o4ZaUZy6c6ZVp
UqmxrUdGHmujOQu74HrWwjtUonVj6CIydDC+Z7+jCBzBNCdf/5vcQyR4UuVgFXvfIa78fJz0IfAZ
zCBQtZdE+hFnHos1GZlKjSyDNWPQ91XjKYm9rKclCu18b3GofOini4wt0DmJxa0ofnZk2MZ9N1FU
/Z1Ii7MpGckS6eLhklOve2pQassB8/anUX+P4cofWXPYwg+duPYhHRd+TSDK0e5oaA7G78ZC91YD
L8jtBVaWcG3bVhlapLriAh2lpTKhsie79Mreg1XrfKxjo8+HG1hMZLCgGR5yPJZ5le7EOMzaa5QS
bmzLocY1LSaC3CsTGNhgwvoe7NsHx3CS+k1JymFiQ9ThrPvXo62qQd7S3rcM6LB86JluFdb7Pqn9
4cfRD+n7NHH/j1u872VAAn8SJd7v+yhTeFIdyN/q8mC30LOPyc6xbAqnr5Tn+MUlc2bTN9Xg07Ac
yWOzI651S1qAAYK3VB3dDUljv4XG4joL35CjGH6WW9CKtiGs4eJjKzeNnYKrO6u4Xvqtazc0edWS
cfkVXYWKyhE2/x6qKVuvzbkikddJWrBEUEfhYPStlUGoURC2DLyHWSOy2zsRgYTz9VSJ3+Dxef0V
3XpAFJmOO+fhIxARjr/sQR76tuVKoZgjbee+zo4Dk0+Uq9+YeF28cW+4MS2NTaenFfyfaNmCKjSR
80aF8O5UuT4QaPCzraZVjW0JQ/IiHCOBA73P6XVNPbLYeh8fyFW149CKKHJRVWBTKnaJ2vP6PU8F
HKf2YtIkNpC2iTyyQqEl2109jcgex5iGxn42og/IgXRiuGpvtBY7p3JuHJzR+4etG2j8Ca7vanLM
CGMxzacykKcfn+qQ5Ly/vBRV2NaPC1qj8wK60byrB4sA1Xisb862uLL9sLPmMUS2CIJxtzCcQR1e
gGDswvZRKE3G9XPNRtKoUeTRyqGspJcGaeLB2HfpfYmI/fi/8DIUxzliBv5IaCUr3RVilROCVSoJ
PN8KeiqBZBiVSzp7YxD7i2uo8M868bxj0IzNZAV+Kx7rNWEsqa/72wdtwbZz+cKMwykljYxksJIc
Zt4hHtVy1AcCaBwNUxBgAX0v7MerA9cZPobcesA/jQlJjVXJmVQBfmspnqs11VvXtPF8q1xZoTHU
qOz7NbyRnx6K1FtMqeET/veRimc0AlMPHpwFFwA9EPHv6vXqdx8lSO0iJZO0JfdbJVXFCb6NEXax
ENqtJfVvB0Av7rz3uKYD2zkmjT6AlHTaHp+uDBn2sa4aattFTOEIk4AKYVw3zVmDFh9C2GYm+X/k
oLO4/jVRRxhKaZKebukfWgYrezCdBuMGFfSWTjtxHQI+AhxiftFGt1IhoY2kFf5Yi2b+IZOsj5wB
ZEqatTWksYET8UH2TCIy6SUmhV18eSEbgWnrkMrs92y1QuYeTY08evjW+Cx/ed8fpnYvfowlVOC9
dKQjrqzOfXQ0Jcli9oE0kJOnCCaGHCrj5Q9q2DJ0HQJ2UAGHu9R0O2GD/1TtWXUfCJ8PNNZivro6
ZJDurANk6rK0ZzzX5gsOGIhm08qx7yf1n4T4rfSjNFyD9M/6/LZItnrbKn08w2qpy9P2xN5fHru/
AlZ+i/1NeW4/0SmC1SDSEfqVKx3/uSiBoZjvnEd7D/RF/uJLbWvYSu7Ad2wIuWsBlO4BcdReF74Y
4uWgIzjMOoNrePP/S6xj2L+CLUUeVhQVHCShMevFU8oCXMv0QD06efAZlXUvjLNK9NeOb/boyKqQ
2LSmpDWaC+a/0UslaHimIwOT+VaasTDCHcrF0q1r/fugVaJJeLsIGxSATOFtz2kW1+GOBBArkTBy
nRgqaNZiNqH6579XsqZJvZtwcoG/UQOTcvbSxF6CnJZry1iv7ILh15g28JgKyR7l0z23JEpjO4cN
yPozZoOFSGknB13XIkzuNl8JNwgBqtfX7nM7qENpZIxa1gFJxuhLF9kgvEq06KA+FCILY/FgP97m
scIFQtQq8f6qqkh4/CiKfyjeHzugeNfneFlLvWBa2Dd4eEsBPk4YXIqbTXBekZypCZ7+JELU2We+
mxUXtvQF9v3ikG2iuHsjZPk0Q1eY+fwz3mpBhXH4933tIokoqOcV2axaGpD5mwgqZbvek73bCkkE
ktORrW5EaFpqennYb1AF072Zz950r1POogqza95GiDidNmYHNHgXDWNA0yMOZMqYUf109JEKeieD
uN7cK0iwG7HlO9wbDQovaiHM3EhsO6WnuQ+IGeoa3rb28VNBl0aJlmX2eneavMNImcyxbASORq0V
Q/XHdI/GP0zWYomLZKunFqlvpENIXnVDflDuFvf06mZYnmsmLtvoXwiA3P3FK7w5mWJv4bVJXNj0
JYJZi04Fy0EKOqoqERRuInVYWd2Gsvo/cO/XZKKuxZ9X7ou0m6UI5ypzqgXV5ABixL0g1wO/CNsb
j2mu60y6Ej9FROn9oZJPGxlMa1/qSK7RQOzFaXBly9VMdpcj8xVcUj2bYRWUTckiVuvetPKzgF1t
V+yI8ZN8gULafV5Thcka1WudVZ0y+GWnD/I4Fy62w+iOl6OZsGKBFJApL43harEId8ShOu3LDRNp
mGMb/1IYoBJlWbVC+LWfOKeFb7JavxTh/3HNTafWKy66V3NnO1QjNwT+ew1u/JLeuE8vi4Yyj5v5
DHD4Y2MMP5u4dcaHhsvSrbuDOle7c9QblZn4tha9tE3hT6a2cwhvAe6+cCDhNGEoGwNz3199e2u+
R1fTB8QPU3SJ6/rg5Vm96RdhjEJglTCEiPZ/3bQlJwp+SgF7aPgd3oeZKq3OFeDmWzQ/QMKh3Kj+
qDSe7hNLhIFkT0CUMDh17g+M0ASJUcXqrXABXCYcfZKYeqaGq459EylxE1FYwNROa+3RaSzf6vpg
X0+CNDGNRLcJ1HjT5vK/SnegUrZgTMFIxGR36JRYIpvDISj242/VNW0CO4v+u1LFG6uJ867o3z5q
o1Nuo/og8TM1rYApSjTFcZ52PbzNR9CBJEf8DrvPVyv8msjr3+hXAoZ2V5yI1HPKjFhM3KrTvOiq
ybdn+VDzGg6eDVGzrPaCTQmy18eJbUnmCf0Ur7xwx3fy9KWD1MMFiT4kSzSTdFLDo3Tv7OUckuL2
EYfD0C94ErZrngnkKzcuE345gSOr9Dq5sTJn447bzfvQ2ZbW3SVpt5jHwHMlVbSJV0Q3UHRBsqB1
6u3UGn+7CDiK3/lTJTsvRrfR4eH1Zb/cLx2jFaJ7P4Hcdk/s1qTxkGDMa3snUSjL8rB/PiRn7taj
KoQ6q2gVNa3QxuqQYlS8B4PKCotuy4YC+E4vDVHbYdGVI6h+TCuYUmAcs4aDpLd3piWWfaQEoHUq
OXZG+b/vW9n1PqXT3Ceg88cHiqB0CmZ2LaDAUhYKmM40x9gMm9A6GQAvZmLY3GSVZOsKfySRossq
5rVMMW4pmPXl4e8jCRMAY1Rrf0nHP2VZOEh7EQBNx8zMmGCSaiYNKNZdwftYY9RlOnqdyB2q8dbS
knhvr5hKDuprK3aAigLubjhPAaWGPxDhsENgjK0qPhAeTiGscwRZ/Rk2ALlLfvBYH0gi60+eeLTh
POo2PpPPChBNxw+Kd1FAUpf2FAHOknYdsRlqCUREl5Igu9cFJ7W1NRhd6DXwkJj1pi/OMWsMPhVN
Mi9PGs18M8dT8+S8Ui6n4AjUt0/NXN4kCl2lnSP2Do5vgpfmzKur76t5iVlgvkVGSSbXQAOZjoAN
lCz33k99qVixmmtSdLyY2rkHTdw/TKlO/GrHDXwl69meFD7IoLgvhvQbSfKKQGern4ZrqwbQY4Iu
dbuXrcriCMSWevbpesg15SfrGe09AF54JXgwLYZ/rIOyh/CeMQr93tC+X2R/tnYD8tTamUnUg/yw
1E/AXa7ZHcfskYgzl2eltSuH/cwvvkr2GBhzdoTalmhBy5EHUgmV/PjwE5YZ98+ljWvN6URTOXVp
4mm1gr5yNJXHR39eO4VnDM8VdKqvC3cWBxUgSoB0R0nwVrcVexB6PfjdXvqi3gBF3vpH/F0vOZV8
Um80L7fKvS1GllSR8oyIENPi4FUQqXCgBu7j6bTGDfpFLsy1/ByTGP/uiPQ04uc6mwCMkoi8NED4
zgeGnYvNo1H4wVG/rAg++zeEeERJoB195DUttX8mWC40QUy1V/MCMyI/bSz+VPUuZtBifD0knzZ+
hLmR/IfBHoKZwBrejGMAl8hKQ9mwMRbOM2omK3jnqqTOXjfsWQgTCzg3IPfvsfQw89IzuZ+44y2u
3+MedICvPb8Q9dkJOC8HFo2Zuv7g+a3DqyD6xUo0V+lJuxQ0hct5MYaetsWWtyBWD0s/iQqf6DvH
ykAdBHy/aElQi4ztJ+w0JTU9XQwHgDJF35KF8em71Bp0Ml6VOBdu/nncWDmUWA8+uodl35ARcra1
PPTQKRbBMzUXz9bx6ALCPVlQyQHmybkcraIrKeGwt9koyCnw1kFE7eSj0AzozNIlwIVFQvr0MVBx
+s/EFSKvkU1/P2wYvVOyWmYt8788F9rfNbDlG7H/Lrn1vML2xOfuak6j3Kzh7ugxw2y8uflAsHXE
z/+nwQqjYXncMMzRou4tI5/Vh+KEYwKkoUqyXzy2cyQshUfgLGbNKsMagAojGIJjQjtj+NYrRGo/
xV1AsZPMS3YvGi+jiVTsE5hEAWxns7gDsp5cfg92Mc0pXLE4xeB+5b/+JY7U98TQmyILSmyOwRl2
qMCTXRKtOJdyAhTzcoOJP4YfdkY9BZJYa5QZYJF0udejiGl3LT7L+0YirTatS4Rlt3fOsbWPzJzq
RmjodCeeCJ2PY0FWUsxhtjyY7hppYvTklvlchIIl0caZQ+Iw3ArNkg+eOKvY7tDGILn+sDvjCQLB
/0UnejnA987jjZRx5juSUknguyX7jTr+ma3icD5Azi0/cO7J29zWgxkkVQb3A5eUnxg6+uIUCL4n
9UOBzSUozo+J6duu2CAeyrHJZDyoRmmZvlL9kw2tP39EuLFWdGzlpJwUMK7GJV5KMOzEdDPIk90s
fwDRXOXC2PTMq/eD4HRWYQvmiuQ1LK6INuhQ/1QtK3Cw/tf3t2/OmfsQhjzSJFfccxHpGZNB/5od
FHbKyLtkrUTh60z81B88sEinHSPUixGcf97mquI3cOztx80qhi6ojH6MHMwxrWpQ4B7L1XaxUsMy
dY11mOjR+6nVN2ptxQn42LE7yTq51neUYL5SktH5rA55mHP5WAvUUf15xFFrJAt48/LLwjODoZzY
UaCSSqivea2yTF5rb+Kom2qsLhxZJOZTsXvHBIWlNwjF8dzVX6fKDofAoL5EZp4qXWeSDNXTi6xj
go2FTSbq8QgDbMAZ2O57PDgVqXMaLNSSsGCqZc2D78EWjuGTj9AxoGcU5c16YEuiNlqru5QuQ1fl
XIeP19HYL0pL1Dh5wflPMj2Rk30c9g3jtNBPuIR4wLRTs/7ypWu83rCpHevC0NGLvGFECDhR8Dgt
qCQjMJp3k0TC0k7H6hu3R1qBDXkxMkiDjV6a7UIjGp6A8zHzt4MeGKJtP7e2/csV5mHG+QKlvWIw
XhkfwLlMHv2Bd/esyGhzZ0L3H0PJer6ANekniPPl1z3ROa4ceamWiP6hxMkLcDTzp6wCiTihbFEB
sSW/bWga21zBjKtMKWa3kj39li8qQnPClyoxcMVJXCJZ/U6ieWIarjZ6UsalTg8ZCc2v4ThkH4yT
awMGGef7fU8Mqpgshqf1DnGZLlRarlgdep3nKTftPwVKdeadThIygC8bNa2cWxhwOb6vbETvfYEy
QrsKlS7VdwOvlS33Esjf3aEgeoKiT2v6AYgIJeEEQnW1c+/HisPIhJbIJ9XcOhaNVzYYrjdVnc1K
/2a/ZEgq1VwyB+czhM1gthic9XgTFRfcsgy5O2pWfAdoglpsS1QnXg7viUg5ONIOI3joTCVj7JeY
HrHTdNkfNmi92snRARWWm/nALCTYyqMYQ/IxaQs+rUOJNjannF72FvhrQ/EBWqfuhaG3D9OO4IWQ
bs6w66z7H/GXuJT5Ro08B9R7OhvqhIBVfRYmHHzX1cRhvtVoZV1LGiMgjtacfmBHRBbExppl2tCc
rRYaov9MFSAyaNePBY+cGvv4uo7sd7bhRKAyhSJRSCn976Xi8Bw8qDdAJna0kACtdQpCRyCJi9/o
ttZQ5nQ=
`protect end_protected
