-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
snOZz15/e/URKoNCLpx4S7EUPcb3+yKKy64yX1UVanvCcIpOTpC9pVyJwZGkuZOkyBSK7i6sGgcd
2MS1CTrfseQHff5q3vvq9rtAAKUMRaCKHXuec94DgnK29Gya08hT18aB3XkD1sklJ2sXL6kHPOYL
16OQmfpPyTR4VAZPtJRnkCYL746QwGutfXLwCwjKMnfHi4sw0SuP8qnMVc5wFCByxhN66Ky/OQHr
qO26XapBkqTqy0H9IaPflzdiIHa980/XsDjtQj4LjPnpwWvxT3x5uKFLzfyAllCXbKd6L3RDcSlE
CfrLC7D9b9l7DKP5pUQ4bjyqPTn0Owue3uN7DA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17024)
`protect data_block
dykSvjFPld7+qaZUQQd8hDtpAPNkBL2yO8zjAqvycqWICitJIQmqi4j+rmTFIlkUkyVBmWT/FnNW
SOf9DEfdsm+7aeMM/+Me2cqvc/jkRcsA/Vvjc7mFZIP5ZZRmu/TX3TziA8ykfxcIXjXwgA++IAON
yQ2HDYNyuJBzPS9bBbAgmwDG53rz9SvoQ3ibyiSDJGu5udB+T8vJqpO8SEdzjvxf+TdpqmwURY4C
78m5glrQ1dUah4HH7HOR/uagdn7fSdYihiz989T1eIw/iFN4tDJWg12wgbjjeUJkWZrhl+6Hg/8P
CpAx3Vlp/PDS5BEclVl2XzYnGZnbQhQDDwMbBa+8AzswZIzaipBqMhFaFPCB0jrq14Jx4LLXNbnW
gB1RnEFrmgGPn5qQRwWUy2klz8TicH+lO3f4Aw8wq7ncQd0HHZhVz+sAY5E/CwqouumCNEhalx/e
ppzBkFTjJEII6J9yozWT7zp8t+k4R69L1diJJHJZ8hlBs1XCJbeQ8oDwlZI8uxWmcT7iw+YE7DYo
3rGwtHJSNqVwGPNv78XcYKZ9PJI4j6RmsDD5Jc/lp7AR9YFgT89DdKZJWecdRgTMkUu32w7lgtQu
W+ZroxjRWcMuTJql97bJqxO5ANzldS8Qw6IC1BQPmbH3woAUU8YAuJJgI7KUKSur+65A9bG56zAw
maEiAAC614vH1POWPWlwR8TbVegmTNwfvrTKxIw6kMoeF4GRws3t9ftSKulUp90TB+6UOzIGqq78
3hmzVE0FI4KXW2vVLssoAY/thQL3PKScQFzjGKLq3L2q8FaWtR9kQjmjZllUvfUrjupmX17DcTd0
AfYnP0iM700/LKADLOfj0dU3x1/lTdxT3WIfqg4ugSiRyqMfj84vmtFcW2lDu89yS4iNLvM5b8FU
kG45zfOlozg77T7XQVxY+2zlvI8nWOII89d9jRpgRxMac/2q8H/UjYBTaVPMGvcca7X5Ek7fh+dp
ifZg6JhrvDGCn6lKzeehw5hWSOjce8zLHgybUslDI27+HOtp+AG6Pu9lj5SN1opi8GD2WGfu9ur0
a3oLbb/A1nPq/DQwkYJW5WNIr/CakLU8YYPFX1z90xUqiHmAlDyyGu3xzwfOT+/GAE3aXc63mBye
1boaOfS5O3t/uVpgCltoRoMfHtHl58Zw4HiEC9V8A0qSZHxSmP6ryJxV1UHVo3T7DZk35+chejc8
mw7RxygH37x5YMvSIJ47pDnJdmLs818gj7HTNlZwZZQKKIiIvzapYe9gSQIWcLGHCMtVD/XeLxC/
5lfHjU5ttJ1dc1TzKbRzNHJNJ0xe25UDv/1VrUDecSBTisLOXzmtu5molCTtHiinDCEEF3hf3ppz
ee32PYbN3hBtb0P8V5t5tHT4MHWUtMuifrDhhuPYI+bioPk4fBOqg1dGPma552DM40IVuSNNFNH+
l6+GfiU+Gr8QkUCaRSxrFBqqJSOHVGq58f9NiFMWCF8YE2caG3tTni8oxsneattX++RN7H/V54a1
rwbmkME+dJxaJp836Gs5dWHewrRANWyNyyxTqtyOAiUElMjktJGSWNClwHCMo4LVzULXWjzl4J9v
19BJYcjLPsjnQlPXAXu9TfnMeeiGhei1nWNbqWGrvdfZdhhUm6+OHa+6prifrSyqJbSLX2dOHwg5
TtWhatw86I5m8hIeUlgqbhHXogaoo7pGH9YZiPZ1202rek1Ald5REXl0V8iqapd3Rmdkl7W/q2XR
z+BtYvH3I+cKdwY8JZ7Qu9PbdHcycoAAENYSARM1Aljc5AlTVCml+xB7v5gZ4sUSrr3BhKtIXJYx
cC5xitb6POfYF8m8KZkHvfVWVu00e/PBIv9P1gktUe4iINByBQWb8fnPreV68Yp4plmexueDt99f
er09PIUsmU5T11/KBwrJqxv/CIH6GRST9oyyU0J4L6qzpVnXJ+BDoaGl/v3/axMENoQXajofbd5u
M/zf96G02DpnUDqmD0lMKmtat+hHCTXwrisMug7qyZbui4ynyoiYtOi3FeR1ZT/jDnV5GykktmR/
k2dHPazuVl9eG6Se2sjsZ+S8JnUfXb8ZdQmrGt/BQ3z2JLP9Wa5rxpynaism1D2j7koF4gNmi46u
fatbhApUQARX5BIGswqAePHSpoKUhhvqnCVpk3qdiMvWzZT3xjplo6fP7S4k+CmoF4/rzOLQteA/
AfRHgu03/Fo7+BHm20lciZQENzBuAP1oT382+ookUp+BWvvOO8ofCM+nKYHnwAVPQ4NfBovtKBqC
Kl58Vwwg5FxJyaIQOOfX5xKd9CTBYLjWVczSR9wGc3ActjGaF5tGk/jeQ+QtXyGh2PctQvhZCSoD
HL2o4W7hQ3XvzCiyVAPI5Dy+RdF7odb2F2iNgzn7+pCeYF8sSjHraXt4Lkd51U+a/pvkdcrSUKLl
8aTeaCizUlQnkaWe3Pfv/NeYwjAmFZmQeNsIYHrb6lAJiP/eQJogppXF4n1QIwS0K5OxKOoSu3TL
xpWdoTDKoLkUluCTyxhZD1XDTQ4gIK9lMGncaZwXhf6NFiYH2DC6gthDGHZZrx89Kw9zNJFMLk51
g8Ia7CKe+Icqrjz/jHnwCQoayqrogYXN78r8zwX+zxm3OpFdJISnxY+CClO29FmTOQdFbi8qE7zY
ZxSHIkZl2Y6nP3Ut9ByLCaKk1N41uA2miLUCCZYh9kPLt89nYIMtRIqFe7pq3RxzWwdV4+k82tDu
HcpWsKsbFADgO/p2NQatFoQafIbP2Cv/rU+b94y1UvCJkH012pUdNxbT6kd8hBzMHbBeOmkV3BtC
pcLbxgpd8Z6U2Rmm4KyHIH7b9VRwF8HSUATrqLZEYgQg6H8bjGtjnWRk1/u1RYgCM/ayQqwF1QNI
dpJsZnDQCo8hOW00hY0S6WV85EwyoJcVRj0L9KXYy8nY74NLfozonUR0l8nmHBq8CmVg12F2EcKE
H6MoTYqUrTpuZy5V40vcUjyi+N+Sd2wNnRLtPxcnKRey/ljI8TaRgClT475jAH7aK7vgVV53eCUw
dfJtsistM0qHqgiBX9aT7ZiXT5o/jz5xOHtubB96g7b46IPhPyKF+aA4U7yFD6LIBW67+X4oUVN6
C+wHUx9YCf/9rbR2EYyH8XN7u8c5HWD4xZXpZ/VvtNgVLUvxTokJYhfphPOXnvEx086Id8ZRjemA
81Be81pBdhg2LypHO5ujwrhhn8QEff7LrUY+C0v42w1FRIPrhBwllzjMlb5c/vRY3oY3sWlRcjqC
kLye2Q/5Elv/fbnZFLstLhlVH8ys2BjKPaQ12S128a5plOyBJ9wNhCC40WPfgg1EdSsDK5hnZT8Q
LE8HK0w4dZtCk+9FiXd8fgGRejJ/9rIfZGQCZ/adOJ6RIe+USbuuGoTzQytLe7H8UsVSVnH1PzTH
TLYIUL7X41sGRd6kPanHRvHPzUd1Qi3b3S6HVzmFzTNy5lfqkPnvLsLyV2KYTC6chBcMxjvvApVE
kdaMt+hdqJaoYad9SY4JLIXpl/xSySsFrjz0eJEh1/2pT5S4OZjjHCNF7B13t13mZi7MkBBzTh4B
MfTRpd1mKvnrqJbVQaXRZwNL8pn2uustjuZNk1Fvx/dXUSlKQyd/D/wxr5TUMXBP5TL85M9SLpRR
paEw71pv8OFC5vt+a0lGnBJM29FETofcMIpoXBQ+M7Ge1KzPXjWDBH0/NnOOfznHE/ZoeignogmA
8AT0O73V5e2cOqSmvORk/LwevE03DTcWZRVgvvncogNjXcUKSxAXljmoAWYIY2LpjEIhlx10ZWMa
0EGnKQBSpmXOvoKD+Je+Y6W2JBi1SwA+HW0qVnCjpDygrxDxlgA0FHCauZJxbzExxFkNmR4TdOji
wAaGZwV5COwLnMA3Ec6OpGUqmYLRju86fSb+6Li8QwtlmCSi58YDo0k/9TrCzI53Tz1mQdqMaDW5
/+01UD3u7e9Xetn0oiKsBSLDI4yxHXVjyf7wKgwo16YXA87p0J78kjM3VtHG2MplZpiJUj5w0F0f
8IANo6fifLEru8fqrY0Iy1JNMgCL+pltUG+JzUVzTfpnkheiwiDLPH48GQH06KmeqmyzifaejTbm
bO4vD4vppuuU1a8mn1w68iqEAmCy+7erpej3NBn9DFQYP6GGoT7HPfN7ThZAaaWiOmf56207K9DO
uQEBZe9qaYcNfXULKwXV7+BfsXzQMQ3ooMRo+VIx8LfPQTkU1pIChxdobNPKaf69nZwJnUofsb+2
g6o3orYPhSZoDn6Jy9ZEjsfGHtnWQTL4ZZaY6O7/G8/bZZ5SNg+aaRYXrreYva2BkYgi56ZJik5h
1hE80rFAQkO4m9ZKzCq63MlHhKppbe2tC740UImFUjop09Eye070sD590qhiINRHjw6jgRkUPkdA
W+n8CQvw9PK0omQ2udw7daldVKjL/DRPlmQaRnrfgVCs6qq0DTfwaW2fTqwLqhyALkndgpQOB2GW
EAhsLTlUxDb6cYdO9utsX2pBC/EufY4ukvtKspvZPcOEw8IQNjhlt/qE1GZLxEtbtuLS3e4a+7bv
H4cRC13KKdMTa5WNhRdVMe7zwkIprf2I3y8yymZ6fTG8cMveXT+fwXtF8UMwS3I8o7y8AMRi1HsK
bmr5NiDWoFnZLP53PHo9g0BIEtqji05ZO0GakcA4ryDCfghdwzPp8gbc3Xs/jZzeU/XUj8CG/VfX
N8NvURb9OUcGqG4CwW1EPwc4iOnZnjYEvTQDoEqO+GARnCoAN3uO2nISZLahNYEoV9gXOk6YqndA
SZO6Qx4P6Noly2M35dbfSpB5+82SBBrjYtOqGMQaWepSd8Qkdo1ChLbkhkIXyY/GeBhx4IWQahTc
bLZsRUDD0AZX01pkRwNTKiwgXCYMduW62Lij5keqZeiD0W7FPMlQ7laOfvo4lZUkyqu9UIQqGf3Z
uFD1Dqltne2Ndfek5oBUisQzPr0H5+kNdX7gVGdxKXqxoDXrwOvsuR5HOrHRolwj8ycjnbNx4VY1
QwnbHhk/x6Cl5DltXftrzrqGW4PT+iPGLUOUeTeL8BlpskGlj8LZFerO9F+fE6lnh92ILk2e69YR
AGncCTZCanT9V3CZPtAINHcPPE/y17d8Rug4WseLWgDF8UlFQKPS2gFTm6QDiIBI6Lwc2V0IK9Jd
Pqe4Hhtcckf/SMATCBd5mN7bdvivQRCNXlxUWVkl7iGutGJAe9KIBKOOtieGwTa26Pf1lwB4ynyd
1clougnA7s5S7MkZDlpARWu+FyqJWAMoUx38e0jelYB3KheCR+LatAK38y4/vtK/gbzHd3sxK2aQ
82zGthH50jA3LGXLuHqhiWE5IjvaTCvExTcdAOTkgCLn4772wPh87JYerjSli1oRiOLQHBRCD+86
BdNKV40B1h8DwYnZMrHkfMEonZ+HvTbFcmVho5k3lH8zGQByumoQQhzjGNed121XaMYMkzcqKsKf
hctaOSLINT6d7bU2dAlsruaUR/LQd1v5kW4SVc9/U97NdmkrAJxQaHkxYAF6o2EgRE1XK9XiJklP
sWszuqjx+8kXZbB0Xe1fVm+s/tAA6LNkViONQiWPjaavEAIvtnBmLJavz9GXYdQfcEZlUvOeL8wb
kTzx4r0ytwWbJimp3/tQ3jCQgtoVDHKjy/uBcZVQn9T5iwswh52p69vOg78zP90jpqlU/B0Q/x+A
12tt7BQ1LBaDi1MrUo8ydW/oWoYUFa9Luj4SuPeHe1/Jw1pIPb7rL77e7CO11TAHqJLDGuXXsKQ2
IcJk3j4ypV2GIFGZmKkpHUK0syXN1OaHt4BX/2cLkKm83rcU7xAnGReVqHnM982obUyXtWeL0t08
uePlmRzHHJzmgfkkwcFFaC+6DvfnqtZoWGVtwKMHUfUzojuPuVXeZ7F4ncXlsOOvMQIU20dcYBly
EJOGQQnkAkF0v8yZByNcVJlWyS6nwaEBqP6VN9if97ph/LiynV4GZ4JGK34WyFOPOI7tc7IsZ1Wz
8aAZyNNg8FGSJaSQ97D6d2bzAux7fP2rspPYJMyTpzF4fP8+hubR9xIFEKznLxEk/rWNrE2XJrRW
xKQy+lusNU1m3o8iqAWbS7zNLJKbf5ptdT7TsNwrXWFeuA1sARN3BZbP8kHw+gKwK/X2QEpo1InV
JlecdYC/Yxs9gdkCqWPLrs5guOAm7CUcSbaz9h9MWzm0hwVpt0hBrmjhcpFjDhkOWN7oeT4l5RlP
0HUkjtRAXdDcFNIotHl8zZKGJ4eBl1k20n9I3q1kanGo0z/KYstl5dK6zr5Ihk2VEgAx8DPeDb/1
U8olgHheOpUBQjESCbHilDFdelzEOt/o9EaPSp/S8zwWFQH85srp3q3kEoXUO0ff3ey2f7AeIRjA
y7/Pag/mU9pO3arXHRpTD789bGchciXm9JzcOyi+oUA/Rc2yuIFhWZyLx+RXDlpdJqg/Bc4i980L
U41jUvd9S6us56JMI8d5kU0WOaXJ7GpervBBkAK+yx92sPqWKOXMXcOjoo1i/SqNS0Q3hLtOvdDd
o+hgLFBtltsssu9WD+G/ppxca8pEbJDzbVxuBb08OkV6j1K4OSolDIsMisiQ6Pwnbpc78mHK6MfB
18N56xI7zoFvxBITjs/V82mRozcblTgq+qNA4xkPW2yhppTHJrXRE9hFx68UBU/dFSbebNfRVC9f
3FWauSBsjYyA67yv3u1EwxCj0VLgRZXp6JMIJrfhFwAxfWVUCTYACsQmX0RgQ94pfxJKlk4+4maN
H27Oq3sZUXTfhCdBb2nDIPDMnk53cAxELN0o5Kt6m0rJ6w/qM9YxCeRCr8ea/JOZHttOqBXlBi8X
8bJ5hmnG6gJ0SjPJa6ePLsRJSoT9Fzbsm2LhdvAFr5qUIaqLxNv9SxjA5Me0AnT/imx5UcbzAZqL
hrLjBijd0QQl8qy33f92LEGB1xqDBdbjAnTz4zKYPK1pmDvRevdLXDEVRIE2ak5UWDF0Mi++dFlj
wufsHMKumJW4lKz8MUhPhdw84AlGNFe1+CCi3/zBHS84B782dgAr6Rtv6HEyENCnkhvoqF/wmeJi
1TUC5Sj7uoGOAl5iTU9lS/df9sJfGYq+JaKFGH1KeWa209Mh/BeiovxnHubdEkL8vGSwtqmBxzjs
jU1glCQS4CgCuNx2/QVuFtrR7j2cKXI6sK0RQgbxJ+4Xlm47OYvQr0FHqDiHLlqki+76knPu/q4b
V1TB6AsaOVv+8+FWt0nTwJlu+SbdLShwQ9d9nJs0Jp9dYwXQTVaeqaWtB2e4qwlcxL+rIwuYGaFF
PG8pKmkh+uIM6xiURID25FfqukU6RaM6CFXnUwMR/SYojP4J9LRK/UTY6okHhAKMNIO5qKpLoeIY
hANdgcLydFsZrDmMq6zFYcA9751WW2LYTm04gjOtQVqYHG/+Y+I+6URrxcZwSNZr3uYtDzVixvVu
qKNGhC3W8iDO8eu8bPfjoTBbCZ63cIeZIwcYEfDrwmu5JvKUJx3oSJ3JBdUJIJgvB9s4u4/utRZv
8qghy+3LTevjxZveI3JmOJ0Ha3tsqGL85TLC5UhR9CzGUJvdDNGiMaRlPSF0Jk7VcLpyN+Ac/KKz
sjIgJU7Ob2DPZz5TL8OLkg4IzlPuhTaqbtyl2XnqSMg6PdmIvnkHp38Jz69GPlQWcX8e+C+f2fN7
2gMchpRgXC77xPffmortSx8K8DYJDHixj1mbx83MeXWDRRWQacFyG+sCgzTgNGTo44SOBYktA2rx
eULp5s4c7WVFUb2y46M6fa29MECQnIx4kEmXnVRow4BfrHyF/4nbveWdX47Z/3t0uadvHULTIrly
t4xxa89vAh3EQGBVD+ilM97ixrjNohV2+3wU0gWyyad0ChRpYPdUTLICwS0INlOyLyD56gMJYaCh
Ca7VSKrAhfR4zCE2gU+yy6Z1FFHX8p9jTO0fEKzuFifYri983YQdIX03vSLmVmkipc/Ajq1KX5xa
C1Ock2KSa+x/D9+gBHW/Y7EUdLSCER/FyD0ajk4lOcDhXmPj7GeheVJzh22Fa4OXGaOJIvx+3Fm6
F4zhyNEi6fUPOSdWafhh6oQDr6x+n2W2c5EIdTCz58LzYkl2DLhAdAPDLKwWTmv2esShlLqSjKP1
AdDnasr2y67efoUysxy1ibu1rKcpEj/mxsi/uLF/RbTvwDkxvCXuQIf0yXH0zpfbXbDSx05O/kyJ
yaQBciqtYy9C6D0xuobEG9BU2/ZCplh2dQplN8eRfL3lIl7kzNkGmLktIdgk9/8gVFNomSl/4Nom
Mb0h3zGNketkNEOPhTqr6rYwkrGXrKryy3aOnnLTZtpe4kOwfrCeKQT+fDRRRmafAdIBK6y0Y71I
5La7GRShjBxgIsTYxMGfdqWTzvxy3vnH/KG4nRFyCHG6UqtvE6Api2rSUh0ueqz6BObVKeai6FUL
MToV+QhTvKmfztVjteY3R7PhQe8mRUueaB9zkO1cT/IgB+Go38KDARll+k6pGzmMZRe5QyLaA87f
zDn0klSyZDj0qNbMNXNsu8085z1O+zjt8WNRF97/5AVFCEaUTshlZdkWYlm2uo+Ks8M40hEiP6ZL
uEKrNYG31lCm4R7l3EUqfYVwTaAd2AinbwkAvH8mQnyy4TTFlqtcrY0GeDzYDPahfu8Ga05v02Ho
65v0hl3FCW8gsMcs7bIMTVyIwtOoFDWpPvmlvEC6vHbVq83jR93ZZlOMJQ1zdPMRsbtY6zJYUcva
HsSurYhnvPvtn/yuHUXUHczHmLQzUcSUnwZbQtUuc//rk5iUoPlukdtGyxzJ1rpOTOT/qUxKofPo
tgkSPv90xqj+o2iT9n2O1E2xwuabi3yCHIwOQh6FwvBkXVc+hkOrqMrTgYquJoa1mjHpC+iEX0Jq
ENQPvtZua5zvZaSodqVejK/MBCaqSwtgD1SfsKT6cL8nBR/xFbd61Y6fMySmHyw94w6o3S3URxE2
3qVBSty0p9M9sBylYspPG/anfWR1JY/KCvnmObzS6crXljUGTlLEbX55oG+iNM7ZDgNrnKSrIXsb
naQ5820/Y8UbDvGTSE3beo7Ee4x5+vXViBMnj8VInSAi1/fadboRAwSnyRi3y8EW7dplSglLOd6C
D9RZhMvt81vkLYGy3x2h26vE4PbOjaiFkBWl1Of1hNLOEehbwq1SGivt3dDn046fvPhn/Ugd9tnj
iZhqLbYMRzCFlZKr3WJ8Uq53hOf/6syAkQGOYkJUmrwn1j9Db7xywFRryhO2olUtS1HXvOJ99yWb
K2o+vBhbA8ZmgqLki+EuMIFaILfJgTvf2TVAtXmmoIaKcc+YgWhHWfqTEk3FKuLTDC7qlS+SHvO2
tyubideuWbt3u9nnQuQLC44EvPOZl/xq6eyi5S2PgN1VlptvarJZSr34qA61Z59tb2e0cMRdBe5O
E9HKpqTLEy2JFOWWU2xUAUCN+c+ladnrJwCrSEUaL47GpKOndePRtoxER4y6tBM0eAcDT8NdB10g
7+42hAKoki1Kqmvs4AulZRpqxdEkokxzOA4qSmU0ZWZKWGwMYMLiCjhu+WrW7cnTCD9F40AgF0Tt
8jKLdPozaK4if9kZ2Y5gME5LeaEtL2KglssvU03l12TPpAI20LPYAhslLLzM0lfd5u5juBOaNkQa
SYuE5x+hz6ZkP91RxaWehH7NF+WuOsb+xb946X3FTiUqs0BacQbC89a/QNCOtmhFjOP8uZwG+Ahr
k59ysP7LdGXgIDntWb9rl85vaEpastH0h+w5Lv/2KG3LN3unJMQi2yvpn65jFzm50LjIf9Qiu/OU
kt7ckKkTnl+5vut3xPyfQuV+4NksSG1r2NJKI4tCNA/s/odHpOrLFBulXL4Emby690aaLacBtD4I
1gCh2fq4s9LiRhvCRPO0hmC9S4HiuDDMrjPAQS/xS2z2nhzRrZ+/4axnHThHXmfrrp36no51LNer
DHf/kbFTE+4j5Ib77fBchQpBUjKTG1ubR4oPTyK6MFNGKJ6Z19jRd7bMB2dnO4EwKaNKhhFjKgFT
D73IyfSe3HAOa3AT2NM0FoLEP2/dT//I/G3zJIj5IfVcC32i5OgcmXaZ9b9EsrrqTnsCWVDN8nGx
BHEvT7MBVa9rWnm+fGlNwmZoii+TsqhpNRmJE+NJeRdK1MVtLF4bedL6V+PaYWKGyHU5L5ezdzRd
WKXSzJNfOyI1fRoMqQSGftC5v+wdZNR/zntyjplFq/LSOkqaE+4z+S1Otn8C+eqgBbtc7v37tzYV
kpTd20MiXBaxvRM+KR1TdoPvPCtRPuu9AWF5dekhnbMQLYVjM50jiasSOufNX0QxMDrquq/jwWrh
mNZNKeZkkq53HOIsd8yXG49CLuFSyplmSTVL4rhOCIZfIAV787TzHri9YYC5wP1Xcl+ZGitzdeea
zMtoJq3eIiQDriH8v6aTkJfunrZSsI2Pz0tWZPTHN36eOhuUVon+NBDw4KA+dIFZSLtjAAfep0Ri
YhH2W2bzWL0oY2zZ6EzVaZr9uGq0nrvRE2YP0TFxmtxVm3u7QxVA9LRB0a+cEwKuLes3E2ELGgpX
R9/7DLgZ1BU70DRrBkku5r9lW3Cu/llQle2rOgKUV1vUEyXnbwqDTAK54wBtmoj0JOCD+BRzGOEr
vrtz1cc6FuVuJLO9tUOImNwlrLZguIOB89g7m0McQc+55yhyNkXoGdeT0AFU2S25GXtE3IzpL52P
JiKN2A1MJ2CrhZeNDzIKUhSCVvQnRO2PAQk0pvY98PoDsGrP9PC2dBJPLOewF53KH4orZ0n74k4K
P4fao1VR7xncYF4MHfOs5lDswO0dCG5kZQSjGQ6egwiJR1Cc9WI/4LBgJrK0pfbwIzeZ7x4TMH8o
Fm1qhiie8afVuCfgHH42wrNN8uGvdhRV6tQLeqT8j0FP+AmgoTXYipHNPMBRi+bnXCdkGNRFyUU8
bZoEAgfQ3M6+ObCMe73gRliOhQSph3YE9WQTR9qcogxr7U+8RKQeytjG5taR2v6BlxFP/Ldi1Cgl
g1dJIha+KIxNnHAPdElSTImluN8geHuHQp9Z9sK/QnmB4rR/gCOhnCPrdn07esxgGb4w/5+xlfh3
GptT4kRxPEI4+Thz8Dt35uB6JSFUSVSTeFG3QRTpUDb/iTlgWUVrDDVKGryZZ2QfRnvV6ybWPa8R
KaEP89+6FQ51RqziGjb2HUVfE1JtE8B+ryDhx6heHSWsJVdsx5i9AQXHTBvG1/UWsd17D7e2kB5i
L8Rto5XI6wwYLF89FM53llS3iwkeEUsY4f4/lhYAmMSA6tQ0eEQMpe5FKVmlI/6pJoiN1f6uRh1W
5lR5AJqkGpHmRQGmVzO3Hfo5Jj7mLNcc6ot394d9Ug7bYtT2JsG8ZtuW3iEgqnctEf+JlJwD8rCE
O+Nv1zENMrf4WQnFPqpL2CaCSYnBM3Ojz//PAHG/Id0+PlgIKk1pvl7ANPPX4MEw037IvFVUylmI
e2KPs3CGNRp8rTmSGkXaMM+4Rpox6XHlAXVjInL1aUVCn+zEkEHAaH0uGZutGDWmtSJzYeC0Za9L
EWolnsP+5Uy2V54UdzPeyLeSl9W3BzCRx1gVSf4tg/rT0kHWeWo5DDHdl6y1Ihlp62URRbiGJGuq
U6rnFptIE9QTN9JwfQxgJ1EQ9O2oStwJOwwJupsogUIsJKNcqhdjraGBZ0lNA/RxrnlLBCojRssi
ldOy7kQxBNNkLOQkmrEEZmVBLAawVSn58Kb7ahnR+3EZP3FNNJ8WLDR0vzfZVF+lR/YyMdi1u7lU
O6NtmCjG02U1lKodyoHzbicql3EgbvuNy0xG53Ew11TJyHNrXFXOwviT/miXoAQBlWCpWq+HEbXy
2SaNTPcVCSPOOUyqm02iClO9hVs3IMHZifsmBE+ytjcNPj0v+ObIOCZLzM28GYM+EoBgpYpGKZhx
Iq37x7rK3PuIL4Ok/XdRk/dmsjV0m9AOSbGfl3OYrOYBcduYyQij5pjL7RX7Fnou25KKGGOIoRAm
ULvOwPFXznQBewwrfCp17XnNdWLtTcnUZ1gsX3kDGsWAld3fE8Z+tI+OlseTAhhHaIoNUMZ1XGNn
y068lqaglSi47Msx3KuwvzBWTgKNZkaUT63TNZsbipuvLZbxFORigX/tfMJcm/UbQ8sGJbEqz1se
ToYFktNzn77v1DZCk1x4AKVxEGWkBsk9gMVEuM4+WV2BDKEYRpDk41Y1zW0D1FgmCw2NsoQY0TDX
9QUIOfB1jd7RKspRiPJs/jJjwnJMOBVUhAlQprYG/gOWI+dA3oR1lDeBFYsoRT5ZN8VREohFhwuX
8moLeTWFJrIbw8I+tgDHjjRfUsHbgHoJ11zE968WbuBlpnYfYLUq8vvjJC61OV+w1VN3i5Q9fKjN
2HB95b1rFm426kvKjgxD7z5A/aqPBpFopKuKrYI0AUQBsdLZMG4lxo38lxqomaLbG/SHcwqV7X+/
LT5QeNocveE6+X+0wD7zPCsH2kQAbkv3GhLz2mrlVT5yMl8WuyB4ZcerZBJkhhkTDU72Hveae+2u
i4MRXZE/j6bfpABAcBieIdqjmtLxbcpDZvgfvHZ5UiwfRzei2lIQ5HshcT3vHGPi4eNK/o8rUOEI
RBZFhBi7/7LjlDFtYYFbHHTN0OrcR41kMfWK6kUWmzaH00cx4r92jyyS/qggF2RxRf6Zk7cSCRW3
Na/+DoCAFWVokZr1SLhtTeVvp1UR5ULgX4YEECLXJTpXGekn2F9ANp9jt+tcg/os0ZVxsKVMyEPL
vqDiFQe1YrTz56wCaqbhRzgoyw3i6aTzr6eRXqDZsbh3EFTnXYz4BRrR/3+OFV0yQ7Xa+de3HZhf
enGF6kJXaCpgWpJY/ywqAiFcIxS9yjXJqikzr2LuwvNAioKwXI2PSVLtz0vlAthFEW6Wjk/LmNyl
uqg01Q4oLqm+2zKHztbWwEOr19oMdtivSV8I4CLEwFCHkCxrH0+YKFSHoF4sJ/q7v/SdnNCwNoKd
1FI7zpMljBLD1ASALti4rRfo9IJBTK+Bkn1x2Al/z5THEyGIKGE/NRWaavShadRhxJLnFw2Fj3A7
+pj/0nfm+irD3acB3jcrQnR9iSHJLap4mhMoyMNSXVd5jz+I5qy5PB3ruxXeTyYrqf5H2tqoZUSv
iKywAcjVpAdruzEsZS0Pon/wKVrj8R60DqqvkOtlPSPeWqVBFyC7BPe3QNavsODNc7RktTp9m2PE
p/qKfhIbv4a2I2GjN9zeWdE8zvfXBgdy9f/IR1NSEcGzJ4uJkXVhTnCeHBQpTXhKKkcNbc++rejz
/aNYoOfIEMEtzTNobgPT/MUpuiRcHLrDC8ha2jK4KHGdpCScC9nTZb7lO4jypkChpT3F27RHoXjQ
wd9a4FIV+83ZKxQWmbJMg7GQ6+330GOOwbLIxauvIXmQxseaHmdGDg9fHG2wEslAhoGBQ6zeq+hd
V3K0/iVwUfg6ro9Oh5brySGpu6jlHyN0Egg5nKrMeb67PJTPeWNzp0gk2ZWwlTxyouEwRShGwaW7
+NoYsuqr4K+o9ICJ8vtXNzZJ+JcsRIrN1jvrwbTyJvSt65R4XRpEDNiDSbLzs/0XeHKrLahtVYEk
WGXj4Znw+GD+C1mdlrN2ZjQb1UWui0A3NiPBNlHMSSmzyEH3JANbFRlPzU2aKjsKfooTtRxKLCod
J8fxa4fZledA8qlnI2shLLWN0euqyWdz4BpJkNbBDVSy7jNwDVuPoyo6IUnYnIX5PPpAWqhqizq/
hiRlcchC5aEJN1t52msJ/Wvs1u62N2UPAEtKh73ewJsGcxdoEDeM9aB2x6v61OyKve75Zf6DLOCe
4dTT0Y4BNXymSU97BMCh9YI/xeDY9e2ewXZ5b2thruXzg+SIVdlFGkCT2+dsB+PPYoAAIQ0nHYoW
4mHiE9K+NFsjMfzwfbbGCzshjREY1/3r/x5XtBcOvmIO9zYUdq6NQrb2YElvlTjU/Es6XzPlopT5
Qi+RyAY9xy3wM1JRipMyXqWtAQvzHDc6UDPzeTE9lDu4mKXA1OwIlqSpCoL3vLOqi7UwkvYJDZgh
Mp94nxGNT/fQE3TLfCTSAOdMVFjtfaMAD0+2hbo2JA12gP82EzqynUowqSEV2DR+aEWelkbjr7Zp
rj89SQYSZo2zYqrz24K2TdNtEsKKdfwzjZc0FJvaR+kuv/FUN3Qxdm+AoJxCwm7sYB72n7ZT06Go
MFETEiuERu8UUJetmb/Z+6HwQVR2goy5DRyRDzuFGXKbOA7uIXpKQk7P0Z5wd3hZumBraACamwKz
Wpuk3r7ayqNVMDtOStRcBFzeQNJi9yM0dCWCoUG6u3eLtmGAew1mZSzNPEdzAbHoyMHYiqhgDnWU
6cCt+Wbk9FQe8tZB9QQXC3V2s7yRCbOgHEQCtiw1Bang1jPAAOeHrBfvDtQp0Dmg6M+IAr5U1xjr
Yon4evUyKWE4+NG4Tyhte1ZqNLImmcpvxeLezJl4CGwja6gRBvKan4VrghAtYQZAoJMFYwCStl+u
qUMkHAXthOqOhuILLij3dmR44o52DKWx8koV/GzYd7I2KiXx+cy8+4Lezu38Rp9Dbk6FgpHlGJma
u7sacGGRVE+32CpMCJW6ONkASP4IdRYkBLRtaT7msjK0uogIAf4ZgGdxPUEVuhk4GVe+WfkTjHZk
QAnYUwqY10RvSfGUBsfd8WPxvnD8dzrqA4pSaQm2zrha2IOgWR8zYRaJUlvxxeqB6e9OkExQSHY8
Nbye5dYtjQW9BYVWh+cstfI67mWVhTusMTngb0wpIOR05mO6zCQV/g9GWCJJbXm47xXuv4sFkMD7
WotgP5C1ygKRzldCLKsGmliReInupTeheHba/PVF1WBW5UjiIUuX04A2pLH49k+X9FbM2/ogFWn3
P/s5obdKwoIdi98urzgbWP6VTbiT0NN90eaLnZid5u1Dom7LCbIe07QtVPyZUPBKjmkYqvygVL5B
KQTWv+BgSWkfL5A7Uq2m+hYpUG9mLn+tAaqVVYLvIgPYuxxaTJ721eTUAD8AOEWd9KXih8HPYrJq
LUVs9rKXmeov4cB9x1lwkZD8T1fMdl/i2+1O4JguepslLig2mV9Jp0di6a/EXyFkR5CcTk5Wgheh
uZQUp+VdiM2HfOAmhaKMoc9r7fyHUJz66Gp6OMWCzhFHWPngv4DTxhRnaXwCrWd0z7yy7ej7BBha
FsR2eYsAiWZ5LSH/zmjU1veVUoeUtJKGuJYORyKfx9OdiRK29tI9tY5k3TH1BFgnB58XtJ5qMdHA
cmPX93KnL5c7aIUX02p1SxEuC4qRzp1a7LCYbziAc5Sgaweax+FM1q4LUyeqBYb+2DdbVHiO+OBG
DvvZJOzy9pEu649k8fhwZu64Yon2OH5w5EevFLEum9L+aMjBkBrzvv0KhkkIxWwgyjk54bJPTYJj
FVq2l/ISZMjoRm7AIhrtt32FDJ6tdHsb2aq+t+1XFjfS+AM4pKy+lCVOYwT8H+s+U3QaIn4tmEKd
CA/Xwbbn2gf9aZHfART0GhMP1arrzdN9IJ+Oe/YQlHulV8lvFRbFMoLSECOaAilltxpBgVBey7RM
8DfwsaKYiFCsr+4xtOLhUSW/y1Sa5TTtJPGt8LeG3bULCJOHuLkroWrDR4M8RyoUsxgygpXFsaAQ
qn1iW/KVTPTcGIj8/cVJ8JJ0EKghyx0h7NY35O7gsiD8cd9Y9y/Oy/Htj9LsCB8iJ6tXeOZOTYX2
/3qiUzfgFEsjupe/TTIyz54y+wiWUVL2ghtLIdiUgK9Oyq3+lez1ADMXCdgWdCh9LKettXmXnhQN
OH4s066M40LKC6OTwR8lZBxt7ycEesPJ5chpAKJQ9ZuUy7WqFDV6q1JgzYBSnvRw608PvInao5py
ukMjPVJDjQI/h/KLaTzGuSFWN3HAFESTQZXHgqG7AMLZBxi0vgjZk6u1QqtRy8KktZDcsJk3jl7a
IZV1CmCS8dumhUnZayGH0WkwI4N989CDLTIg02BqqHtACYreBX3IL98XD+m+LxGqnT2LvP+8+JcJ
wHse2UVPXGRENTLZbIRjrfMqhcwzgetBS1Tutsb121QmWaepYopZ+iSOaV5i9ibafdoxiQ41mQOA
n0sCPzysDF4T620EKsnR2dBeLdeUabMKQJriHAtNgvjoIyPmtNSqHGu+5K/PkvyGA9t+efPeevmz
xtWbtA4ER9bCYRN71iF27YfQamriMfJiEljG8XLxXTx4Hm5cLbtpz9gJxuJ4tJ3UwU9/A6Gn3oK4
OTYv9TXyUP8t6v124bkiHFtj70vQS451UNEYEGVc/ujKOrSpehIYWbI/9kLzGNaghXUO/Nd38fbq
k8p0zEko7gLVr2byfzP7ABXQH2np7EiUeiC5XbounYSP3acVM3iwXxzdqhaeN9fR8gQK3WeStIKZ
66j1P5Q8+uvxz5pwWFlgoW2WK8mxK+IQV+KIwf6PW4Wgk9InysZGC75zTdB5AV5DxP9Qene7Nhcd
0qg71Zx/QlaNRyS3DslgFIYdnYx/DmQ1o8hp+2wkhFIWM6AcQkivrx93e6k98DGbgKNQZjm9/mQL
AO5SscdCg/ApcY2otuTLcbGcRe9lVu0zLbw+YuHwM/4I5EwttVPU+byZBgDUapQf11SiLzXQi6ML
HsdSj79IlszyLxl8KJugYzq7UCvxyVOaey+vZApYesoHRyE/D17I7bIyoA9FNwgRI3dwhtA7Qc0J
hgF/Wjt2pTjGmoI1M39l3/9JbhL0NiKvIOSin/qybJP1ynmACsRvOEAfFeb8tEy2zKk1Ch+nTEQG
UC+3orLa6tkmuoU4jPjkoPVYyXozUkgihSmc4Klo3hN1yyytssRDkJUUiQjZs+b1s9b5LO5rxoNg
83yurFp0doux3uVs5KUED8n2AbYxCAipSdJRQLQAY7xLchIfhSHhhoQGcDdVdxhFvHsVbSLHe1J+
Y52JHzBe0fnTMGUH57qNbZB86WsdzYt+TN99iwjwsWu22YHTzpM4t92qvEfKRhPC450GKfZ3xQyM
jEkkWkcwZWiG0q+2F6K/LSYC3p6BOf8S7u90rD5El+wkK1IV6T31HIKdA93XUDs6X+o/+fy3hMDe
lxxJ0jCt2nMnygQgkmgGPaYABp6cIKOkI5iyCEkfJAmeq/U1zYluXl7pT8Ab327tf8YJFg29ymDU
tzp3N2xtWNaxq24O+i++DE+jXP3AAX8pLF8eUb6uD1zeI3ZGV1URSRyzjRR6VlP2QtP8DZ6Ewmdv
yPFdqiVoZhVkb/62q1z5TxdartQkfTRxtb8v/c/qfzxpOMdLF1JSykAH8qbe+thK1mY112c7+xmz
JE95JHoBvvZ8Yntg5XBCI5RoSkIXgCgntKdi20rBW00tK7teWwnamp/4B+A/zFHxXqm2N6ABH4kl
qe+nbmYNam8ou7A1MXavTVszhMPgsWkMOCuGqr3rMjOcE5hQ4wqcd5RKaMXGXRDRw4HS+p3fLskN
OPNiqJE1HbEfEa5RXRyFnZS/kbPeEbyd3jMSOLwbmL8GW4wEdlSsUAAmrSTLzU27TH5UeuZQSpUU
atxsqJet2RNFg1SldiLKrQ4/wtMixXl3GHTNaw65hj7ekstdH4Sd0Z1Q5Z/ArerwdVWojrMQP04w
aOJFsO1Fc7Y61Hbai9G03Q0ccXk8HzxUnjU7jJv22jLZl/5lXHmO0L5QN2OZv5HveO8rBShZTo8m
ohsc263cfFDCUsLrM+zCtvzvSTDYVY3vZERZzgivt8wbFh1SOd+WHZbTKH4MwhJZTv0VPuF+Oo/Z
vlh/pRHJV8x3obQ+QpDO82BH436jnGNrEIb93CJDdrHcJBK/3A5KpSrckcWUXoq9gftly9J66fEB
3iU5o0VwqpeoMyxMTMojWJhCF4wnkK60MLzmLSqAVMMA9DH5+LTBFkH47g+H6dEphkjcDwpX0U2C
mdoNOl1lzbk9VOv+sMnsLsbCEp+CEmWtKlrZtfesUrcL+qYNIERLAdyv2oKfJcmMemBXcG5/Y8YD
NY6BaaqcunR7bVyh1uUgHjzAUNdatqtDC9w8NdO1dIWPWnm6wGBVwTZzqGJp19DpX8lMq39bfPpT
ZJCTm05e5e0EdlfPTBQxs7LclZMh72jjUQ0Gy76KqlDwQZMsqjFX3NDTUGesUbJayRdMJpYL2pL5
LmWGMixZ6L7MqOU/ZIii7kop83+BdvJKFgTtt96R4kKnjsQp8BCOOT9PeSmSDJAtefZ9l9qheICG
hhkzgOIgUh4Ukw7GcqZaVSHsWJjL58n2oz7IZYDcJbtGTGhT4cc9YtNf342Up9GpVkq34QV51wlx
JuO6jRZ4E/BLpmFsnpqqLzqIZYPyZJ46JvFg5oGs8GD8I7pc+Vwz5nxXJyAwCsBHed3xirTVytPz
zg7txrz8/qY12ziFXgR4Mz4u8b22nEA+TrK0sslY41vJZLpGURaNoRHaW+xTFWYqL+77SlBgY33O
nz3NChrThtN4Ll/HpL/ZYdcW5Amjsd4dpx8lQdokEx2u533M/fWBD73xjJ6OA7Ou+WZWEqHOe05U
TcAlEB4Nt6oP8tbi5pWds4zlYLrH78SGLvahvNuJGpseuG4lQT0njWEqRYgohJ8fAFWZJIBk1UQ+
drj+o9wuY58j0Y6mPMJB6vK7AP8d4cxvScul9M/ONYaO1/N8zgOan0SHm5JbS/U/6iK9O5+iaxPl
xrh/6X5gfL9KaGQkqc0GNcQJwvdnYs1l+7BosECQIUnd9Gowbexsu6SKm1w1a4ivViCJPti6NZ57
cEXwEvyqPYERIHSBRGBWWQqJBajr5euts1nihAPSGT0POhHDhxB3R6kxCI1DVkinnq7JlpL4DT4e
KoTdQ7K0Hi8YHwtgtFi6C7EMza1ndt7aNjOetz8dI3kouQhB/IDsfD1Eg4A9WKn071lL4XoBpOHL
j40wZRgsv3it55N9H5y0zXMFIx6JeGpDJwhbGxU5cc+jjJtwtK36JRZJPqZdzGXjUMvWM5Ha0L5D
WOsx89hTvhe2WrnXrnqHKGHYhQAwj6wq18LnYuLPsDCISBiZ38H6CPw2cKrDbBi3TutE66mZpEi3
yhc+UCp1u0tSADpPDpHE2uSoX/JAON+GmhRyt4JLj+MiYLCGOFqXCHUmPQuaGrFbnAHJEtKyHQ9M
ksvfw/crvofsxiRvcvPeiyt5MbVeRaMxduXl+kB5DvXu9r/D2EeyBkuuHHRbTV89aRAOwfWQyR2k
IHkMkeHq8uM1BNPB/CBNcI8Sedg8hrGi6c+CScvGoWe/VhVwmOqDzheEgIqpQcSx7dDqsBebPtWr
7/sTT6m3YcBoLfhm5ajcc+3/j9eY4gnfPkJLB09fLRSWlKtBYXMW8a4fZU6qxE28GDrklUpxeD2j
DCPRjJhlAPvlttpFxREGe8fb+esHXaDPWF5/ZmjS7xQVA5jwiYVVQDdSF6noueMN3ggopw7mcKd5
CW8GD8Bnq3O4eTQN9xkSuFPe6mN717aZHVfvtC+awiIC3jZFLX+1s6yZDN90LvoidMifzNOKoGxQ
esIdZF7wYwnatN+KpHiedqZVRSQ52u15YOq9LRpkyXQTikJaRxNXhDIu84GJxoE+385ebTR3LBti
oJ59hmG7RXxqhc0ZxX9V1ZJi/hUi4fT5+5pUuz1AZ0pLDcYfP85FD3J7t4bcMS4GL4WK4uwhjKvc
m1DLl2Ddto+JzUYEsfpH6aca1bIHA+mi40KWVcv9w3H4tHgjGvCRy5g5ZGHO9OFF5a0C+THDs2eM
saEvSmB39HqovcNEanR4wmzsi/PQ9ezrrLqOaCSDM660HcSeCrKA2U6HD3Y63CJVFB4X/n/2YIq6
ObTVFjorCevpedcAzQVeXoIRU3N5etNTuyuggZVUtda5rbp3rYBR/uBMtgqia3E6r2kyd82X7JGk
E9GpLjDoRunyDz8DZq9ewz+O+dLEdDFYy5yU3JcE7p4Wf8VEEwOb98ZDMjfDMJhZwHi+rTHGr6u7
8SeKNXOy/QYGBQd84vcvDPvuau6x4OqYRvaiUVE18SPzyWjcGJ7i7ALg0eFrhlU6O7YO9xl1pKTU
Ac9qmuuaaama1mDhDnhoTDJRkwbRmFZVrCfh9LLn2YNqc+OCsUpbfr4YAGa3cCl0FDMvN/7N8WVM
5ybDdGSTM85vM/zS2CYB9V4D9v0uAsDjQHaMjDGzC4WFp9LdKVGkT0fUEPn7kZTtGBsvFtw2zDGk
lX7tSj7qVYjaG7Bmady+SlPAFJFRc/kntSX7ju3JPEXxyiiomcE/VE0J7fAaosb61Pi3DOHlH4QH
G3Zz42WHMjGZtTtZILiHTnwVc0KjQY8ap6tQufNX8XdudXDqvEJEPfx5GTWJJxd0KGiZdZyKl1L8
ug0J81P0Y0qHbyQPs2lAVGfjDNz13VXIfPf/OPVvvDtpdJdpWIJEEva5nNEAmf3+COMMxDoMpZzg
zmAmJupOG9UP5lBmJK+aZJQi3Rmy4j7ea6m3Y21/r4ZNheZ2YnvxYOOZDCMCRCwqmChujgirjOFL
3NS4IppG5zvuHQxJPgww0dPqJiq5A2/JrLWxaPwFgDU0bjIAgXmGLS59aRjSj/mSoW7/cHBCw23X
GcUzRUcIW2ILBRHoqUGr4F71f3kQq0Hb1QdE9mC3pS5A6bRiF/rZVubsXCMpb9lIMz0UeqgXx42B
zTruLpSuAJH8i/lf2txHVi69DQs+ARx9E5uxpb7/4vTSl4walb/6eBhxkuz2EyhYVttGr1E8YjD1
dBbKtFJM/yoYEqbRUVcVeqPsNpMO2YvzOFGKVeSpD4cY/TfV3EGPzwrd37GFID0wjcElhQti3iqk
1ivJPKRzrvFn72e8QE04cWwQ2UTFZCybOSw9WQwai7m0wro6WN5YXlsB2cWdKn5IPGBI9iCB04gG
8jOt7QhvvzdaQ6oHVBoWleCcL0de9pljH004J0m4BDK+i3zkmtnTS+KOjaEvVMQoPhINpJrtQo6I
7TipzTV5clOD4TtY6nyg6WJcl0BCk6zlicQ3LzEBIQB0dY/UvQ2SJ87wcyTnZ3OassxEL5sKO5EX
HT9mZpHUY9G7/HSLAsDyIQ2/W5pWHVj7Bh6LHKKLchyHRULlzae6VY3Kx4vjWOOG5fDCo00Go1sl
iyfmvTlc0yTSjP5bCcf5GTs61011uS3y8q3X+XifqSDF/87nHelChRXLH9RrUkqtnT2dvu/v6Ac7
aoqmMA/7aldukYoX3iOoMcM6IA0yiEPpmbA3N6FzV7zO81TLYQ3VLtsIJbs3hcW2Jm5XW+6wL6hp
VEA8dKTEGe+Gu4xqMcZoC79eRtVd3gtYAGGQoIfp4/7QAI5WqXgdADozss5k+8kvwY8Bsmtv6kaV
CPjKlFI1M/PS6v/dRN88CWactoQcx2Kl3F1mXVa/KeL//vxp6LJwLbB3ezjDL3wni+P0y8ehYH8Y
vhoiflnnc2sqKyp8yMcfAlKTRdvkwxnLihjXc/7oiBWJ/VrKeUXTdQUYyrAX3b8ZByB0T2kukfnm
HBceKq+XRFmo7mKJLyRTXbLEBI2ZcJMnouVY7A+HQdYNDgD/2/2My7ANQtX9fAY03Cy3W46fCK7+
P0GX76e5L98TYKJuP7DrlTpnoHTuxs2V6nve3YxyIsoJuoYQOynHMP92+PbN+9JgJwFGYTLeQ8o9
gtqpADRm54TW2CW6xB+AAfjJNd/vHkFRYTHw6uLqQ3Y2+S9uDhuZF75hh+NGCC2UGr1CvU+8Boq9
DCEOfkCZzYGNOLcKD4+MkSyMLHR2G5+vtYVcFjY70D2yGzaMahryqK3q6QjoM/kPBZVT2L+sWmnF
tLtRRwWa0i360sxUUOYfSi9ofxsfZTLh6qidHgNjqI9cuWUgbr9DDV5jA1gAY5ah68u//Wl7k0pr
kjuuudjfQvZvn/UM599pUTKp6qRlQjW9oAo65BZxpSCv/jlqNiR/zQTdnuxgpKcaROBdt5O6kQf6
bwRR5RYotuu2h6HUMEvRhQCLkMSMTc0Rqx9/9gBkhZYk0FIHXwCmN825rq46hfYyscKewiITxmkC
tQGEHwcwSVRu164+QTc6A/M4bso5AlEmN8Sj+GZtJFip4mpHLpL2CPlEoIu+Z1pT+i/LJFO8T3IX
OFxkkrgJagsk+EOL8RU+6yF1y/PMYbPcIuti+snnnk2y/JTorpoB+LnHqFv9+JOx9gKLdDpN1SYD
tHY1L1pAd3JVxod/wll7eTtUN6+BBcb7lcf2bMoLZm6Su8tBALr2O2lafJ4TvxUhtYruQ0ySA67I
sCyta+uBgR1srfCKnDxdBRZJzGw8cBuXXMqmZgS/HpzuYSuXAcQ49krun63vAXGv0klR4oHPe+Vo
5+qhZqZyRvbBP4g76A1GdA1ueYiyT1lQF+f3muExznOMpZoSBwSKB57GZM7sT6cLQczTdIL2F65Y
314D8a/8EemccXiL4q90QmUny8aYmoirrhjLFHAoD07669oiL0zwaHMLbyrdHUO2HIzWLMdngr9P
1uKRWfx6qcX09Gx4NANpszAY0AWEtbiKQuJbjHu3cgXHtRWpVt3rwfCQWFyE3DH0tz9Zpg+Pa91u
Lf1ItTAYoXGuMZ4PnHJJTK9W+vWNLG+RHMphYviJHYzdZy99TVA4zJDHryEiOp9SiC6qc32M9yIf
wxkOCDQ+ezG1wW81Rr1byCTAq2gQLlPozysUpnHVn4yqJNbArLU=
`protect end_protected
