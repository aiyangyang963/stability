-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
q63D+ddsGrq1oCGumt6/FyVaQQSd9V2K+Cnpv5doK0ew9GoPw0ywZc28xBnA/sbZ7PKA+mwfKyN0
51119WkH8+0P53P4nrRaBkMOD+k+DwnUs9L5K7lYdQB6qJ3vdOmeKedbflD3is9UeOZW9TD3fnVO
O7Z3Eq9dlg8mZtCEDnS6G71EZSUga9l9dASumio43QI/fXF9XsXTwvyiDlohlxl2e6mNzaLdGXxE
GdrQdpMHLlHg0JFa0/G5Gz7RK7/l5i6Jrn/78L6RtVbNC17Q99rezsru3owyjJ93dXbPxrt0mJCr
x7ouTHMpQckC3ZFMNxFSt46dQ1t892nmBGS6Bg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
KCD1HTcByH2AqAiC13L8dbtFVZgQtLCblLsDj8jRjyNjRRI9cRjQhvB4o1any1j1vSWqDrcnGeXk
tPGqImIwRuZtueqynjatNyLVZFNMau8Semsc6/TCkmXezZIBo7KUSiP5Fi5FKKtR3BGAsvb+g5ao
XMIvHfIhT6piRUtyUafZ1FlsCgGBaJ8oXwygfrkyjfFsEG8un/HwiyzlecaoRssmsbtEEIbhNFFW
b8ad6l1ALSwduckXLtgm3oPzlrQbd+ghwmRsCI6gFb+GC5Jj7lV8nySMT9rNlmhDdynLmPPvBQs3
zNljzYNZA6Y3VY3b9yZtQJ62MzapCsB8lhGQMFPMKIy/6aohbk6GvACn1Ah4nJz54ZLPIsEIY76M
74UEFlrBZDACOw8Eo99S8/IR6tdmG9nZpcqU33J6uyWrLgGUCaeS28SeyvWCYG/Oh5SzhELd+SYp
RbFvIgIL+QJNbh/Kfi34DKx0TtWPKFhVf59uOmWaF/lBStf0grCczfVf4ZCQn13zk3G2i+GQU08z
AvDK/AwiBf6gjrriUR8/cMN5+zHgZ5ncw3HqvNswPBVUjFuAU0ViR01Du3+arIjs32D2DuEHlWcr
oosyFnHD7F1IuagE6SFY1UaZ8aSPkcqV+YUyx7rz3bHoT90S+w04NWFqG6EiPhF6Rw29YXRXr/ju
4ObIzkSdBWtap8tkGyWeXfF1fOmUH8B9TtpXhln+xwRWBT63+L+PAJ/wDGd349Qw1dfMRGd0cNw0
xmAT2xV0gNCvkrAEPv6/QeyIe3x7xR/buHha2xAs67CxafNynElAVC6Tcv0IP65W1h2wgoO5cMPI
wSA+h+EcQozaKY1yUynIf9E0J5ot70IdVwgTXrkFH2Eooo/tEXeHmuHsFbhGgcAvI0ow2GoWbULv
/1nrfSOkWLF0AjL73y7XGP/bvnDFpolkILKdNqxJrmHcPL4veDsYNMxegINmBGgVFG04cqrtW1CN
AMJ2qWJwz/Ip/rxYY2T3E6uVPTiLL9e1e7vsJ0tcGT3dIB5qllk15v+NPrIpZ8MM2gLz5NtOU4BR
gv0TCS1Xcu0qAE7m/aeLXplQ0kDwOSVamyyHJG4axWMtxnoJy8hq6TA56w/xcS7BUljrW0jBCmn5
TMjtwczc6PTff5sXzLXfu0xdSJ/+Xp5hgUBGqH3RHJwYoT+HA/A/Lzv/mRvWJFsPlO/IS4LYCLQr
GGqZzQYYi33KbrsqGmr6CNucTarauWQ4cqHt0Mzdc6tlmtCn354VXDmu+Pm0lXwkpWxAe+W0ua+y
6nFmRdLd48k83TZzBRQuMHufYSafe6Z801z6zZHUk6+YUGoHRaEgsEexbgim+ueT6Aclk8i847QV
FPrJ3louka0kXxNYMTB7+kBOl6FjI2N9KXJkQUUw4uVjVnv+G1xt5J8pi5/M3Uy7DvizzMLN1QWg
ZZIKJJNiDOy1rymYV+0DqbfLTmZZbebruKnCHaO9qoc5CfG7HwvOFxWQmRSdQHfQK9EmEHkn0FeD
v+jv80X4ELwRURE75BVP36RlRJyEWsJTcqiw3DWH1zKbZ4gcoA5vI0UeZjh0BeUvb71ccfiqaE4V
lZn8HXjvkTwsPWkrVS3clyIF1mdYGhvFQnlYWjeIdXFHHAPOZzQ2ah7vAPrIPbd0BMhxpw7UBGB/
BdkB+8UV51Br3EjmkCwWV3vbmTN5a0REIrbTy3N7ibjQFYonyQ8Wka5nt1akOAJAM72tQ9EDTqSU
vXxZ2ILqQAXinZ0Y2uLywnKTYvMqtBsWdR/O78U3B3DnMmfU1zTIUJ9awRucQ1pp9Yg6aCs/BNt8
lfiq4mdtsoCbt+M8AbU2UBlg2a800UzaHLjmAI8mCWA5dSxitsegwHoAdyvtxFkV8F8tlwTXSrlE
aH852hgMq8uOzFehjhriWLQTbuhuuY3ZFFCnPc0110pRwIusr/CKqKqaeSE3zbppbzptVSMEhCdy
KhOQLmG6WYsQRi2+FZKtIdaK6DRLsdvjqML5Gv13uaw9gVhAKVk8kJjx5YfOutLo+qxl/JFhu1Gj
hFoRYZGoh/zr39YSVUWigB0isf6I89N82gwcWKjWPNrIKyhHJ8ONQDA4xU5ISbSCazcpkdowv7Wv
6R4DOv4W2n8cvxuMan5ISLTTEEEeccCjW80kqq4/YW9hrIks+ZZorfYfJWrbb9Nkk1ztQKq9F/54
6heJGfdqFE8NJJEgfbNIYuIkgCaovrGumGmES5FaShUEN4zm/E6GUStaaK7fjZmuWNq3ck3Cy+MQ
oi4+PesM/dnMVgf+D5lnteP49c0y//rBKDcLR603opI5vpqAa+7zwcDy5B7zjiqIVapuxjjBka01
6LAWPufJB0GCRRQgb14sW6prrcB4aibtXJYbNzw7eRsV5twcHYhCkmu8QUwyNhMjGJzzwlF1FHu9
Hgg0UA57ACGYtLLrZzkvJfabo04nFQ3ylX3WYvDL8VuJTIF3PUKODSKgjr4IGwupQJZGaYYSyOW3
ZpslXvvikfWA9vqu/g16sYrE4SbkRwJEtBnE0i2AGjj42AR14KC1Fk1jvys5Tz77P23ifIfx8a36
ctK9WizpD8npO+hxGHPS0ntDyqYkNPW+nEMSa3wL/8ig9MRSuIC99bhDAj012n0IOHXeLxv6UhA8
ENXyDF8wOESkj33th+kK5IDBAbuMA/r0Hb6nwAI0vOm/yxHlrcYC2F+XOsmwdzqXaxMgyuC/TuUx
DZ4BheRt3EXY72RqUAlEp0hIBzi8Y1rDeSztMFZgxeXc63XhSTVpeiPobJRzL2ANTZ3aDaHRUBQ0
9A4xw7q7xOqvB0xt0eg04tjuqADnPeKz0jfvQsE1dM8mKRTHgF5aoWb19ZdR6xw0MbEQ/NIuConq
1A9vLdT5X3PsIaJcRK6ffq31l0Vb0F7FnH6P+C5LUJIf5A3p9dFZHwpNkuP903OjowRy5ibzUUfA
ZezN+4KxQ8+4Vgvn+2RK8xL1rYZsK2va5nA6hdC6L+2vGXcax/xsUs6C0TC3USYaJINrtp6y7W75
7/XnH0kPqInyLeSVvaQRyL8xtpn/rqkdD19hOg9E7FRdeKk9RzMXirhs2M9oc0aTMqhXJ+RVemJk
JBDHHzwGocUCmc4AIy+xbtHcjrSHNS1bLyv/FplOUicVnt7pPBHYkyRNpbFaUB1X/RJGPWPomb2j
WSt1N3j2c5CPoaXYtlWwDB3t48d+gPovhE2/y3EhE74DCe2tt4vwmGhFJvIPFq8z3WjUMsbHvSd7
rgoBSRCJaf3cr35cQJFbfzagX8qSDdXxLSVvZUusZYptadQ126Am1SA9HbfLpm5n1YQo4sW7xdPE
W1z9oKQkvfM2x5z8kpQVj4nsVU+50PynlOVV7RlQwRXR8S95Fw/1s06E//fMQgkjO+nGm1QMIq+/
rz+Kz7RRMiGWfe1JBKkMfa4rpH4iGJnAV9n4XvViKQ2SsOj6GObjfs4tH6ehTEvKsABDxBoP29Fd
dzcPmCOj3jGwND0FIOmCRRthl9AryU1D29dUjE8/pXw7C4gGAQHmmlCKh3PuKfjJ5BwiT8x832ZZ
sAU3jAtPRuUYeqigvjevGJjRcUiln0eR851AW5vwJAiDN7kvAECefXuFTbYTjz3sb0VG/izelkfo
fhWORj10aR29dIcsids5AfB6UPy4r7yMlyM9i/FF205ONdRLT9hpmafTGWORzO5B5H+B5/7yel7l
KNg+QbYSB3rJILfQ1l63aX8NSLFv9wfVjNfJJVs+X0Bs/mOJPkKl1axgCoimnOKHroZza6EUTlmI
NEvyBiddj0Sgt1P/aT47HXrRmeyQsr7ROaqesu3kU7ZwFhzw44/5O1arL+J9pdddayplcp7kkRuz
B/MYTn7SlxVx05P1RWqpOgyrEknV653bn/FlgyAhKqZD0sufcyDgc9uzURDVdCeJz3lxs15Wx78O
oHcM0i5L0eLAKpHbqE4iYUANeqUqs8HW60rMWCf7/tksgZ4e+SR5zh+axsJrR+TzRtv3OKiAvPhs
W7Xut9gY1WFqyfnelCRwTfupfTPjISdcQeJUuC77EPP1R++/ecGd3he5i+d7NjmSY/g9608FC32f
iwhtY6Wj0g7dAL+UeU/t3SyPNokGkYxZbPSq0yzwsIqApu11Kr4w8QeDmT6XMTTxj2AdpIpZmgoQ
etr+zSQyC8zXGAVgFQbPivd32SIDWu2AaqKPderv0MrF0pTW1C4IglcoJeRLL2paOy5LXUXEFqsh
2TYJwVgY4Vc+lZmehlOWu6fRn5URt8QT06+wA1FeOsbyl8d1MbqgbU2xVLhEmEV5RO0WRDlsMfcW
1U46qvxh9zf9rlX1BQytD9SAInBxKuaP7jgqRcEPJi/6azApmqgLmSnbcQtruO4qRG0Dp6IZ+wGl
XuTcvJr5lk0vbCe5pUrjHAaqvRIWhyjYdEMbn0WCSM/JQEjU+6XegPe+qscu8pPtyFzIbwcELfMR
1p3XeT41duouLlttco7AMjH73T6MuzkD3GK8yDx1mX+UkPzbtHcDYFp+gxsYu+swI1mnKj2hu1bl
vJdaP1NEqeqtuV8u7XdfhR45thX5rZA79+f+sMPVELd66/gUzWiFISPqC/sRyzmZRDmanWmVVnIj
z+LcssUw2Ipcb1w8YBOtjqN2/gKMd+IE2gAXkPvd6KEBcku3mMg1eV4ugjsGhSPovrI2O8HMv4J7
OIFMlkkD42JHVe6erJgJQT1fjTWSOiSd8//Is+Z4iSUdbGZzawwX50jh+F8FHEN2MuKdw/M3ev1e
vmiMpsdI4T5qX4pZT8Y695DixzKyd537GN/OyLglBo0UTZHuJdud4Rp4NcKVzS28u1ViSfY2WJer
boiT28SinqKTst5OPO72RYadDV2jsgtEcEYc6QQtHL6mmjCkFFZxVniImMWxtx8z0TQXM6KZwtmU
gun9voCcJbfYpLId4al7yXvmDtI4MaYPNgtX0SwKbH0A7WdbVvnIvYpcJO3m4T7+GZSxLni3QfNA
48XbmnwLj321VdTs2i2Tg9Za6F7C84+PHdJkPoaD6hEpE8AaCcoKVlj5VeSTOvg3AZmt0s37Aoat
tA7nzfftVK50F3dtekXo6EQL6xQNORp8hQtxpO97BvSc+dsQn6hbA5KrbxxNtrOHkNnrm8wuoZ4F
zA50+xxVbCORuyzclc9VV6DzctIa814HTW1z0vpgJG7TokykCuSXxhjnF+72xuNqjC62Dv0Gagqb
h0YOCtEwZAiKUqJBIguZ3MHJ/ZHX+L6zHQ6bcNVzfxzssmj9rOBxlcqaV/p0a5N/XJa+QVYVV/Hu
iLhefUNi9JmMSR8mToGk6byTuP1nQb3+xKPadV9eVqeEhXTgYJgFeX+8CKlh/juFy16ArFiyFVKQ
trXyHiJ/MRmswvI3q6BSngkj1skGBC31NlxcYset7ABIfImqsy7tG8Q6XmDXkRqMcw6e9ftH+/5a
4h7xw7Aw/4O8Ls1olqAp/xSNoFZwxr+B6LfePvg7S7J5vOp0lxO+d8xMzaadtsZzDPd5MOGNzvp3
TD5l9XbyHcX70kw954EC8Y3o8ZWxY+bV3rYMZ17OzMX689vzNueg8ekdS86CBZmOoJzlJf9j7eXp
zUJWR1jj0kGMHChlqyHcfn6Kl2GVgE2RMW2iKG2b3ruguNgyV3N3lRLnSwqh2QrMCqHMbmaBp838
rAMcj+y55at8dfX1u1BSSf7DYzKv2Bzfirmj32pTnChOw65B/948SghzP91ypGS2qXVTG60Q3U2U
PoyELUWYJGi5GGwXvhzM0Bg+e+ZtP2Q7D/uyPJXcELt7fMrg/aQhsR2kAgR/MfGbilyKzRa+jUH3
l4pnevEhutwI/UIOkA95MCzJd1Hpb03LEXWyuX2Xcwq1aSnYUt23u2ozCGqq6XUpewPhpEiLSIC4
QMLMLK8p6YwWlIT8E+hIy3Z6oqInh1VCu4b5JCYiQlMlK/tE+a2cyEaDi2GUAeq6n0NCxNMtLg7w
KFBnfMUS9JZz/T4qavflHKIDemwyHMAyfwtveeECrzi+p1O5Q9gh+MyHKxDqiWU27DxPVAhJqcs5
6UVcn3oc9lbVg24PipsV2KcteYgWHPus9abnkhaRNNM2axXjKRf0N0NyzFigO/g5Fr4KGiyggJ+D
/HlHqffx8YkQyBogWUoz3nCUl7R/rZXLx+FgJ/pqz5D0aPxp/+9XXRs4yT7lZKZxHghFFGqvrPM6
8yRbAvjci7YS48l6zHnlv0OF4jcKkLO/4TAKTjAfp+z3o8CEH+rPGqYP8OF0ifZ2Rv/cLl5Ipe7S
UIjwpfuFZ0JuN24a5CP1qPROSwycw+HM0hR5qifX6kGp6eL90AFIdGia2JkzOGDx6IR5KXcVsAWN
ufUsZy08zY951OCGCWreHW/YhIT02a4duqO6RyxQaOCQK63Vyl3889/HIMB6D4UYd3zulKF448fN
Q0L5k3NPKNPj30C+AsIIc+okGtTKSsj2OE2hUkciN+LNit3l6LW0le3A49Qy8Kob19Ja10dJQ3rT
NWli9exiR6D2oEGIVY9cvmIyouUV66YiEMDT3JOKr0H+RcW+qJyeFwUfIYmxnTpOkcg24Uf1tJwJ
TD/Zm6MauTpxFqiVnCor3ktUTbAEdEuHqhZ1RpV93gbj6t/ZLZuz3xj/7H8EAfyCiHXOh6kyOa7j
/kr/rjs6q3VcdyR0T8kJW8TiDcrep/74VSEDa/+DDCfz55WO/1LHlQX/+LmARrM7S1ga6kRxu957
gWwIxmGNnHgvkCZI2P0FVBQMoXgKu+gpm+DkqPz34K8pUxTfrI0ii2jBsZ1aW3vaxvoxBajXU0Mk
V/7/rJNBfaSPn99fJ4S4YCkqNP3Kyjl6o4UEJxp1MUdXFoC22FRsnKsEC1QzqEmkkPPUZ/q8rEHg
5dpftePkfsCB+EwluXlLl7vyfZ644fUGt4ZFMseHc9HnJYVSrLPG1bW8/YqBHNEf36sc6DuU+Y+V
MAvFbTADj/kEi0aD0dZG9WC/BcyqRPU3S6BI6ipIXJggFvsman8vI5kNggwFtQwLIKiLwokBix9o
JB9vx6vemEQmLBHYvfY+8GcrN40j0E7xjTwytGmhHVS8lHX5odTP6QP1L84qWZirbwYlrfquKWpu
j3/m/pO1QyG9PyXnNnkUFxme63bYUdEDIN7q2m5mxOmr8yeaed2qH0dUggk9j9/IdFUDsJZsKlBn
M6/IkhWLJytmmiSCAeuGyYrJKEtwvxuc73z7tlVnXBGi2qQ4vJ8E52CF6X5kqxiDltCCxYTUY7Ii
MuDqzqd4G4k+X3vhYfiEyUksyzLrDoeiZnZFVLHMesSIg1WVSy7JFrgQ79CeNqSFVQQsy4pn3F6Z
AhxESzhnr29o6hOaldTIlZ2Vg4oxsE/LYlaq90rmeE53i9gD7uPFu8CC0gA3JRBdpXwL+0LPFXgU
szOugVgXYdP800nJjNnz7g5qVX88POTJYHOR4GReT2NBPHbQF92CMMuldN2J2TzEm98MnpyE5bKZ
jXLnCa2rbrh+tgHKtc/Jnbxet6S33qPq0HJhiG1IIHiVk3LXeIYaxqsY7CeFe/RY18bwT/olWjcK
QP1kBJ/3ILVPOFQYZO7fMX2FLnemzYIzxhyojDaAy4I3p0v3ZD4V0ADJNZCm6zdK99n3lpgc/GKe
OLUvDsvoT/hGTyZpiQhKO0p+mBHKiNGtuqxRem3TnGLBD4cIBMKKW1aP+5OpEpIDiTCnC8V9a3Gt
LXfv90/s4hNRsVbiZKml88tvFBU7F6VMIdq2DuVUWQ4ScOPyF1XsootS1KCGVc36lKr+oyOHM0d3
3ID0JTUl8ltBV8B2nP7X0ygWwEpaPL731tZqJnYwfk0/nCBU0ql9iXZCpGYpJpJwwbjAwVOQBD4V
fY949YS7FmLUQvxo+yChGOduRlTReoIB8QnFOsDPk6jq22W1E5pqSPABgcHfg4obnvT6LTeq6doi
M0AUqYKtYRgo6IPXLUNoNfOYdVXP+nCsiXMUROgrgunfmKBPBKHqMWFc81MDDPbJnck9F5xrsalA
KKyITy7fR1t7eYpAMwud7w+7u4904kD6BcyVcqhq5pY6A6jpluVEnwVLjmUup4V1A6e9GvDbL+ti
mJSVVNLtPHValMvvCKYWuYB7tN/2Z4rDOP3/bQNb5yJTWQVNsYH4F3qFPNkpO2w3N2xAM2l/IHL4
G9p+Cm8obvo4nfRaHXZaUHda/b1oojWTB5HSS3bufKmMOmUL9C7aIXlwnoCTWhIMjzV5ciL8d9yG
ktDNlg0Sm9Qf5ymcJVK6WwJERO8UDrZmDcAB9jh3MUw2hjZ8oIIUD2V7ttKjtXDN60nGIhAOPNLu
2PRkPSrW/sm04BtxgaTE8NaQLrKSTlaknke8LwzztXpMdkD4G0vJXMAvHUQXQph2pgrCWC+2R52/
I+0s1HV0srsGpTKhpTU/9/UdyBw8pMd4A72nf6YtJktFWZfgXm57+8cvKEJ1b2PpKURn3k1DaYs4
GA3gUk25Z6DfkIi3XCJiqe5ggSBVKlae8jau7Y2PqMwt0RKsYl1y0w5lMfHSrFDqXVPCDwgQPTef
dZ7djSNgn6ISpBvenqR6fpqhEIkhvf8C4LBcbapgF/1/E632RG4gSFLayRyrSFbVd6+XTz0aqCuc
71LkDvNCGvyUUbo4Kq/Fc2ZjR4g1ZAtHhjZd/4p9fxFN7ZUjPq1Vdh0SU1BrVL3JYS4FaWYjYE9R
Mwo2wiCIPBX+G2o51iUD64VPiBVcGL6P1K8ZSji0a4ydZdMtELPfnr1L2Vqeryczlp7pOR9IPtSp
GWzsLmYow2VbdRd7XdLqFerdO5AEgH27nWd7I7ou+Mt4T5wqwZHOB//iPva1VRWxOoI3CrTWTPos
kHo+wMbuUp88WYwPVYnC1r1m1gOa6C+wV36KpzBQFtxBDvQRAJnrMJ4r8gso9gTgQFi47ruo81Fj
l9HaBeN1woSezT3piAPV3d8El7psxDLhXCP31B7qVaN7tIxhLOpNJZ1wAQXbUvW+QTXMl1mNwmg4
aMrAOpm/X/hZOk8VVKe2nmXq3GuIjtSsXt/fpVq3zzHxa+WspdzVsqHi60BcnWKYvkT6ht2u03/v
bmhZ29w2zQboxZANdch6UGtKCpm+6MGJtLQ7dHm3IkWXRx4O/PHhQ5zg4Oug7OMYGak1r9kC6vM8
QFPmRrPgvGovqzFbFYsNGeIQ7/I+11RFzL6i5Ji01L8SVYSKf4AOwjDxKo0SnCtbqB6kDKrHJvV7
Pk6zoR9T8qvLxtJwND33qg8BEwVxR7J9WtNK95A2XHCgvu9Z+yiaVDGI/nq5qaQc2swHMREslW+c
8Fenn/21mGd7iDYpmOnz+r5Wxgd4ld9utVaSoIjcnmepGKZw/hhtWJqPb9FfLpyAz3tyiiOGtbUr
wkBMZqsM1cGo26XHdx7uQAOIL0jpAsiLapw7Axnnpw/TZ59yAH3PotcrtxCO8weB9Nm4/llFrZBD
VU28icQZn5yfZdqR3vJNkr9ntK3T9Uw9t3Cs0FxLD2B/mREU8U09KsK0RF5cH+kLOqZoJbzMiSKa
4Xg/AfYVWPQj8VOAukyiukHLVj2xYoNy4NdRDeVvMVZnRfTWtgEmb/8d/dRNjzcPw4BzpLMffvKS
StgAvzCRGR9aIwbx5hf2d6CRo/J/+LzVp8rZJxisEF9erYrJQsd+M43ZSN96oR+hxB+8cVyAITZV
jJn3fufPOE/mrjBm3kqiKbIhVpwS1CbxNHbMZQzKxCv/BU5BP+RZ4/NNGViMZqbofYB3eaGMTVvY
vpZ1tTsoy5pU4yd028fBeJ6H2evJKTLnObLhuEbsVR6FwH3ZGkJ3wGCmul5ACN5FDCYZDPs40Xy3
1r/43U5Q/LSKyJNIxqhys4TZp4pL51/5x/LUx/drD2hc+ASf7/VLwq+X/rEY7SfaDT60II/2Qylu
3G/oJ5DtwV5tFq7M1JfDlxTOE8kt5/8Jy4OZeD9vc8F78RHS/JZ5ieFi/XgBwbgRNRiRjqAGF+rg
m63kHqd7THomIj0U/CT9c+0womvI2Xj/IU+69peCKXDTZ/fp46ai4YBQCahqj8Q80G0iIb4B59hb
xaiIsdiJ184MU150J9lPSELMngUsjNrkmRhN+J0nUCwOyzt6uJ2R0ozK9PJG7dExSAv68JKMxVGq
xdeugfOFiM2UWG0zdQEywfv19L0priIK9DFNziXePPBYHhRkqUAVBZKWGJqRaa61E6ugej5C9TZJ
5IzhpNjn3XVZH9fQvyFQn8g5UfP0KNIZGxbah/PedEUVH2xkb7jtygphFN617ZfmSwLsRkUIMQZi
iQnVo8O7gk+Lx/k5+98IibDdMIAIW5C3crH9dEAtToGMtmtRxT7BlNnjGdYHsMZDC9H2m07mwD+S
IPTLkNlkGRAXKeqzzP9Ix22sGo9NnSnqs+hTU42UKtb8qBw7Qat0uFS/tZkC/IEWFNC7Df+lndcX
+MzvgYNP7nVpKvAndY7UfPNTV5pDbYC0TughxqteD4HG9Hhpk7Yllq4XA+Uy0t+vyxP2y/PVwNO1
mboUHclnLiPhDhFBsvHjNz8SN4nca9LsFJUlnT6IN/av7FGKKanBjtYgIRlpYgmZQf2GNS2vN8Gs
Lknljd2ETuCnUIShToSpmkfk0aiRuMWD1d9d14wYk0gNMJLpUVXlK2uAphED38GiLU5MqpL3B66d
fzCu8d5SaQ2sgYhAyxMhSf27r7j37W9rug7nW1MzOUE0kugJWhqlJQbozOKmQhZrTZNyj4kNpFdr
hsWxPdD3o9kRoh4n0hOhmaPg5QOjv42DRAhI0/Pq167f5X6SIi//oiOlzE2UepUZxm5ENWQKzZXI
PTWONFrNmUxzrI2e6JMVM3H0QCDzqTajEH8UZpx/p3NbJ4d07SDyzY3ci6b6KpqBOODQb+f+PnnH
bCLPaI9IMcYg90k5UHCgvEkz/J0z2o9N51fRRHzyRh1V3u1n3Gs0N8zoA5is9LMlsQaF3J6DGBsy
y1v4Ziwg67JeIUbIPZScpi9C2nq9dptoTx2shKHsppCy/pmqw7Ei16R4ZW2+UcEHozUDZ+ORgF76
m0Uo8jeqjhoHz+xE9RxuvG/QEFayqLpNZaVLL1jVqvoDEJo6KUZohuRISGYM+JyQYouxrcB0zfJm
ONbXGULfWiuNQORfEZKA56dN/3wYYvKzwU8paIGZrkXpjHIqiwD7Gj1v6FkYbnXhJ0LKg2Od8BIU
Lr+U/UvNBtqx38Kz2ZSMcT0dVi9vUIv4Ud2WEXIOVO0sey0NdSb2EOL+rLGApDzZrJvMf5GDpLVo
PLkp92vhezTVlBu/ARxQU99bX2u65k2XwHl8BB0Vxsb+xqhrevtu95z8YNcz1Pn4hu7mOwgzXxYs
ez+bxPC0i+PPtzENbp0k5gp/zuiURk5Jnl8u/VBaXXOzHZvB11CLNCfDlT1E7suqTo2GUppvizFB
8aD4v8jhHjb3GDu8+7/tHulLb9KCUh8Eke9+QSVs6qwA0RALowQkdrbIGA7Kh6WtWc30TAmrc8oD
mB1OWkrhM5KIgRt3v6ZUl5tkpj/O+0s2+FsQye/daawDPaWbZo8yItxbZL056de5BifGYLFkYUez
jXs9lBYY0wXYO9fX2IXyjMpUNYky0jCIskMXh7sOoFy7mdMA8ORvJyT58HNnnWTGmdE2pDMOKfJN
5i0E1+q+GsHz3298kUTe13mhROtnw/DZPmw7psRbqqwkgY3TLzFVagA583vGoJE3S2Fjvopi/hk1
MUXEl++/48t4L4LTM2tv/kwT6z+HsvPYfLDQIu7BqfAEmG6uOBHBR/lcPLDiyXzWCAg1Gospa4DL
i+sf9VYtcGdZerrxvanFJ7TWEAP42INFc5bcCp3vHRlC0WGNF/Nvb8V+a05v46dNKlrd1nPtxIz/
TbI8F6u+IQ3n2Y/6dG+1+NgK64HWPAMg90P0GagwLzQbY5ZmeK7B+QDrZ4BXltXYgbIuP/fEt6Mg
z8qRLK0ChOmPWONspwxcmqZ/BGHRfsFbUhKoPKAlos3lZFDSMBSL6CbzJ+amGRfD/E2W7FN8sAA/
erRDqNomJrmwTtYE+G/cp0BMWonOjBIx5PGrY9KKroMpCMuLtgTcx57ZmR1lGYAtVAosXAfNzw16
jvgb3MUaJs3BAbXoaBRMVBYmXddysvkBVfHA4xa0JLR21euxjEwihXxP+cv/oXSiO95xUdN1egYF
eBotiIl0KjGWeW56sxzBGnl0e6nzfnqDFkD+zaEIVb2Jjpi+0rVSpfYOPpn0bB64ehCBaxVXgi45
twZTM17bfd2nyzi0+VM2DrZTUTGpxC3+/xOqfI5fNoDbG8jiYriJQUc4F0vUC6oHrb34IMOJTjZP
F/x8Xn/OCrog9WxwENU0VT65XgGLzDq1uWv2B75vM9AwP5JbPzdGxVenLR5kBc0yDsoaAvrzAUOK
8cudIKNwXYjrgqTVPgSmRWZcd4pm5Uo36mxJPye3ZXeFAAxgGIwVkJBggS1p/FVYjDVMh+NxNlDn
QPPdfFWSoWmMrJnVXYZ0MpWKW8Rgx8hRkiFJM1wCp2EANUyvU23jrb/d4DJqDHyB7t1KBfVqMx8m
NtZF9iaIBoQr6/F5mSrLgARJGG5k2jB/yDtOZogp8dcyN9RlT6gsVLAIdjWRcN6dovNLNh+uSbtM
y8WjAX96U2CSF1mTrQ+UUDTFyXBKLZztgJFDl4kHYAsB/OlMnL6un288ABwZANKC4cxvuhe+XMvG
Fd2CbwSVGJywfXmEXkdUNIN3om8o1t9EBgqWIUBvxgkuhQRtIj4nXB4BTCgNC/RpSr02XjjC0w2n
OvkEGkcQe4fVxtrs+snrPK5IQHKm5qIgE6UoEeTtp0dAcSuI0iN4MGgWD/PLs3FJyXevNpP932Iq
ooCEEWcxGzQCB8fJn2eO2Pd165xqu54JUnwC+68WkMRMG7Aiy+WaTrMM+5e3mb/e5AFbaFBYaHf9
ZRDpdewhdjzUOobVRFl7UVlFlojOFwYNMcMtHa55BE+JcASd0bAohc5AJbNunfVEI9t1HJwZcFmI
m5ju1TaOevmX00nf9dQ4hFU9vOLiZ1aL5pYAlryu9UBjzByA48lQ/0tilC6M4QsGcD5Q/W0UsXiP
ZYbitVcbb/Bhu4gIw3uYLhKH281Ue+2KRW6BrRTs4DPcCKF2xMbXW34XsoW5mkZEnbMg/0+f594x
9qIuQFO2bk3hjyHeo4+Js9n/kFZritiieV19L0Xe+2LnLDzWI3jzsaeRgkCxYbJWORSrRmAbz3Ar
fMVXN90J4xeWJR5EABA0Vey3bEwZvO9UWd5x6WTJLn63gOOjCSovA+QrHmM7rI3Nn71W9KPfXHOy
+76veqU48DxnmtYPeKGL3i1LZq77PIoVrnk10Z9ciHfnmTco2M80QSkps/mMxKW0jANSshhDJrnu
srUEQUd8KjO+yUvUGphAYq9Sn9ScyGvkyLwIg2lZ903ywDgOR+Tu3C7kuUJNXDwRUSdFq8WJ8+1H
PBbzXVnbVsJh2ten9YGYMBfWWhY8wTLKHi46LdvFR2mmrwVQNYUDkjN5RO19CoSu8xXcN1AQrNib
aeq85VD0DBE3MyiQgqVzW2Usqnw91gwhE0c9qEjPbDdmTTf+znNTAP21Ba60cKfw1DVpv08ygOvZ
65v2WmMWUv+YcZJv1lmhHm5W/9WZ4nKBPV/MLFv5A5SWdk3HYzjyaseyAddACVLe7vS/FVvEnOlT
i2ZMMD/5n3Pg/jqwwtxw9Wdc2xt+BlwCzotfDSKlDCb/wINRGq2l1fUqn1BSx/pqhclFsQbTYIUZ
hW488KlS7nnv+Zch1KqXsw39tVZTE1Kd1e3gKAp7pIT8DbOsh7fzO+li7o+dqtP5iK3d08JIE0M2
qS4kJw10aOAMHJMbsI3exQ7mDaH8tADXZZQo4ZI4GT0uC8Guk1zqM6f35D/aonmwRMUbFdYTpD7G
11mDPaaaOI4JVGro+lYzkIpaL34QIMBXY8Sy+9nnnv1/lq+BvZAnXJCrfosFx/zMgiqtykCmw912
Zo1K5ud/HXsq2ZRW/AtlpuxAgiGXd8xnWbR5jbaodozPocinTF9dyS/cuRlutwR2beJDfU/za1dI
GKxln6FTJ25T4mk9U6wMloIb9+QzIy+RKEx5RXTbdiNK7GlXB7NabSyVClc2V1KfuOtpaFpAfbLp
KDXLYqX7CohWt1GdevKA4MXXwLuH3x6JtNaLyoRIIgTSmG2e8HgVgrI9CCN0Kj8hh8DrrJ7BKKg1
GVMRstqVDQoGchc/PToT5Ox6QieFT1ZLpS1u6eunJwQCIIvHtueytXeX3CMI/UgGVZrs8EnwgQ7c
9Tz4DVkOwIKy1bwrKoG1+l2uVH788Cr3248LAIRlYC/tih0EIb0Gdc5fxld9r/GhzoiO1ghOIzkk
gXBf7PrQwPWKGBa6v8CwzQUA8Ez9xQM7euQ3pi4EV//lT5G0RkG2ECxETSGdVT7naUw/QLMp1Csv
xfWfTmq9s6TQo48mz3l7L+84MslgTWhUY1p3YjhpgWfZeYiazTdTgH+OAf+wSnIfqPH3bYdRerFV
FIovZDfdfdh/Lb6wZvnE0xTzu7Jvpal3zf0MCcffVF+vhSJuVWy3PkEIqjjeKKoBzzHoPhHlBj2D
R7bfNPGRAiw1KQ3mI0SRFMAQuolKaG0nArd10homaQfzDZfGjNnTCcPzjJOkhZGZ6+9JNajWHyNx
AGR95c1bUvvpYyF1X5CYYjzGXuHim2gwhOKP4l/ccakpIc2f5dce97NnKi1BOSgJG2vLQ1S0z+vr
pRBVXrvdMApUAEQMT9Mp5e/mSlMGjLFa/74Uve8PbNIIFXrvmTFHiESoaH/o8b6eRMyL8HvETIum
SpMXodEny59cJcDsyFQYrHoMWcD0kqOkITVJ5qPGgtFplqrNqxQ5QbSZ3pqOVPCnYP0v0K9sAcLv
Y9EMhInnTwlb3S7U2X9238F5AUEdX/2vPcDRaSVkQiH7Cma95YfckAoni8fjw9FfrXG03WlUCDUN
mQKtR5mtEKYj2F7XsyY69S4lRg13dd2Pt2Uhi7clnyvcOKmYan7gl+lUglFZnLBAQV7n+bAdtiu7
au2886WboNbqpIXc49ekpAZoa7ZAJv3A8geQdx18NJsGfVK9QijBzymPK/tH6Jq1kDVfMWYVRnrK
cU01DFaQu3jGtlIaAy2wzJ+pkL4PrxwCBQhqBd4fIoiMegcveVvJjG//aoTxLN11U3kRu28Qaz9s
jRJ0fWeR8cBAOjpN5d5G5NrsTB8NRWPtb/BTqfw6wpSHpeAzuvd+QJZLnxd9m7hUBjD7S/VsWp5R
xxDIocJGol9uFqQJAr9xKQd2q1SLiM9izviTszLupghZvU3RW8Q05A8QN+UOMZY4LxskjuDfYJrM
QKiOXnCJZM0Z/k2+2/R7imX6tVf8kxo3A5+sV1VmxUtjMP8cPMhaE+swr8IKrqwg356Ivf/M6hZx
BtlB9ymECeUOnQQs37nxc1b9G98gukbeFCEQtUweGp1LfdgG4saFbWJixyxMWqMYMXBzPcOUlPGR
PoAjKJNH2RR633w+YJaQE1GOobjy1r9IO/65FcBjMNqnsz92dZge/EZSQAtulGhKo/1w7yKX7zwd
gzVbuf4vpL66EOe5bLM9SluuR17SlWojvAfWMfuP19LcJr2GbyhU2QipWLhPBIgktbaXw2O4Hndc
p//0T7H6PqogPSY2UtjfREG/Sjjv78bBwExvM8kfLZ3zQHfG+Iw7MT/mw7oo7VtIHXIbH4WgSPDC
rckYeJrYc6kI0GVHEpN2x6fLSpMxrDl/miBsJUmAQFAhUZUazXVXu57x6unF6gQOpPVlDufiNScs
zD0o5aJ/Cy71580sWMxEbdhGtg2irfPTYGaVMHsvt4V/MA84hcwKdhxtJVBDJDw9kcVIWAcwogO9
Yv3anEQNvrvRq1HTsmMK455565FFD0slT+1QJ+uPPZKW/c6Pv7Ari+yVi37Py36TcGNacMNok84p
OxPrzC3mEyn1wBkA7zT9o48NrRhySTAotGhk6Hz/c8yb2Wzw8vmYmN5vtgcq2bR5jNnTEjP2YFVb
FV5PCkg+diPw0zki/OgM0Y2WwjnLWy1nSSEsviTeIBuBz96pu+xH0EE6Rj2Mp5f507+HEdac/2Bk
XupupV+bdNDtGhEghnbN59XdAp4HtelMYYpFZ6U2kHelXS2WgGr1QpjbIFjP6SSLX1Al9gkrfDlf
JWGfEKayd9xNe1R60KP+9W2ZZY3sMrazINOlz6c3y0/65E7jK3oYt6XJSvNkyhWQzghCYFppLaIZ
JQzlFC6xyNvf9JU8ibJO/7VQmMeyN/KmUIDtDDQa+XG2xtfj5TqxWEBewd6v5Xz6JDO6/10jmlDh
+id5nj6G/IfYp6z9zVixe+61vAfEidJzzBZg0jiHoHsfpp3sFgtxeAu1/oM9T+6Hj+CaR+Ud3+i3
EHRuI19camgj+2jpfrq4s6fgX/myTXc/1XOfzuxBDWWzo3B2QurBpe8YVPABlmd7+tarQmcyGPur
2J6ysjDmbJcvzmMlfe4JDnRvgztXkUWki7YpxtwE8x4IMzwMhARerg8fZuyGoi9nDXfETXdAl360
p711UClnQcHV46/OVArmz1XINj3NPojIiePGazOufL64EVB3l/K9eyLVo1700tVg7pmUg7eyCcLJ
FwAttvD8F5+LdSUrxy1+lckoiC78Jzw/dcwBtJI1WtG8aPDpdmjS7H0ICom2oXckSE5WCEUFJI+h
kr9SBJmrNx7LYsYg9GGWR77afSOWjd9diAz3Hm6Qt6l6NuTPqtkC4Ce1pE6U+DXuVDVZxqvt26Ce
VJ0r1j1Lmbn+ouBSdJyNQvZStZMQ1Va3HIEe/6iNgpAzwiITdZG+FH0drrsg1FCSukIBw8pu233f
AWd64CWzSf2mj28y1AhbhAAI+3nh9EcMQP99sJ0YMQ4aYNXmoqLAL29AyrKxWDW5tkQ+rbkNOWdb
EsTLGLX8knEI6lWBf3Z23maNWXak/VGgG+V7L/uCF0r+qNM6gSMuwKsTyRoCOk9ZbEFmknk1kLRD
VrcyXdvFz/2q4Amc/fPUPgZcV971X8A=
`protect end_protected
