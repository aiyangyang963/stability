-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lqAP5YjK2txCEkmJQ/q7Wn2ubsmoEi3OjmKIruxHuz8Nyt+BFKVYOkVN3rxWN6aqKoJWhrVmU/8m
+CTW/LYrDZWZJS/TIfFRDWLWxB5xNB0RpK5xzvcWYF+4868NSrEB6I/yUeprmfJn+GYeb2g3StbG
/R+u/6M/IlYbO2U3hx70AIIybDFY8L/6areO8DKAaA/SPDxJnsC4lPFk9fyEFOi8AKBGtDpto5Jj
DxqfMbrYy7fkn96ELCxRh/OMGkeL6H9P/WnY5gUDydLJgIz8Pi7Xm0cjcfk5AWcnDUNzKpjCv2Wz
A85soy1ntLZDxM2p3RlRAm279p7z8EhF9TGUvg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
PBnL7wLXrwayF/wBRdKNvfMHFpi76oQ1hX6jAZd98x2lArMg13cKs/kPb9Q6xNtR+hVlU2cibyH+
z9uL2adQ+hr16TrFwyzyaIol8+9OYQVCoANDqqmhPGsFKajS7UrpCm1EB/aCFI9elXIDcv/6mGql
uSqSV5hTNcFZSKV979wUm3d4mep6iy2gbz3KS26yv4dUcXBPyJGRco9Has6U2C/JkX3wUvvGVgQF
jFCM2pz83rR1J7z39CUvy5fx2dT+XAQxdrfqbk6ifrbruz/fCfs1/+jXa6QRB/g2PC28bBUYTVrQ
YxiKOgzQlMt/ouqH3p4oYtHmyB7K40rkPZFrPSFPaU2odpK7pQJ3vU+LptVlJdCoxQSLDOnmKi75
F2ikmpU7zmdCfsVNvpon/Es8q75e4tVwH36XY4Ub5CLaqZt6MZCa/Pdj+GXqOF4QfN9iGdh4XA/T
yUW8rfnblw8aJ7vVR5SbeGyzX28vhMsdVb547uKc35rrcJ+rQ/6AtyZbNOkGwo5FOnU5644hvzEV
Du8EPc68dNlBZBJrUPWnEXObUVxam1ytqr4Bvk/4nwXjOwpDsyBFivpR+vMChlTsVPx//gJ2aiPb
Ef0OxHgshiWiN4b+HB53UIzXXl81sgax1FzfYrGQB6+/cC+GcAic9lAewHt/MAW+APmgW7DC4Vxz
ikkbqNnh+kTaxAxvcBXcrdwEZ/z4tnoS9zrh2vePjxJG7l06i/1+AkLsckaLfpF1HRbHtmQz6aBd
gjeHd9bjPrtUHssC/nkxCX5kqW7vC02eYRZ1JrgAmDtbb8cfLe9Js0vrs2FBFh422QqJmnzX+xlJ
/Q6bXx4hhXQ2pBgKXgBWSkjUBA/9UgZ9mXAxoHv5J5661nX8UcbXOzia2bpG/UJ37z7u3imA9KUV
hTZsz10inDjIJ16fdfbIQ7vd9yZeCqgvqMaic0EH1Mbo5bCEkOpskaRH/eUGYWkrozmmypqoR1cX
Wqk2YwR44aANgBhoQTRLd5wD7T0c+njiRDGhnKtMKb5NnYYXVRteTiY8BV2MyoUa8mEoWOhygcE/
WRZT0VKBVW2UvPo2g/TdzmJbgMipp1NmA+ZnZeHm6BON+ke4ptxZRxGcX1bssIjpaz0MXFNUwUXu
F/Oida5pKWhBMMiEY96gUH5gw/E54VTat8HnRReyge51TcUend29kvCM/aoSuFReZLLrN6zJ06gV
Z54IzRn6+bxjkSTT5+3CF1+N1qBZuHpyr18SEfJq7j5gKYp7BGR8UO3hz0yw3ZclKzBESe2AhkCD
tSgGWGaxX6KHVoqgsxKmy3Ds/qAI4OWAGScAD7oJi0fmSUpZ50RdcVBYotDUz0obsPT/koIA/f5R
v7uPTG3OMuoatsOiJn/D640SHpKMRsQBWVvAWZ0z57cICBoXigCf5Wp67Sez89y4oQ4WsVJtMHiX
gpPlXTNQiA7Mx78sOv00T3VUT2j0XEK3H95WjNPeDbHHh9ZSXGKfYgLStCKmEScND55XVyEiXyvU
/rysy3fxtuAm+/C9hMakuMXc7NDwn+KxzUhdIGZQ8tATPrewY6MhM9zV0u+6ZJtC5Hn/ie1on5mr
Hfqh4hHu2Q52Wv4z6b0SLLThiPZarVLmIPfnFH15Yy9dL5gW3MS6NkpX6W8+Er4c6UZvAQWSk/jQ
haD/s0MlP1yqNMN0odSiV9yQuFwWcdjz0zY4cXa7mXDkjvarmwatW4MkwghiWhO9/lyAbcMLSGDl
UfoQLw2H/WWdjqtbnEOnjuZ2Ovp572KHn5qbb78KTlxY2EHmzRWJo+i4Fp+k3mh7KJA4ib2y5cdH
FOPLzEEAUjuzGMyiboyn5EwAsgN6Q689t7dxpe8WsG5NNjT3psubiIZav/QpMC+Np+qXrjyyREMn
yXj0B8aMEOJTAtg+vwSZedMFZzzsI9vttMy21NnOyCJvPAKLHWlt102adTELnmrTDwvFwQP/S/n9
BaswttF+exCJvzAM7sQdrIK1bBA7e2H58rmXxQIKp62dpUQUoeCjOvc1GDG1Pc3p8mp9Z4tAxAZf
ejDaB56v5znq6nbCX7iVeA4uL13x3UG+vhkrEDpbJGN//ihiMgytnhlUnOr7+/OB98Xj46UbxOYH
GRcUYs0os/MmoqbEI4lwowc94cXPEmpFx7VZLSBVDoAJ1jAmvgLn5FH1RGopNpbFlFNwsFIIeKlo
Vy1XNCL4rrIvc5Zo47Xt+6F5UALjVmvJyir6fPO0RmEwSFSzJ1Z5ROoGlo7qdPT8dpEYjZfGzMi+
A/EstcRd0UFCr6B7oloU6Ss8jdgIJhrHgh9MGhcKO6nckR9FB17LL/CTq7A1EXkJ2opjYyRyG0rm
jCl4ovvoVJqdekgF4/mLjq0COo2gclyE7g0LXcDrZ3/yahcLU7l5Mz+5rhsgeeNMNgjlBsdX98cV
NYLYl6PQMREF9Do36eWWl9W2/fFZvT48BxusS3IpfouhZo3rRZWO9xU2qq0LRNoCjBe4bmspQtuq
NmD6M9bD+e2AsAYdzBryzUlTEDV9LSiDtkPxZ/I8xSkBxwGxrCTI6HaLfNy5TREvu4+JSubDW2Cg
IZAIc2ox7XspmJS5CfdoUYB3HNKsHm5hO3mHqWStBnkzjLz99dNg4uUeYI7+CEMJS8FgI3R7xjF/
C1/+vnq5l1F6cNZveIrhDaWcB79qumuW24HjeH7NqV/SKfhEHB4wV+p0q6rVyDT0kcIa6r2DzVlc
UmmN0F2bp8q++oNPCOH4prybF3f42X6NtYoe1d5/E1sKyl8g3IbBTnph5LX3y4nasx7vCkGzOp4/
V6WpWP33FFW7oJWHLLdN0GQDJo4lODrkZjnujhAp9WmUV7NVGqQuXsd0uqgkRfwN/ak/2VrBJv5s
CnhOsSAEtfH0GtUXDWvzCeoO6f6jfdzQVfWXtgio8lyty57q1dhu97IAn5mrfsV+otKOFsMyB/QP
ymhyzrmNBKtIaqBDYbNXOjObqcf76F13PKI/GQ1FI4iMCo+6uQn2hrUZ3eY5Q/neJA3UsIco46mZ
nR6GBIrv+r/KsfP0dw9yT3ukM15efW3PprlXlIYvmMjMoN5HnDh4pof6xfTKb2amNARxrEw7oy1x
+/E/xcwzE+ccT57SQ+AZY+GjqSDPfGkL91X2DEGCbmqQRivVntvwsLBHYz2fwVyhMH5Ek6CJ3t/K
CX5BUY4bHHlLDJGEyVO0QbhDJT4ZCLuJc0gcGHykduD/dp7cISVXawsNLtpp4TzbpVtF0Byo9blT
G2tT5d/ffzWLGbs6ZdCDds9fYx5cbJwbQ5NXnbBVwAreLjX1qDBQz0pnQRbMnmjej9gLcYVDLn/a
mY+Ybf7pX4lvwB0I8a0i+kb7RU+oWCB8miztmc0/yfNkIXIl40ikC8z6CrHNBElEU1tJSMRVPaZW
q1k4ll15vj5r/P0uoVH9p9sYrePLL9Ujs4JFzTPtEdAQGMQ8gyWzKvp7N/oGI1h1JF2NQDPSVjLz
cGqj09uawx3xpLrP7i8WgUJpTciAmdTi1r91NnaWd9LZWzovR/Bh2VPCZeaVimxVcoc1L+SpJQ6u
vO4e6iDrlUD3Z1oQjHrJjrXbm62iPv4tSNIJJPu1Rj30buwKlnNLCAg5tdNNl53rOvl08R0KO7X7
uTwVfyr+/frOxHy4BJ101jHX8fzokcPfD7nGVytLtWTXNoNQgLDax4lath3t57U90z257fUxDR2l
MJZPxK6PUJlmXCpfe8GF/mEPZHwYwe+YRn/9S56El8zvtwa+d5JxBvASX8/rWs5Em3jpKyejdmeI
cj+gFoJ+ede7dKHGB8LnNaB6d7ZqNljtSH/5cRzFyZx/RVoqeobQpaELnN3wpeQOqZu7HHn7oYpZ
y2u+S0noKFiNFMjhPiplgU97qs21P93y/HgreZhvnneRIlrirG/Jv0LVEWQSOcCvDfxp3/TIgUgR
QSWIWyOfy1q+tv6RT9S2BQyWx+OUZbRhfHg6rKKTVgeSxvLCbZ1nbbUcyDBN2FBnrpCDB9JulC8U
Q3F3Q5AclaWNU0RMfjytbE5ErEDboSbVKfajjibvfppMuBL/lyECJF+iCAV85/rxYgkRjlBm0rWS
VQ3wUYW4CwBAp0q3xo2NIEJH2sFWgY0NqyiezJIPOScK50j+L/xLgzbAXaOvbRfsqOnCdx8Gvg9B
cWzlS+y86pLtrM7RRaQDaT8D052YOsSa+FYdhrcBGV6MYkEIRoXEIbr2mMUbpwXMeGl8bWfzc2DL
q0PFcHlusSkdLpr0lipMHNYIv6u2Zedfj3D64FJkYylHVN238S/UC0nrp+0ecHmxGbJfbsNgiKcT
v/9dGi9hDql/2AQTSM8IiNn1zv5w8ZrT7HDRUSsjtVmXWu6err0oO7MbxxXrFTzLMMdu77QgV6Ou
bDtohJIPjKwLE4ggtQ5NVeC4u0Jp8Gpfl4Axv1GSHGZVXJ91V2I6uOtaBGfiyFvB3RfDCepxFcLW
7VX0GeiysWZosClhra5p2OtMuYCNnBh70svNUaS3+2VQxlS4bS8o1pVQormceC6znYZpsRJA9U8z
42wu14nfDYoQe4pO+1Gj+GIo3wgnZ0SgXoEcyhG1KqU+DE2MO1Yy6YaSLFhDJJlMs0m9wrzN0vFF
62ZBfGOd7h8euDcXGpBam+zBlZ+2WhdOiWcdpo1D4crIUUAqqFlVgy0Mccno1r1792BX3oHz/yZX
f+gTg+kWUgdPD8s/C53uWEOwVxHH4T7NlG2lPQ1ZJ4IlmoNxb3ywcE0YyF5TltYD35ApGKDDGPnI
EKi0hncYncPtN8WvGHfi3JSyBmbfr3+Vohzp6K7NsgoEM21xyIPt2LAUQWbsilZ/8Bn46g0Z7JE6
T4ZB0bobRqtXZ+HiYTauuNWQ36WhQf8jYchdL/iZHk1kCgK2owTzBsVhVSR+h9ooSILJ+E6654uD
vMI+KYqYd/PUKbd2kbViSxLjSVwklu6Wz/jD1jXo+hy/7BZhJiuCxvy9dm6lPPVZ8APRjIw1RhhV
Lop0SWmOfsAzKnPb7oxgpzRYPzSW+h8P71tNDm1zFd4mSjRUv7B6KL4cRBVCea2+HjGw2v8EE4YO
XbZGG90fUgF0Vv9PaA9KQ8OJbfzeM21E8FE06koMj5vOKixUvMn9SxvHBygRLsc1angOnTHNIYBJ
73iW4OGP7DQxK5lIq+rqNLRF5ajIEvIUWEAYAzdk6yHzVa1lNpFnJbe1FUbU1WEJ7t/Zza/UAvei
beiJYi9XgFyxMikfYAX73SCxc8QRRXmkB7oVA6QH19XbM0YlFVzVdJGsn3z4wIjsrdsH1Y1/NeTT
Td6PbLmkKUsfdPsiovVMUEDtcM+9XwD21rHH026Nk4IfOezIFE9fTTxBcc7cl9iW5J/XMOnHX5Ax
MuMqfruSnsVkCIl8/7vohLsrHG+SfSVKHfh+JmnO6gaaZw0oRwH/9jUoSobw40s4hVpcPG7mbK5K
mgXdUjSfB8OLVR6Pl9x2prrfyPcPbsx4D2HUG3UZ/TBp9C+ZQMeWB8lqTP1RONEhhnFO67/Juuyf
rmnS8aGXwkO6RsY15cCB43Qrp9E5/yKc4zZ0emAw8ASF2X1EqHDOd5I8hkmg1onBTsmN/aXXICBf
DM3xJdamlxgDUmOu19X+D5a0QX1WK1SLrrraVItq9qBlIJ5/re8HfLqzxJeHgpjfnHWShV29pDzV
hHNioRGtLXt9GQIj757Ew+F7hYu2Hkjh1s19uGy5PuD6+D6qFH7qKPpBrwBq1d4xFG9D6w25OFaK
cHwxqtkHtgXPmFVl1whXsB6sD3nD45C3khMhGwYSov1IpJWMfnO1vWuX+6CEnjSu5xubg7iDzwPq
Fsat4iS8uKb/hWaKWdq85oTfy+gtDEifErnQg6Lyc7B3F9yF1j6XAfHF4XSgUahwMZYL4m4ONyhk
iYD+x09VHWe7v/uLgeoacozfTlOmQaNLvJ5labazzIrUx/nFHB24ittWjqd2YhKkN0KMnUkElryG
y1B6rLvNmeMjHA4zhvHQh782GwariqIuBKd/2XilYtaYKstlOWuivN6GKHcUYayCRO3lOytzxnQ1
hG845gG0FjR1WKpWJTfoxxd4mAm3VWpGQWmPSibL+NV+nufUm+G1ON4LgWrDrH66ppZHQPlDUXVy
/ZrhpqJn/NvLroF9h3XK3B4tsZ3RIysQZzmXE53ceJoc/Fs8OBVjYCJDhu4YlDRRVACfrU9uWGxS
Eqr3wPTmOt0dkAFbrEZ1NwBCx4mqB8QqOIJDWnX7mO7WdXrDK+3vK9WG/sN+AdD6WG3YeULnr6hx
sxOX/uuPRKXRLTwlDRXihpQ+4GGj0OKHNrZzLHC/pwV30Zp89UCVAy2bruPURKMIeKxFt5TxNz0f
1UUAcFBYa7RST80Ga1WSb2wGsrlC1OTE+7MTREjQrPtLoTwM78quy7T+NjGfFV/3nR3tTD3BddTN
cyYwKgU8DB7DOBvnFgrwF4r1YRsOdWgqJjlP1Ub0WDEtZsS+6dadEFD1cdVsIqAArQNqM7VGAKIw
Wr6d2rzbDNK4gAWtc9UUbqzcuHE5tvF4NSmpSZa+PpdrzfNxegvFBIXwvTLRMWn6OoD00gREe6Di
/mzo8eeBYCDqYG1/lIfW8I9jEHmZF6kmDeIO+S2u/bBRRdtcm6KRTwA+DGL34ZpDQaF7xcoHIGQu
muouj2/+kaoO3YJyfYuE1f8jdtzh20y+TgU+G7tNIC9+HFHp+IBtR0CMmB0Xs6xAXszcJoxPoWdD
7shKxZBvET5afo1eRKgRzSteJhsXeXuuxFxhXsUe/6MEdja2X1IXO4CxJgpx0JhOWF7iUF2QgxNS
5tiU8RArkTovgHPcSr/a8ZQPP8Brt9youYDNTRGf28vnExqXPFfkJSXR0gExip8hQAkCHgaK+jbz
P6jORsMh6RGEMK/eP6uWTNAIbWiQEmogoez4DQuoPt0VjG6A8b1Guqt9ZKgjDlhvj/hazN59QQUC
vnTziUJdxpCMTvWfoIzHvvurvV0CcK3BOsVAxgkUjY8+JVW/D/fFSOyIUF6X2l/1wnTXVJQ8nJpm
W4HhYVh+/eX5N9DTdR0Mw/vJfw/q6jK148qyoFvw0+OIjKq8F48lVlAkUrvQBFbIjYIVlbBopcPj
M/H+qcOcPZ7ZqamCKGFgk45+iz+zSt1luUvEJFPuw3Kfkh1rJy8p3C4B3fYduXGLUrccA0HL3L+I
qhLEODtCn/gx9D/pebXAR6r5oT1vMXsrwu1tVgWZxkGWIWPHvev3y2SdfRvQgzorh+X8B34QuobW
gKxN3VfjGoLrz2Lx3ACNoqg91Igbp0eMuOuTTcCGti0/k6RV/4F5s6NtwcE0tw2RuDSq5v94tEqb
rC1EO05Z87b3XR15JT5uVG+bbZu8QlnixXxv9ebVdra1vsHBKYIT+ShL22CRP62qi6g7MpKeCp2E
OAsEkpFLkmmWLYD3ob1gJd/z174J65nYM78WEiw6HtypyP7BXIpe6i1UG+5iJiBt4ornYEbYz3a6
D0y7vVjz+qYS1WXeKfAGl//D4iIfHnl8iCCo7It1tG1hpgaRbd+cHtUgN0IMSr4RZWg7xRPAYdhc
9lrC9UCb92CrC0dGeckcGnWbsK9XWGLhs57//opN2MyDAHWCw2z1do46sL+RL22jp8imx6F6jXo2
a/wPApY1atCVzJIrX89pxqO/IUghxt2aYvmQGSAekGql7lVx//CITjk0TiQ2FYDqPXf92350KObm
uGRyWiiSfmzW/7r2aRUmyyJKJOlSQqBaxCN9KSmVHVCfBJpVDzMmr/lIBCCjPuHUigxqQFx1hb+G
0XM5Qrnub8R50rqQwS1So2FStBL31bldR9MPEsvUf9W0TqK5RtK9Z1GQGrTVU/hiNqNaHOyMIPFP
5HNUDs4Cv3syAfATJirPmTOdQwAaDYNT/4ndqirCj3FfINwS86AkhX3q0naI+aNEcyB8jhf2kTnl
KR65HeRhrNprHl6tXk0SzHzJs6XJSneCqUPcvrNK2lTR5tds8uB3OaiGoo3E+Txc60ItqtOOUYkb
YD5PNytIap7SzUMw8veTd5Fue2IH3Axsw5h5xAz5UXt3KKNurYScqU5rQOxuKmU++1sZn8UFc7yw
Aeh2jUC8XdqwTql6WeV6eXgBEhM/zsbVgtoOHm3KVS+RKP9nJSPMHxTkw0IR1mY+ZUgTfXcmry8w
8pStiLrxQROjDtWDJ/il9F6k1TVFasIKFrA2HvVntnwXreJtGX4oA8erS4tcK2kI0RU/LMD7gyX3
rQ0joC9letGfFRqAstKE7JR7QSSMHs1FxO5/QHPhey1JgY/cdFMbEqeWPmsZP5qunJuVRqEkjtqL
sthlbbY5TwZsxSzTsh6sVbMOepW0Fi4yVHkJrUU0tRlqgsaC5zL4Yqlt58jGRMSaKtQHxOanTWbc
h7Rkfnvx2BmNabBrQC8RuXW+LTpc+GIccseVmqeAL8TW7c6F5ZPPQlwZCVOH7eOTWrQFOxRuUf+D
3paFnJcf2Cjnyyw1RjMhKiM3Eh/w2kP3oX2SKc+Yf/F0XDT3BoYg7MwDIYbcuLIXH/GlpOB7APT6
SZkmrnUUXHE4oCRgNojf6+pekWdAOg6ntvjNbb1QPjudbDZobDah7eTlyrK88ILL9LKgXi687XOe
AD3A3h7+7gYm903HMmWSgvjfgQowSD8pvc7oin/88ql/H+d5DIOny1hQaxOrr7eB5km+b5Ss2FGh
ue66aQ64QzcM+UrCSEsgG1Gvr5Sf/rY3oXMZ8Ny2wPDc+hqF8RsM1RewE2J7zf8Xj5e+yN1vNHSp
l8f1PC0kRZGMqrPrrFG5vq7mSlMcK7ko4U7knQTNcGa4RIEiE8w2z78l1GKzjPhS3eSp/82WlKjH
W3HVDgtfXEfNRc/mv3DPAgLVmmSkIb5Cn03RxAyM2cqX2YGhR6XztsuMDbqxRkpuAwJ778eS6WrY
PZGdSYqG+LdfSOBjKVlglF3UWNkGtYn1Gg2GPkC3JSVSwByTphMIrvX+0fwPsV5RRUVJcaXwzbgI
1q2boCFFYenYus0N/uTWAiiPUw3pSgidhymTut2kpEERyynOSeJz9X/tpd/G0H1JBnhLudrCl87W
i95QNvi81rKeCfRnWXvDQ5ccEK2Xh2Hh2+kF8nuEXNfqPHX4uYx3rcqzAGBjG7ahPGjoym8+bNCU
ra0i5ZONWcEgxOfNtK0rypQA4agEdvzlTaLqKSvG4LKuTJStZ1KcnnAnV8k1FnzcurCvJU+0OFVY
ykGs9zu2wqf2oLns46wmkiD1QivEySatWQT0kHhKkbBXpj4XVnoWqOjQ8mxT6hAYN8amiCN+ve5J
s9z3XmDuq/6OH25KKo907+O2tS3p3P6oVRfhOf/qcwUrFFOA1VdI+BIKiYYaqEoxO8RcMeEP+dza
/F33xURk4FGp2XMHIiHMD22SXNKLH7yxyZLIHrKcjPwRfJfbnXV+n1JIS2uZVJZ7VlrQhVtokJTi
xjlAqbPXbmRdHc+LMO8Y0RZYAwKUuXdlCov0CRysLmDPskcouvNNVSX0rPIaonIvXtwCNu+fTloZ
CXV4Ckmu+hwzxyDrRWXAm6PtsvrEQkhJ0USfTDKE9kpyBstv9BsEZNQYQROCNsPdTIKp5jtNixac
CL2i0pxTfi4me2WA+JCXIkqE7e3lFHcQzH1BairdIwcS2mpYR6bEwNogzobwEf5zALFdscxceNIT
PucQ+EtfvW4ocnNHNBK/9jrL7y0rM5hWTc5STgJDWU4gLvNtk7OCw4NoT8jLKZYKHn6K1JKDKUlu
eUDFVRWePgr0Q6RF2JUsAf9oFlPXtjPSMbwmNwu0DyaVvj7jxnbHW/KHqtkH4Iho+Zq+vSieORLX
YZ3fVGiw0Ivkqpj186MHW8ckvSJEp3PjuH3PYrzI+yM9aRg7HAYQ25rbp7DgjQmjgN3ZCOhipvny
8COUch04EdhKD4Ovhwuj4X780TPHyCKgJLJ6EniClQehvJ7emu5PMmnPij3New/54ug9DGHE/6w9
XtfN1QG8KkB2EmI/k4JYl+v0qeUtdvN1zx4HnPXtecxR7RxxK269IH54wq5fRptaGGO1M/VuipOY
Bx3arbZPMluFRN3d1E2wwsonD9MMXaZo4oCMb5rqYAQ0rleWq2zYudAitl7Pc+QmlJ5vZpS/Ibm7
jv77pMNlsrefuMfukLR8o/0o/Iv319IUrQobDm9DCqpfLaxJNNUTZfskgaMBht4gyFrQMstAuKv5
BCiDFImIFGGKoMRPqzQJkOIkZBjXog36otiKpavkpomLg0Qup1qAdZpFZJb/e64Ahli0zrl/Mxu7
+IN8U9OhiUgsgzLj+M9t8Fl6Xz1RzqCx8jWXpvR+zGQVqtxwLjYqBaArAoUSkVHBT9PU7sZAK8vH
qwDucCTjhmRKx6LsH92zVGMmf5J5XFt5DuVNNRLLAWwNPOJ0vS6m34wS0MFr7mJuU3WMhBKr9rH4
NYQpjSsGlj6szCoHKVK6TfY9Wg9e/FvuNGm+Lf2oTQul1bXilFHEjipwji9SKItaUqtLm6WlFerW
BR0VCwYTiZU15aD8VKg8yfIOvkkf1uRFxWSpUFIKeeAI0GCqWlhJ7PJ/VpzNQmduS9Qwv6dG/8eu
vjZvMjzgSHyqBUB5OXhPmIGcp+pLF2j+b8XoAuvExsfZ0TvdQ0VAs+J2ehcKR8n94jRTxANBjbrJ
KsTkD+ge0StLcYUx9eiCkQiWwDLp+PY5wMfsGhUOmguhIBfujSq+dLWbc3y5ztJCtRBWanbxPp3Z
BrNUKNdvxs82MJ1JsVUqbqjvaO3vWwVwljBdups5iJBUXwPE8gyOhoWESs18AvBpoHigQz3CRyV4
WeBXFXbB4CqwDTC6m9tyQp3iMNvaG71UL5iLhuJyjcwZ3cHaI47FsYdUXU0F2DNwopSqH7AT9S/v
47XbqM6cQiU9DvyKwVtl9c1PqWo0JREkoL/tl4tywFn/M8KYYwaUdPjko59mraVY5chwuolEJgLh
Qa4hLI87eS44fSyeLp8c9IrLSy2keHs2C4koPYpCPoRjVOMftJaO9o5occHpw3V/NLjSxg9VxMN2
KS+v4Lz0NltLNMT7aBmrwsZ3gvxvuHiVR+vOIXiIXQZZSEkGabXeaoOUCKKsswVkPDrH5hZw7yDb
Ncn4I1CZcp2FfUNH1xkJvoq6PSoWgDG3oq1LQkywsKBY3lhAZhKoat3NQJrFUExWSMzKa4BPsREJ
b8dZ29BrouqI4mLbHs85NwfqztIHdZ8lGkL96k2BiNAsUKTxRJ6Hs7xa3hiHrB2GulIDucR9TcL1
kRVHMZjeo4ySulef4Rn0F+1M79eIQMnKzN30UM1OxdPxn1lQ9s20ScGDd2ClFhWJ5CjY8FR9/P5H
Wr9ItVu/qPutt171wp7t/vgeqO5rmfdjJfPfnAR6by+ZqYthtpZKSryzktveu2uaXv+6B6SlMc+w
LeNkKoNKZyPpdQm52nyz5IsKJSnR0JJTejLzG5G16Sv6nmDA6FD1IM3/uZt8yzckdohahtZq9hTH
PIVtwMktBdtwK4L4jjmDqYrkDvmsCKafXBHfM8NzWn8qqRb3jWvVgD/ZQ3GQ6mtrkydv+GiXxr6F
imveZI6Q9VrN1QA1Rq3cwFSU2afb6d7JN7YvaaGmVVkFtJUCo8WBbX9zAFIIB5Ub+mDf2RsICt+2
how/00E9a0ushayLsl2Hi2imWo7uqACVASJ90d0oWQRirxiIu6Gzr7+1Wb8NdzMNNpqmtwOyBBpl
/elGEDVuQjgErY9c2VzAj/3SUaaDXJpcDuHVP97TC1VTndOPrUm82LSIk0a2voFajfjRUYhYXGuO
2T1N/AK3kFDJGGs2a1usNkfbilU1nFJEeNKplxbYzBJymEVbEW6XGVaXYj0RHjxA8MG44H67Qcj3
RB2GN9gAmlafpNKrQl29zjTjW0yNtKO1VLmChhLc9EjesLXbY4SE2RWm2s7M1WVMFpKMvKyKAXgG
jfI7ylfND6RoAgcXzNUf7MzLdYrhM2MGFlGqwo+yD6ck32w7U7NaN6c7DBRK767QdsAcksNc3Uuf
ZgAao50wS3coP7p2m5tghjerZP5/TdM6aMCPiCthl7FSxYxFcmUvQrlbHSHC4yEzkw7A/y+4Zf8m
oC+fBi96Rzy7yOtIv3h8Wkr09bXbGNQQx04zRVl6DTOZQ3MAdKFCGoKPd8yH55NG7MGzYQH1evcR
XQ3XxNI1y0+Fl2MC+OZsoAp6sO9+KdrGB8i4CQKM4qf9f2tJho6tMuZ8R2DTw2SgtOC1nU+Yk0bK
jS/4/r/Qpfc1o61PORHi+0QgxqRpx+e/AJsjtykxAT2SpUq8o3UiZZKDt1D7ILbOGy/nBXXRGxZn
ePt2HX1iHGYryMa4sGQM7JL9ZSl0hxYXRIw9Vx/37W40mA5ldwfYiDQCc+3btDj2NH0tK4tj2YEH
OZrT8331BKMQPbFfEDGM+nXBClaSiONe64J+P/OjQF+kC0vswUyFMB2rFYIzPay10BbbGzil70St
J/brjyZpKYXB6PVXC6QjN/XDM0O9dzMGrOkd28wRIUB6fMdwe0DsjdAijhO58f622IgviVHlRyNc
HX7GXIfnVBcZQFqI137dBJk/jBO+eXGA0Ss2GxHqkWhq69rEB/K1rsg88TPWUxY02nHWFe/mf6vF
XEsGbIBS8v4coR9AbkMrg8gX8EGH/yz1LuZOJbXFFCGsjfdqijYwvPUfAo6CXEBbp6qJOTzG7uZB
zISMRVK2nZAICiE9QJ/T8ylTcjQsJmV5IyXNvhQl3gxoNuBgyKLC6d0TDpIDI+NLYmmGYaKd3maI
P8XKdcZhnyxOj+C2YH3wCrjp5uMgNC9m507RpUQLJ120KE7BfmQDCQ+MeJ/Rzk2Z8696tTFH3pk8
i34AVE+ksxP8gphYU8KF+0WJvfWx5Y6+deV513Dotrl8JAlvJ6yuWsqeBvtyWH8qob8jTc6qV2iR
t6cbyG3bYcYMogXqVWHMaxY4LjNbaAs0Z9mQG0cW5/6Ha6y8BH4lUHzVdog3Q8A0TqPd9M9we5hu
/hqKoERfXY1TnpE4dSMGJJza2uN7JQEXBKMAMvBZrR2iRta7LVW6mAfy2FJC+ZZ8AtOX7CQi9M00
C+PJSBG/44Ejb6xb+bm87eg8lCZXKiYeghwFriw7Xkzg0NzKUexYKXjhpDDIGe5B93NeN8NiODxp
ZE9o0Nqex4msG54QTtxFL8KwCgRZAMckzbmhsY24Fq+wWcLztSzbLFV7D2rKfPxY5l5nUoTXx94U
ZFnIitR1oPn5GagumAMF8foBY7OcqSUg7EUENi2sk4XpehVIETMeyHCQdDM0YXG58c1U1JG/KvD4
/lSx0EV2y+l7iotiWM2eueakGXLCOwfb/leBm5ING4I+NPHQ7aHmmPMIYiCmpJi/TkATg+3ioXn+
QInrx67thVDvlG3HkDIZBxU7TK0NP4h3ycmBcZ99S+DuSDSXZU5mz/DsYSzb33CjAl3Chx9gzIFu
WIZZ8uOh3ssL8Oerv+P/sd4zRuloqS+oYgJVKi8WuVMTmDjSq7ENeXZx0Tx4TjmknO6CjMDq4/MD
B68nYY6/XKt5tqNBIJ/x2Sq0kg5xIB/+F8riJfTrLiLivQVba3Lth9Ngxt579hRRclYRt+0=
`protect end_protected
