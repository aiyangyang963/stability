
module issp_dat_abs (
	source_clk,
	source,
	source_ena);	

	input		source_clk;
	output	[15:0]	source;
	input		source_ena;
endmodule
