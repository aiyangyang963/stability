-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fjU5645rESMbEK4pOtv/x3lHJb5Fv9YG2Bd92c4Bzttj/LlBgl+eoKmfgQcuHaz2D57TQdoTJhVY
Zhgx4OxBA0oe+7BeBZRi0/5CzUhbDHZEIeUzZOAOLPqVgnMY3v61CHH/k87BqRY1eRDTRLB1zOE5
12OyY/eiwaXVT0DHDiMTlARe85dI92n1/0BCCKQrp8G3tHXDyUPKBfWpVVrmAyQXGR8qoCkyVBIN
DNLVgGWILu4ggFbtnIudFoNGnXChqxgyHlE0Cw5f1Gq6Xd18GfCkOPju3w1/Yf9RuH7SEaQoYQxb
5cxuN01S/Rk7voqFhUAJlfVIkfJGcMGxgrQPRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
WCzqecxCAx9cJLf3GsB5DSchswz5i5dTAn3pS6sYTnSzC+lRgftUOgkbmN2kWbV5hIACWMyH0XZI
OxnCYxYHqWLtMJiROQ+OR48QCGce1defx8Q/EgqKAvr/7igzzTvMM2pELfoDT0UyVzwWMBnVRurr
0wVHc6IPGVePOnkv91oOtIEQT1b0X4Om7OK9VgowN2mR8i2fDdRAziTbz8XcSubsK36DMdQq8nE/
AtuiOvQ7eAAppR3BGRrqZncGnilLbyEmsONdQQwXUUU/9XL3ZkmB1MlnvNgPwwoHk4UP9P5M3eKF
HTjNcRnbfO96PlBanT/G3OIVjNKNygH283QGZoWbROSLcl5IOdjJAX8+cyFz6NtULYL9Bvvo9cX4
FnwS8/JfnEwBnxLfnCRGRae15sI2k0+FNYeylEnnCvByoFcyYXkmtGjSZWsYFrbvYPNNT7MutCW0
ivRgdKwfrQiHlsQE9mguC63MnYnIE8jIqeXbF/4Zt7DRTkK8EMHoPfn/A88BiJ7MnQF0WVwbejQ7
UWLbVFt4qKI8gb4+rU7oEt1SwuFrKqTcGsPLZLcy25k/yWSLUDHZmSww5sG8YaByp5nD/IT9kphH
VH9695opeISgYOm2+Grz6SxVym92+XnN7HWyJnAScYHUo/tDCFPnSqe0tvsGsfIz521fwNOWzaHs
ASM0uIIieyj2/PkMk47xIFmsHOHmerhMHqzkAcUE6in4DviGuhGBwB1m5m1Ir4Arfi0NesSyeoPM
rgig7Fd41yK2YJ35Gb/b7ayMuh5j6Tl85ONgsxaxPvYOo/XoJnXH8y0CaH0UwSmTiOvHG0+AcER+
zgB270C7Uq4YbrtrztWCHbBd9RVow4MYT00OaAQo1dU+YKHCPCGvDuJ8pKTewRGzW4s7cZcrk2D5
Z4IWqWYxYf1r4ikPpJ9SDUcG+IxE1rx5/VQ0cpWJGCcOYIavALUPyt0ehGtkGjDAnRxfYLw8qzfU
BtE/zmT318KWQItcKroXH3JKncl8YMfL2OmO0bF7nmaRO+Nr0gZLjMTKA1AbqDwp4460gZtd3l2e
Z96U7aUIHO1cGTaJLOKxr4Xp+UIqtHaWo01bYCLNbB44rETormcZGGrTGtmvubtS49DaOTiHEzvr
h0nhuAZjZ/amYpxbWODFLx+NcDS2FH9j2xnFL4phT1dOJ2M1QbiBg6eIS+4ArQ+xfr0U6aA0UhD9
d2m/zLZ+5nfBK+qW7AU+xjgtUyz5WM4Zf5N89DX1Co1G/2j6k/iwnLbvDVDVOQLJb8O5u7UWGA9W
VGP1Tz3A0RQi0X3wVPPVP34wHj1C1uwK0+N8b4BqohGzr+g6DfFlYnwhghzUVbDNN9Qiu6xVrZG/
/VQucc4gZu6osYVfcIYE0U7yixsGEyTlDQEO38aOY3K/8eDqvBo5erpSCpDQnblzBbep4gJ0t+kP
8YAHlKrb7HTg6ScAocj7wv7ep5jG83fHmDPFc4bjfpwQngmr7Cf8mSUT7uXKISlNu1FBFMivM/k1
LssaXNyHYWaEeeHYzQs3neppbc6TF3XsyhgmMJt6EU7vQiyQsS39J0mxNm3ASPCL6dJZ2smt26k6
SQeoODRnvsscYn5mfsph9Izxyo//mSm8OlbHQ/fNMIzOz1O/U0+0ZvqTRpIcQko66K7+21T9Sr0F
lv+8npi9L+hlDTpz09PyGNAuIVCITcUjlMhki9kodBUAbjS2375AvuL46vno1+EdqL3BJb0zzzaB
0hVZ5A7o++qSv1mmWCi27c3xQy37Sza7KaC/3FvE9Wu+FTTMPD4e+f19pNzmeGPmaywCzZP7QQr8
p/gSlKmqQ1LcYbgixN/IHLtlvhOaYx6uTpr+Rt+rbx6Lz5KqmTfCu8TgUhMYaxKljOj5DYFuyUII
8ahTGhL6OFcgr2qZ0+QaoNEG8NGHhJrUTsVUdGLEs4ECAmPMIQ4gi+RDaKGYsvwbO5lTfRi9gTiV
zzjFxkA7E6VkgfQ9ctuKrEWv3pH+lGOMtFf9EWW1Q3j/wyXbWm6PaIekjb9AnxXJiaJsUOW6Ys6l
3Egkm0H14y/0v9/gowHf4Fmt7rKLFUYSvYFAbvGyaSoVn7S393yX0Lb90Q15xa3gWOHOOZh4CdZZ
XeBw+2cnFQSxcyjOk1B+Pw7jL8XXJC4nUZpAFjYjzQ8v9A31xEqGDZhniUMBT/aL8UPQ9n4LTeGJ
yPEzZ8j4DpRHovdSBeF5F2SZMhmSOb7HXR25LkSsFvbK+eYV0yGEkCpVQJP4LjW59FH6t3BZWOvB
Xg+A6YGCgi/TALjVkxtybqr9tNm5h81V19CTkd3T+9NnMWJCKp021ptXxxsLJnmu+MdKnG4p+TLC
CtBpZArNqFEOdq3tvkWxyVcyR242NZK8IM3SNncs1yip0NEN4Xu4r/fUizluLWAVgJmGeugXsV7S
a+HhCvjqK25tozLWvriFoL4KgooiPkbsgZDpAmSuIjarQ9UL84X0Abu9ENsYSIWIr5hBl0KcdkRQ
y0A8YbLpuwkp1lDC7diXAfyH/xqYZh8QiWV6uh2QkYQDAm4hzkPQzxrAoeF8QBr/wwyD7vkLx6hG
9kCpD3rgUQqyNXViNynVwN+yA7JtPH/wozTIhm67M/b+loZWph9SlWNT7pYCuhAGlG4grQSydjK1
b2Wb44zNNPGlUKsXpTI+MAa0SXi+ihLBlFPEfrqwvDi27C7jZQ5U6IxKVHsHFRbNyqn7a5AiFMdT
hc/Dd/yzMLk/ymxrFczHHscATMfAlDNWmONyoJr9yXu0ukomgHkREbXosMt+ue2ut3pnLnwiZJrH
aUqssrrSnCyrxAYPpFbUdlUcxTnJXmNpbWQrhDvqCbHDmJpjxZKZyXSXvHSLGZSFac3RXcEfnGsx
3tvvSH+isXffeShM1xJm9959l/2WLMSUwoCZiopZDTB/BPWNxPG1OAw8jS0zdWXldJ61fwya2Wew
A/PYXqz5nwl8RjpnH2CCS2cIM8XXatc7DZUW2DgFhrRvX5LmABk9F6VWHMXZYmSSEKqUZcsHtKum
zUA2OEc3dG+Z1Y7nEK2bu4mW2bXDnyZmvjt7fDRKg/m75oosY7IUF8aHGZil+nf6MPaSZCbeYB9t
dvKps1T7qImjTiXzqwmHGJ3/t9c8fvlgHwmwEcYavwL6H91TlI0BbJhR8dH4Imtzoko7/56nEpaM
/uZvDaPx1GjsjfdhkbERZa1K5VWDXgPe+5uIgSdUIfOL6YufUw9S6thbe+gaYpv++6blJgTWcJCP
RD6ya1LJQWzFEfLkd6MfqMtePDuBlpGM9htKcWNRVruY7OhJTcijtrJatUTWTQT9SmBisej9A4i1
8lRqhzHFa7En1JL1hjyWQ7fYff2v5Gxmd9TGo8RudHZM+hK/8x9kooY1HDCqRT5/yDFwnUrCsUrd
1Dpv4a7rQhAgoyNyqhyz6+AS18WIvlJGI+ua9zq4B+90pFlC4dRVC+WCMQJ0uyHBtHxTFxsC2J+y
386PiJ4k4+LvUtQwi8xxHMmksNLoNO1NGvFsXbz9R2mFwrhbF/bv/VE03Wnw78cVlGfC4ubDv2MV
Kp5DMEIIPa94RT8t8cmQcTwTBxxbUDVXNbwUZWuAbLozGWSX01EadpJvJIwLBRgWIpvsH2jGVkh2
R5MzIvGIFVXJEXPsyIm4/opJRCjoi+MjyaqCbdvQbTMktDxldHKZtjqkHjEN0AB5rewQW4L67OnM
1k/1aRI5qyF0f2lmldsmAmGnuYUPDdjtOTjf0JVQTVKiiPyvHBMERrhQYanmH+1HDa5owtKgqerG
XiY9Wk/PTRBkioLoShC+0GTfQfre0dRAiLuwxQ+cJOp6MHHmexbhQnb7GoEuwaK+eVd4D8xeGGNt
XILUM8LI21YPRWS/ECwZsOnRW6vMPam96tKTwzl900wjuTlG7G3X+UeZx5dyls0bhFt9feFx6RQ5
0GSqh09Gj/H6lNCkYZnqNyXpxPVuYUsPOeN+HwgOaYRFk2brV/Qz/82z8/7Q6y7CQClxCNhj6Zh0
NaHr1z/Coja6EWcZ11zjAY3aT11gg2qOQU5HJ7sLiP5foB71Ppy/peNV4PiaiJT2IfLPhtCBKE7i
1dRNQdi92ZKKJoeXkV4u1Ri/zIKoXLpuI/T133irETtwiGII6vR3+Lp3bWQxwBMXQ1QhWmTMe+5r
a+Q++k2MYW7ZnEIFDHAayWKXR1PPNb0iHJZn2jsN3x0OcVsMX5SAZGB26Nc9uhvcPfgYNJtG08Av
J2q3u9q1sRS5nXQpK4CtMqY44IwViBC4wlOFn8dRut7/0tWLnsr6CU6coih5TnU9ewcnxpn0yUvO
Kp6HdDYj/UZKJeCLsL9A/X1gJ+LoZ79N+qARBuBhBMd0hfmYIUG/YEb0WtDFYdSsie7k2bp05sdg
wUJvuIwPH33mp5cvaK1jsjjkyJY+eTYL+FqbBPqsoK6w5b5JtpdtoU/KQFBF7LV0S6X6ZASTN7FO
yUiOw3Nc8rJFik43RSvqb6i0EolNRbA1fQ3tPelAy4E3sxE0MfwmM6+DznbnqQhn7g+PyYcWgQ36
Uh27oLQ8Z+2722JHHjdYp+qkKhFvmUZ8GYAnNCF1CO9Pg/j9IP0rf5AGIrCaczh04qyVQ5JeZhvG
fma3Gz5txliG5NLY8fKERy2H7hju/HwoMriqY0SHXQF7yu+so3PDVC75jewqH+UghFoK4rB5hT1M
ZSytjykTcdjDVK+xvHfcirDER5wPBWE38v/d1GOMb7EVaQdT8SHUetvhb/eBlvDsesY8grLRMUhW
2i5zmG2rJTZ9+5G+c+2fJrVkHpegh68aLzgQDkk6MFmQytS//ab31gFjFOYEUvzaKp2DVr/Xa/8O
61pr5JAGDoO5p5mxN79SlgtytQgs/ua932LW5aI/G1sCYMPIFGBE+fpfDDc+6iAnjUSphaJRPrnd
gLwhMAYuSBOTzbKhN7ftVvTGJ9jUMpmby+KOS0OM168Ak4gi+sXft9q4A87lZHuogJrQpRSp/+aI
6Ebin9m3uL3QuMYc3tz3EQ2RtMHtZc+gVDPXR4Ev4J/6ycD0AZGGqMZw/6vKp3JD65sWJ4uvcVx1
0tmYZU5uLFyq65vZfycX0jTwbPvcExTJ5U1L5g25Bhi4wMADbaQndw6gux7JJ7mCzdKTzZADA5qv
dLy/lBlP/2O8fW7w1wTFefwFi+8zYCVixZ9zx0CR8bYFRJWRRgPiZqRmUeSVuIU0mYqwXN4yCKc6
gQn1doswuB4zwEP0Da9acFq8U7elKBFOsneCOI/uB/OSMDWAjDsm9f652MlpZ3ewEaSpsX+1pYI0
hWZJ697EDoNxywl9fTp1HV2Lb6OUtqRqpdjq0jodvWCPjGBAXOiZnNzj7KVs5UhPyPmUJgUKoIAa
HrNWAdTN0FyEzb8QPQf4I/yiCAQIOHS+HDK/Ftpv752jPMxQd1UBVdlH38zOxaBfykZpxTfjKMFJ
A2SU+YVs7CI8qSsTbn7A9Erj5XpntolQ2eXC1jfb78Le29Pd6f+wIcsKHZoDc9pAKRPrXbivL9bX
hrUt9hudO8hrHyVwhNuM+l4LPv5nmbc7Bl2ojmFhYQf3cnP2tCseHf0bnNxl+wSOvMY8rQapjMiY
eYdbFkeQn5/c3qRflPa1N83h3aBjrkH8C0ZwB7Ihdx53sgQmuizVa7sSoEQnu2NuHSDYgEcW83zt
XCo4RyDBWzDabmLGEI8oEwsrRUGaXCEOvtDd4tb2x4trJd/WBqaxUKfwY9/32rOmt0Uux9cFDuX5
hb3/1B4TwYnk/al43+zayNd6SGSu7amecoSdvK/lfEVeTTpC4Tz/k1mAfHVOGq0QAWvncP7aCgcK
4faG3kNlAnM9UXYmkde/KlxnTmWqI8Lcg4qNP74URSnur1L0hQxzGkfjG9wIYpZkNegk/rJWaEcX
x+2XTfXec/W4+OeUBAz4fhj9ShwjNP/SB72nVee1lmdBt8FE36S7SSPjVsakbkRXwx0bArBczBWa
aS8V6xvidxO/UwPBDjd6IJ0KCi2XEnw7RdtT+ImiCOQ6E7P/3N9mdtS7AULUiaO/18Lc0yF6x/GT
g4L+O5yPAAXr+Tv1MMEZTvxZnjTnDyC/orgaUg3L+sbtBh1AxPpmDKrW3ywoYGhJGLwNe6hZa9Vk
lMWTDpMkHsuzwtsbg1xcgM4/OWbt48jMr5SSyS82uGyxUDe3tNk3V/Re4vFRwXoZqzlEueGB0Gpf
Q8UyxQI38RGaxc7KGTGaBpEwrdZkfcmcYhEUlt4GZ2Kf+GtfzC0R95jzmhgIk5Vjw1OQHh/jf544
4PtQqL1KLc/iDR1xPzptFU6s+aTulMHu30FWmPwkX58UAzVJOVlaABf9SvrTldYRNgSdmulNLDMS
6IEbTJOOOg0Ce9amGoOJC8C1BejNa5MRqxR2aYw/rmA8Q/8STYIND7Oqx15brjgUoLqOwehRFstt
mpPdYO5tkgtlDm1suBHSXvMD5goRpHK6y6Xsbqud6veq4lOKWn0YJ1osbtnlvtw2pdopfiv1TORv
zsz2ks89RZH3jEyahtW0eWTWk5UK2sT89wXTcJEpeYVEDjhdjNkaspvusPlKzlqXvEIWhA38/uKp
0iUAy+AgvsaxCR+TVHCIzoElGjZ8ebPs6TGscgUKUNY7mMFe/yrWuHKHOkjN6GRfZ4IQMxB6CbgG
g7p2UXS2jjIXyjz2xBjuh4TKx0QMfgd0yEaSlKpWsP6hzV8+bTu9qlColns7iLqXWBAQ6QU4uVlB
zIivuAGaUNg1/3dgDeZ4OFBEsYn6SgIoE4N0dU8PLLzp6/u23bLGxdJs5n1HCe2JU9g4XIu5Ed2u
50Wtz8CGxoi2Y+PYfal+gx4vb2jEDInZ4CgLMsfKBeDSp3iD0QfcVsxIn/oArWfMB0K+fUoCyHzy
gR072PrqNE4uf36DhqKIcdLIa6Kvdrg9VUCuyPomJrVUuoGuZhUIVwlBH9lda78qA5jFAd7FplQx
/0VaIThv5gsmLI+3np3A+SdHLAjLSR6QJfzXVMSw/uxfDjXfvMHSItK6m2/v2FNKI//paQLLFh9l
a18e83yuxiR0tXB8OvP1NJUHytyzPVXWnt+uOWcv6Za9ANxAEVIbljqJg6sXodCkEtsOTyjsnPqk
2pVnKUmZ+8yMR2Mimyyszl/HLGOYnU8zQvioznAVR6BSQ+PedFTfeSHXEE8DaohNCdmgacgH7Xny
/RT/vIOQVewDguVgrQJZ9E+2s0gjHTlum8GQLM/aUvUbf4CjzeA3PqpzS0soT6OTSqbEbefLLVP6
CGfq4gMII1R0k3N/7+wlhCEmXHpx06NhRbNgg/nkx3IPogyFRDXQ75dzTp13bxnJbGAndPbU/LX3
zgxhovd8HPWVWx2uhSWZn4w9RrV9k4GyUwLdQBblwpETHEnDCEK3bUwyqO//fWASIQfn+hJQCvUY
qtknodVWszdcaMvXuex+s1OVNtkUkMGJgPSOA0pS7/vN9Dess1hKubb2tp27Z9h6yLVRt2FwEskt
bJ6o+wYq5V/2TOConrBkcq3gbfanrthR8zFqjGTjZLy90pw8A8FdhDzVS/xP8r79RtwJomU7b+/R
SWDuuDN28Yoax77jivJZvJ96gF5scmK4hFZJ0wr7iu9x4Iv3otatb2+95ftV/Lt1YpBxtzVjoP+W
cAar0mfHz0f9s8iml1mRY0sEQbs5HwX2OngRTG9Oq0WzElNtIuSSeNZUNaTR7RwByBhQCyKwITLx
Eyz4IA4kQwdfZqHHjMj0xVkIiik2uER///0bb8jf2eQmK1U9bN0SIwjKaCtli8PB339JEmIs1lRd
CaNoDe8oDNWzF2xGuMIMlZ0kmh8l0T203EQ42Bvsty+WWfRTicrmT5tTbEjtBNGu1iO28jYZDw50
b2YktaD8lVaJY4qDZ0OCprQflACsiz+hLlNa2DibG8z1bcWWUPKQOkQAZfhmleQpFNiMohQKMiGv
e8DYkLuN5YCWUg3cs7QdBC6tGA1oE9fe2LTJbWeA4JxBQvkR5KrjvB/dXgbl9+jBwIldDK03EfaJ
v6IlgttH3xLICKzDH2mYBDuht2GBngVr+mzJ50TL891AbHyFoyfBVkoeubBiTYlr6vpOB/FxCwxh
bQ2gbwv/lCg9ZyOg/3YYQv3z1kCLXw6mDvNm26O5Sgaojnq/3bA/p/qs12A4Y80CspWIa670MBmv
iTYTqxD5WtXcvvFGpyhQPsY/gDck4w5eNDHPy2jVe7pe/Zt4sfXtI+sBSlQ8zNRTQSaKppmkj3cC
ItZwdgy7irNkxEXTKzM+6KCiMP2UNmfP06ATbxKHi8/ZJ/cwjK47oPYi+zvB+WoE2AN/6Htau5tc
IVeQVbikiIjwfPhLHjQceOjvUMee3m3n81Z0bmaf4Ft6JRSmmJEdfZz+xovsXt/7FDhH0hpl9d0X
qARdkLw3TpMHJ9/O8TPHiE9M/AEuHpAOmsh3ZgMozZx0hHhiWW6Jd6gt8N0pAnj3LtaSG5BnB1sW
QhWOLeJ8M8W8bGguU3VABr3rOZmeiME7ySfmAma1L/1k108dG9Qa3ylc5XfqgTV/n1jf/uMhERdS
phu1HGw/KYhalReRIfKiMMZvPAHORUfdmaZByOBkZjOwYLTuHJxdkD3kMd7SlXPtH5u3GbXmUQHj
MrjudtLDRT/LJ8l8jrS8KsFX9fQ2mAAjYcEkSUwUeUjH2NWo8ZrgagB3c+7aK8kLfGxJg44mSvqE
nurmn5iVN5jgTV/vl3DhOMMRFN38GdjzoxVlxOFaNQ5gN7vBvgXuRdwv8I3YE8qlfzZ/KuAi4+SP
rC2YkFBP/XjOfoXVC4XuvR8MyDQE4dWRJheMknWwctovMu3PRdn3TNnCuv1mrQ+KWMaQ9q5BUCGw
wCaMZvKaJ/dk9U0H+M3DoowTECiN7a6rbtyHCjCuMYQKZj2PKbP615hKQ/Up0MZgrLz71HGCXw2v
jPZcxAvELJbDHdlXMQHjKHEvTWp63pRPs8K/I5/C9b1xqYSok7xgsfGHDR5Q3SPXJ/wPp0TV1dBp
y0staZbwmiGCEkeBNYF8xAoyLvvR+m3cRQcCbd4eSSbd/V7J9ybmMNYwV5ZFFZrCi6CbF8fjesTI
8mZ5nNfZm4ig+OkfPlAHbQ6QHc2gc8XpFl4oBgxWbXah4bq+UU5Ey5JLmoGngsez3ivCWvhblOHI
Lx+9TriZ7SNcPxlI4DhTPS9tyl142OYmEXHL3d/1/cqpOQnbW4PoCc5XCEOWICeuwZreML3mOxQQ
kJg2hc6yt/jfaTiEMzFSi7eUPjtJ2Y1atjbzjmkfTq1T4K2Y+44ng6LEDgPb0PpqtLcLKOC+Yx57
NJPIAzQhJ6IEGaAWHDQIL8Y+j4+Dw94ATuDSVL3Zg2rMaPJaLlKKly/ce/visH17ZZ9/wyGjXEvR
5cLkFzHRYliwu1NMHW/vLRFqbBzUoxlkzCMshE5O4VzZkhMECtLe68viR6oEv7RyJurv/gBnEt2S
6AonMyPKSl78WxV4I8inKylNW6x6ZBKPBCUcvG5VGBvYmmc+R0FCHJeGg/ey3TmjrgYHkr5UXVZB
gy4p5nnGbEQhk1HTG5UHqlcJ0/SeJZFjNh9nzx3ECl067V39PJVtjohss6yudrWy73QK5U/mmXI5
11PPxHnyYDacACwecQzD9IKY2yrkiDlwo6yiNZr+K1w0F1U74SgWtNSIsH/bqF5bJ8EOH9LoJMyR
VUVl4RSpPbYQwFhFb/dllA2OH//D/OMBMjRT+28pGo4EanLYnMP6EtpQ0crMDHAX8/87X4w6YDAo
hlBlUprpR8rLXqS2uzWBfKHFpMuGP+UVttLL7V+DfCyPHpvAP/XzD0pttonAO0qJWSwODLlDP1TF
jhQis289Rod0Cq5bD61LZcxMjKSMl2GuhIVjWhofVzAKNwnGdz3jX6ni6DNlYn33ov1LT+RGwPF6
+T6PVydvux/z5SRZYUjkUPJ/ewtR+f4+4br70WpOvzQUgi4+sSoJ/nUk6o2mdftEbPYgKs5kfRbc
/Yk6FaFw8rC+wSuvhIgDct/dkZulZzQxxvhHK6aJrHQw9122s1HnySfVuR6bAR8Pmmy/GfUjns6J
/KFFIy/VoWpIDv9avaCy7GCvIXP7h1GeNj9HHODK/sncoz+Q4I6MTOMW3p8Rn32tXL3skSSBrKpt
MLUTY81eZSAGB1d+cSuY/Nz60R6D2dLOQ21YgaVeg54ntQ7oygkBQ9YSHLBGtiOWbtx3hWquM2GM
5fMkjn2cXM5s0euJgUTlV9MiAo7UzQHwH/qhe61Y+8Aaab0K6Gne5LYK/aR1PVWpVs/Mqtgm87TV
BTSr6zQoE8Z15GFuEls0rqdhrr2cf9IbpPG8eTPqgoXrtV0V33BiFFSTdTofGqXmsoB41dHdjBdW
xVX+XDLYOsVaiJUWJLxHyDKppv/J/BQRJ3gy4hSXqgShEUfYG5XkNHHRUJJA0lfRygEKD18c24xO
+vQuHHxU/kP2sDpmzQ5bdO3m4tyCKDd82ddnAMDFC5iI81g9O1em1bOn9hYxiyu5ABt/gw54zcYc
O7oSf9BMU6fo0gSt9ObcWYUMktJSgLSMqySP04S3xk++mX+92yveaxR9J4WhKT3fdCpS3asK7tPJ
quqX4lP4wdxcZEfUFjy+rGTaZh576EdN8iEzo/sWx67geTShM4jLvawUzzIOqomdeZUwKcLzUqC5
NRUFMFF/yVJx0VBfuaKpDWCSxw3Zc5WT+oIPoH9GK+tsiKgIAAQqIjb6mPTAK/pxUkUIp3ZmeCVA
Ca1uQymDmhVqGEzycbApW3RvUzfQW0rBfdOq4dU3+MFfQMQGRpstSGwm5oyObNpJKoOftuJqXEkB
Wlz21Xbs88ZAr8oEPCsrbOvfiaTc3ov0n0WMdFNgzhXoeu6RXMRRdYI07AC4BciTpSJsc43WZi2z
EaSSgsajxWzbLjVXUsDVThKEAd0cWXrkV5WO9+Mhhfxo+1xOTHxyE+IaIobp3n+8yPso7FlOQ9qr
xmjS5yBtoo6ChZH5YAPFS3pT3/NI0NfVaNRyV/5kXOFw43Pa+gqGh7R4Vyroi61p0UUlif8OkhWB
RyR7MHojd/TwVUMkVjTIvHndjxuwTugxXBpJt74ZonoR5VoJ9l8G3yCqHna8YQmwSLzeMQIYHYBt
fWbywJDizjMyfbihO1xZy2PZYqQImrUtzckRZiHFrdWyx6jSfYgYpppIL/hXVH4R+1ThkearJc8B
CrC6vamBzqlvDrsGbLcQaumGoX6FvkSDbRRC1/D2pofWJz6oIQmjvQVupaAK5/wP/+r2fk1hjORS
6sZQOJrOttFIHja/DTuFNhL1KrX9EEJT3F6JMqRFK/TABQpzVtT9LnxPz1IbjJ/In9BiT9F4bfpm
o07yY5l5HQLca/U8Bu+Opx4G4D9u/uV1t6NXScnDAPwGfIbWOaKBIofzOIkWdfN5WG2A7ssH/APE
epSN6eRmALtZQjN6dgtBPD3O2smSOQqgX4oCItcAhHxPgW6Ow11riMteSbVSitAO6a7SuEoEDAKj
2yFr9OV9/Z9DI78JwIFZRV4wpLuFyqZwW6G8jreEWILjZXtBfamzkqmy+XnQ/PO4mzPlgJFHnTyy
KhOPW/tW04HkcvQHLwJMi7g+fxhNt0Q9ysAT5Be7s3JHqngGdUzN3EQoF4d55X5Z/WaTn/H4ElRC
LEYJ0en5oAHzWqpG9XEpA8iXbWxGx+DrE5lxdUYixNYAQiVyPiYX+2dUWAFRcKwF9venhSIV7zbg
pP9WB2X19qyXcl7TK2S3cWqW8x/81nXmo9y+2mOSkZnLkk5EiU6RqYgfpgQvMuzwDPIvNRpNahlS
tWDEaAVu5sP1PGfKl4DLF7Fab5BhkRL8mDWqi7csWmzPSgJhIuwLkNaycyjEDVo/8jU5SA8RY/Co
9fCaAC1wiBQzISv3pz9WLlLhP/c6MT02rdAZKQZ8UNTLr3X1PQ7T/jLPTOCYZ+j74pJdDD76SZwJ
GhUkLOy2UCiuMJOM+lXYBl6DYXAz+ZwNOmf7LmPfDUsUqIMcDLQo2IWxEcIIX+gVLEEzoFrnzUBM
LShh/LrxloF7hOddNTCiT+Qy8fg37UlycDOKxuR37b9EcFCqp/frA0QK5TxEMieSEYOum/4EUHwp
8kzmT9ddFV0k8YcuUrxQ3SMJMzOXKpXQeB4P1L1gtbHrXn4E+1ZZYVC+9O5uuH/S/4a32e1S2UXc
mo4ja8aehqsoAUg7QHoNjSkoQiZ0Vf03AzoxW7y6mDGLPiMN/ZH4OmtR5arD4KRvbBFYtsb9YEkA
yHE9LuWjFys8Tnaeu5SJ1Dy9UEwpvWcf5DVKqw/IXY3g75SQZv7vNoClXN+JBrNztKXugzRvOdrB
X/T19wEf+Q72PPcrcTsBQ+5ps9hdTZY02Gyf516qrsqWm5uh6od5wnVlbZ6eS7tbshtn0GDdwyjY
8YYXFaAC8GIeVvDCVG30ekq2nLiK14jh221WHTBHhxH4PZCNWSJi9sH7Ny/299vNWI0OtJjDPL35
67Z+MQP8u4apnM9N94T+x6FqzjmjnbWDgPJpvEi0HkaD3AKCdl5s1ZiJzKDuXndLpRSIkIYnof+N
9RIbUzlsrllV30zpBJNoSYPW8Pc2g8Q/LrqKUSjDcvxDf3Hg1ExkqDPQp2RqiSkWZWYAwxlc3Gw7
R2raFXnYJJKqMo1Ygxrq7DEZzqsbT9f1OaByLDYAbqgPigykI1cYspY+vzMvWmdGoyr6MVBhHlAG
qWx7R77KrBiITl4M/SdckUBs8/8yH+xOUekmLKbkwWPAWVEoidjUldgGMtisD+2N/OXCyPuaEZIu
RYhXZCbGxASl2DIykd9DSBNbRFi4Do7RFBZUaKkT/PUIK6waT7NGoiGd3ZJ4xRUkBOeTjgWjWwQn
Cv4v6uZUgze6EBejMNq1YTHOqRJJoU2j6p04Bbxc2///QkTeqFY02mu9E0kyFhBtWjfSepJbx9yG
dL8J6UlL9LiJzybBPTm9la+PNCm7LZ9d8c7MwVKjRmiBRNd860GjFU4BDxffUhl6rnKT5+cQa6vo
q/Oo6yPH0BCEKw+t+Y/Fc48kiZt56oemHgM9i5bxcz0lktXN8WKUOmIMWPoa5zxCsmZWqlpUMi0k
M5A8i9FSgFn4LCDMeQ+72UwDPjh7/bRz+2Df6y0loB8fSVoTHrIhyThSNaD8ekRdMRuoXxSXYelt
zqHJN34E6md2zKI4YTsjhzlPyvog2/mSou3t/3KkF7NdUrPv/3I82mK2u18vJeakRqoc491NLL90
GfW6rOhbrNTJGT3sDkSsvSziK2Dd1J2yq/p/kyVppzUy+4BH+oM1/PUOdoVxmnL6de+RysORlhel
xVXTgBdPcy4ipCdQVceyyPnBunaoqr/moGGDupFs2/Jua4iIQqdKejbwl8leyef1A8rpbmtfqs/9
8iHJqu1pd+XuFVE8dmP9JvDF5lFIhzt/GPJCttYLHg6lSI64S7RlbRxhIMlBAYz5et5P7rgkMMg3
baXACJYknFCcHmqGJtMwJfHnjwM66XzuXGC/7HcMXGuMN+BinmTH8KyOhr0fvaMngCScOiWfMEj9
RjmL5fe1wJXrtT0tqZ2F+PRiRxqY76UJIQsWw7MbyR3VYqBJYjDaUS+ou04k6TgnHGSA68VZYVEM
tlELnS0c2YPaGMZ0tNpURTV9X0Do9aHT9Jhs77lv6RtZTc6rzVuxQ5W2FfsbLKIR9guGNWiGsA2R
xS4BKma87pRaSKT76NEuTrJRkJZeM5ItG+UsDeeAGTftVTXej6gkw+NDnRUJppac3AK14ZGVDB8V
Gs0VUTkAk13vW6nLzPuKVZc7FUkIMK/EBkRtbm6Ze7vqpV8V1oGnV4snrUpV08lN+R98CtO0InYV
sqsBhg+nIx/uiRwIfJtNfx5X8m8XcQeo4eJTTgRFcToXCkG3SwpXciTjxSV6l7GIm51dwoA9eCGr
pe1ZcqzQj99J5iFp7jBS/HM6oH7oysa07MAxlU3bK4VL1x7yRetebqcteZz1Cbzj1VdzI9dwuVWv
OOe4kGQrNPENpLVuxZVPaUmS8Ps1A0kdMf9YKeIlgx+CwxrNVLIZutlowYHof2M=
`protect end_protected
