// megafunction wizard: %FIR II v17.0%
// GENERATION: XML
// fir_2_10hz_nco.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module fir_2_10hz_nco (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [12:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [23:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_2_10hz_nco_0002 fir_2_10hz_nco_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="17.0" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="nsym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="50" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="0.00025" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
// Retrieval info: 	<generic name="speedGrade" value="medium" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="frac" />
// Retrieval info: 	<generic name="inputBitWidth" value="13" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="6.581512570846826E-5,2.3224682081490755E-5,2.1263915186864324E-5,1.348849582427647E-5,-1.884515654637653E-6,-2.6618803531164303E-5,-6.246339762583375E-5,-1.1093106149928644E-4,-1.732944801915437E-4,-2.5030970573425293E-4,-3.421740548219532E-4,-4.4828696991316974E-4,-5.673483829014003E-4,-6.971539696678519E-4,-8.346185786649585E-4,-9.75638278760016E-4,-0.0011156742693856359,-0.0012491375673562288,-0.0013702119467779994,-0.0014727171510457993,-0.0015505029587075114,-0.0015977213624864817,-0.0016091193538159132,-0.0015803587157279253,-0.001508324989117682,-0.0013913477305322886,-0.0012294170446693897,-0.0010243176948279142,-7.797284051775932E-4,-5.011202883906662E-4,-1.9567001436371356E-4,1.2790676555596292E-4,4.5975486864335835E-4,7.891962886787951E-4,0.0011051764013245702,0.0013968131970614195,0.0016538002528250217,0.0018670330755412579,0.0020289572421461344,0.0021340770181268454,0.0021791793406009674,0.002163664437830448,0.002089534653350711,0.0019614456687122583,0.0017864631954580545,0.001573855523020029,0.001334545435383916,0.0010807289509102702,8.251464460045099E-4,5.805459804832935E-4,3.5895180189982057E-4,1.710843644104898E-4,2.575004327809438E-5,-7.058848859742284E-5,-1.1422827810747549E-4,-1.0438119352329522E-4,-4.327772694523446E-5,6.400272104656324E-5,2.0973681239411235E-4,3.840607241727412E-4,5.754586309194565E-4,7.714693783782423E-4,9.593565482646227E-4,0.0011268946109339595,0.0012630249839276075,0.0013585883425548673,0.0014067762531340122,0.001403645146638155,0.0013482708018273115,0.0012429036432877183,0.0010927581461146474,9.058009600266814E-4,6.921945605427027E-4,4.637623205780983E-4,2.3319711908698082E-4,1.336030527454568E-5,-1.8359812384005636E-4,-3.46912449458614E-4,-4.679716657847166E-4,-5.407938733696938E-4,-5.624890909530222E-4,-5.334119196049869E-4,-4.572196921799332E-4,-3.406107716728002E-4,-1.9298773258924484E-4,-2.5823352189036086E-5,1.479914499213919E-4,3.1502480851486325E-4,4.620902764145285E-4,5.771702853962779E-4,6.501343450509012E-4,6.734839989803731E-4,6.428086780942976E-4,5.57172461412847E-4,4.19155927374959E-4,2.3481316748075187E-4,1.3244637557363603E-5,-2.3386844259221107E-4,-4.930642317049205E-4,-7.498731138184667E-4,-9.898195276036859E-4,-0.0011992902727797627,-0.001366502488963306,-0.0014822309603914618,-0.0015405109152197838,-0.0015390111366286874,-0.0014793031150475144,-0.001366745913401246,-0.0012102582259103656,-0.0010217201197519898,-8.152894442901015E-4,-6.064505432732403E-4,-4.110619775019586E-4,-2.4425852461718023E-4,-1.1948979954468086E-4,-4.754334804601967E-5,-3.5839391784975305E-5,-8.781907672528177E-5,-2.027036971412599E-4,-3.754065546672791E-4,-5.968526238575578E-4,-8.544449810869992E-4,-0.0011328886030241847,-0.0014150983188301325,-0.001683353097178042,-0.001920394948683679,-0.002110642846673727,-0.0022411919198930264,-0.0023027784191071987,-0.0022903995122760534,-0.0022037792950868607,-0.0020474193152040243,-0.0018304386176168919,-0.0015660012140870094,-0.0012705628760159016,-9.627902181819081E-4,-6.624060915783048E-4,-3.8884449168108404E-4,-1.59999675815925E-4,9.044497346621938E-6,1.070310827344656E-4,1.2739759404212236E-4,6.87647916493006E-5,-6.482833850895986E-5,-2.641297469381243E-4,-5.151444347575307E-4,-8.000194793567061E-4,-0.0010981149971485138,-0.0013873724965378642,-0.0016457131132483482,-0.001852559857070446,-0.0019901995547115803,-0.0020450667943805456,-0.002008696086704731,-0.0018784343264997005,-0.0016576983034610748,-0.0013559159124270082,-9.879799326881766E-4,-5.734111182391644E-4,-1.3511351426132023E-4,3.020453150384128E-4,7.128877914510667E-4,0.0010735623072832823,0.0013631944311782718,0.0015653080772608519,0.0016690443735569715,0.0016699671978130937,0.001570522552356124,0.0013799790758639574,0.0011139786802232265,7.93586194049567E-4,4.440172342583537E-4,9.30038295336999E-5,-2.309868432348594E-4,-5.006803548894823E-4,-6.918226717971265E-4,-7.84908072091639E-4,-7.665645098313689E-4,-6.306227878667414E-4,-3.7866129423491657E-4,-2.0110366676817648E-5,4.282290465198457E-4,9.431107901036739E-4,0.0014962774002924562,0.0020562049467116594,0.0025901610497385263,0.0030663306824862957,0.0034559883642941713,0.0037354526575654745,0.0038878023624420166,0.003904126351699233,0.003784316126257181,0.0035372392740100622,0.0031803613528609276,0.0027387409936636686,0.0022435372229665518,0.0017300298204645514,0.001235365867614746,7.960800430737436E-4,4.4564888230524957E-4,2.1214493608567864E-4,1.1624231410678476E-4,1.6962896916083992E-4,3.7402540328912437E-4,7.208026945590973E-4,0.0011913296766579151,0.0017579516861587763,0.0023856430780142546,0.0030341444071382284,0.0036605496425181627,0.004222087096422911,0.004679002333432436,0.0049972692504525185,0.005151023156940937,0.005124472547322512,0.004913222044706345,0.004524827003479004,0.0039786044508218765,0.003304614219814539,0.0025419348385185003,0.0017362559447064996,9.370048064738512E-4,1.941132650244981E-4,-4.4529649312607944E-4,-9.401598945260048E-4,-0.0012583628995344043,-0.0013791483361274004,-0.0012947912327945232,-0.0010114876786246896,-5.492977797985077E-4,5.8799090766115114E-5,7.68773490563035E-4,0.001528167980723083,0.0022793905809521675,0.0029634046368300915,0.0035236580297350883,0.00390991847962141,0.004081836901605129,0.004011917859315872,0.0036877573002129793,0.0031133051961660385,0.002309114206582308,0.0013114570174366236,1.7040646343957633E-4,-0.0010530924191698432,-0.0022909268736839294,-0.0034721465781331062,-0.004527578596025705,-0.0053945062682032585,-0.006021032575517893,-0.0063698976300656796,-0.006421418860554695,-0.006175396032631397,-0.0056517538614571095,-0.0048899115063250065,-0.003946809563785791,-0.0028937412425875664,-0.0018120997119694948,-7.883394137024879E-4,9.160373883787543E-5,7.480282220058143E-4,0.0011130099883303046,0.0011353446170687675,7.846074877306819E-4,5.3973650210537016E-5,-0.0010383679764345288,-0.0024494121316820383,-0.004113132134079933,-0.005943876691162586,-0.007841150276362896,-0.009695583954453468,-0.011395701207220554,-0.012835128232836723,-0.013919766061007977,-0.01457449421286583,-0.014748940244317055,-0.014421929605305195,-0.013604258187115192,-0.012339571490883827,-0.010703175328671932,-0.008798809722065926,-0.006753446534276009,-0.004710397683084011,-0.002821032190695405,-0.0012355901999399066,-9.357769886264578E-5,4.856671148445457E-4,4.116959753446281E-4,-3.6962778540328145E-4,-0.001870464184321463,-0.0040575359016656876,-0.00685113063082099,-0.01012676302343607,-0.013719477690756321,-0.01743069291114807,-0.021037248894572258,-0.024302296340465546,-0.02698742412030697,-0.02886546589434147,-0.029733220115303993,-0.029423482716083527,-0.027815626934170723,-0.024844160303473473,-0.02050473354756832,-0.014857197180390358,-0.008025452494621277,-1.9406128558330238E-4,0.008398334495723248,0.017468471080064774,0.026700401678681374,0.035759299993515015,0.044306524097919464,0.05201508477330208,0.05858483910560608,0.063756562769413,0.0673242062330246,0.06914467364549637,0.06914467364549637,0.0673242062330246,0.063756562769413,0.05858483910560608,0.05201508477330208,0.044306524097919464,0.035759299993515015,0.026700401678681374,0.017468471080064774,0.008398334495723248,-1.9406128558330238E-4,-0.008025452494621277,-0.014857197180390358,-0.02050473354756832,-0.024844160303473473,-0.027815626934170723,-0.029423482716083527,-0.029733220115303993,-0.02886546589434147,-0.02698742412030697,-0.024302296340465546,-0.021037248894572258,-0.01743069291114807,-0.013719477690756321,-0.01012676302343607,-0.00685113063082099,-0.0040575359016656876,-0.001870464184321463,-3.6962778540328145E-4,4.116959753446281E-4,4.856671148445457E-4,-9.357769886264578E-5,-0.0012355901999399066,-0.002821032190695405,-0.004710397683084011,-0.006753446534276009,-0.008798809722065926,-0.010703175328671932,-0.012339571490883827,-0.013604258187115192,-0.014421929605305195,-0.014748940244317055,-0.01457449421286583,-0.013919766061007977,-0.012835128232836723,-0.011395701207220554,-0.009695583954453468,-0.007841150276362896,-0.005943876691162586,-0.004113132134079933,-0.0024494121316820383,-0.0010383679764345288,5.3973650210537016E-5,7.846074877306819E-4,0.0011353446170687675,0.0011130099883303046,7.480282220058143E-4,9.160373883787543E-5,-7.883394137024879E-4,-0.0018120997119694948,-0.0028937412425875664,-0.003946809563785791,-0.0048899115063250065,-0.0056517538614571095,-0.006175396032631397,-0.006421418860554695,-0.0063698976300656796,-0.006021032575517893,-0.0053945062682032585,-0.004527578596025705,-0.0034721465781331062,-0.0022909268736839294,-0.0010530924191698432,1.7040646343957633E-4,0.0013114570174366236,0.002309114206582308,0.0031133051961660385,0.0036877573002129793,0.004011917859315872,0.004081836901605129,0.00390991847962141,0.0035236580297350883,0.0029634046368300915,0.0022793905809521675,0.001528167980723083,7.68773490563035E-4,5.8799090766115114E-5,-5.492977797985077E-4,-0.0010114876786246896,-0.0012947912327945232,-0.0013791483361274004,-0.0012583628995344043,-9.401598945260048E-4,-4.4529649312607944E-4,1.941132650244981E-4,9.370048064738512E-4,0.0017362559447064996,0.0025419348385185003,0.003304614219814539,0.0039786044508218765,0.004524827003479004,0.004913222044706345,0.005124472547322512,0.005151023156940937,0.0049972692504525185,0.004679002333432436,0.004222087096422911,0.0036605496425181627,0.0030341444071382284,0.0023856430780142546,0.0017579516861587763,0.0011913296766579151,7.208026945590973E-4,3.7402540328912437E-4,1.6962896916083992E-4,1.1624231410678476E-4,2.1214493608567864E-4,4.4564888230524957E-4,7.960800430737436E-4,0.001235365867614746,0.0017300298204645514,0.0022435372229665518,0.0027387409936636686,0.0031803613528609276,0.0035372392740100622,0.003784316126257181,0.003904126351699233,0.0038878023624420166,0.0037354526575654745,0.0034559883642941713,0.0030663306824862957,0.0025901610497385263,0.0020562049467116594,0.0014962774002924562,9.431107901036739E-4,4.282290465198457E-4,-2.0110366676817648E-5,-3.7866129423491657E-4,-6.306227878667414E-4,-7.665645098313689E-4,-7.84908072091639E-4,-6.918226717971265E-4,-5.006803548894823E-4,-2.309868432348594E-4,9.30038295336999E-5,4.440172342583537E-4,7.93586194049567E-4,0.0011139786802232265,0.0013799790758639574,0.001570522552356124,0.0016699671978130937,0.0016690443735569715,0.0015653080772608519,0.0013631944311782718,0.0010735623072832823,7.128877914510667E-4,3.020453150384128E-4,-1.3511351426132023E-4,-5.734111182391644E-4,-9.879799326881766E-4,-0.0013559159124270082,-0.0016576983034610748,-0.0018784343264997005,-0.002008696086704731,-0.0020450667943805456,-0.0019901995547115803,-0.001852559857070446,-0.0016457131132483482,-0.0013873724965378642,-0.0010981149971485138,-8.000194793567061E-4,-5.151444347575307E-4,-2.641297469381243E-4,-6.482833850895986E-5,6.87647916493006E-5,1.2739759404212236E-4,1.070310827344656E-4,9.044497346621938E-6,-1.59999675815925E-4,-3.8884449168108404E-4,-6.624060915783048E-4,-9.627902181819081E-4,-0.0012705628760159016,-0.0015660012140870094,-0.0018304386176168919,-0.0020474193152040243,-0.0022037792950868607,-0.0022903995122760534,-0.0023027784191071987,-0.0022411919198930264,-0.002110642846673727,-0.001920394948683679,-0.001683353097178042,-0.0014150983188301325,-0.0011328886030241847,-8.544449810869992E-4,-5.968526238575578E-4,-3.754065546672791E-4,-2.027036971412599E-4,-8.781907672528177E-5,-3.5839391784975305E-5,-4.754334804601967E-5,-1.1948979954468086E-4,-2.4425852461718023E-4,-4.110619775019586E-4,-6.064505432732403E-4,-8.152894442901015E-4,-0.0010217201197519898,-0.0012102582259103656,-0.001366745913401246,-0.0014793031150475144,-0.0015390111366286874,-0.0015405109152197838,-0.0014822309603914618,-0.001366502488963306,-0.0011992902727797627,-9.898195276036859E-4,-7.498731138184667E-4,-4.930642317049205E-4,-2.3386844259221107E-4,1.3244637557363603E-5,2.3481316748075187E-4,4.19155927374959E-4,5.57172461412847E-4,6.428086780942976E-4,6.734839989803731E-4,6.501343450509012E-4,5.771702853962779E-4,4.620902764145285E-4,3.1502480851486325E-4,1.479914499213919E-4,-2.5823352189036086E-5,-1.9298773258924484E-4,-3.406107716728002E-4,-4.572196921799332E-4,-5.334119196049869E-4,-5.624890909530222E-4,-5.407938733696938E-4,-4.679716657847166E-4,-3.46912449458614E-4,-1.8359812384005636E-4,1.336030527454568E-5,2.3319711908698082E-4,4.637623205780983E-4,6.921945605427027E-4,9.058009600266814E-4,0.0010927581461146474,0.0012429036432877183,0.0013482708018273115,0.001403645146638155,0.0014067762531340122,0.0013585883425548673,0.0012630249839276075,0.0011268946109339595,9.593565482646227E-4,7.714693783782423E-4,5.754586309194565E-4,3.840607241727412E-4,2.0973681239411235E-4,6.400272104656324E-5,-4.327772694523446E-5,-1.0438119352329522E-4,-1.1422827810747549E-4,-7.058848859742284E-5,2.575004327809438E-5,1.710843644104898E-4,3.5895180189982057E-4,5.805459804832935E-4,8.251464460045099E-4,0.0010807289509102702,0.001334545435383916,0.001573855523020029,0.0017864631954580545,0.0019614456687122583,0.002089534653350711,0.002163664437830448,0.0021791793406009674,0.0021340770181268454,0.0020289572421461344,0.0018670330755412579,0.0016538002528250217,0.0013968131970614195,0.0011051764013245702,7.891962886787951E-4,4.5975486864335835E-4,1.2790676555596292E-4,-1.9567001436371356E-4,-5.011202883906662E-4,-7.797284051775932E-4,-0.0010243176948279142,-0.0012294170446693897,-0.0013913477305322886,-0.001508324989117682,-0.0015803587157279253,-0.0016091193538159132,-0.0015977213624864817,-0.0015505029587075114,-0.0014727171510457993,-0.0013702119467779994,-0.0012491375673562288,-0.0011156742693856359,-9.75638278760016E-4,-8.346185786649585E-4,-6.971539696678519E-4,-5.673483829014003E-4,-4.4828696991316974E-4,-3.421740548219532E-4,-2.5030970573425293E-4,-1.732944801915437E-4,-1.1093106149928644E-4,-6.246339762583375E-5,-2.6618803531164303E-5,-1.884515654637653E-6,1.348849582427647E-5,2.1263915186864324E-5,2.3224682081490755E-5,6.581512570846826E-5" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="frac" />
// Retrieval info: 	<generic name="coeffBitWidth" value="32" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="31" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="frac" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="31" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_2_10hz_nco.vo
// RELATED_FILES: fir_2_10hz_nco.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_2_10hz_nco_0002_rtl_core.vhd, fir_2_10hz_nco_0002_ast.vhd, fir_2_10hz_nco_0002.vhd
