-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VkEf2gTPUvDE9AsvqNRzyQL5kuAcGHy6OoKXMOFYbFV/LHmU99Mpw2TTbOhpOmyCgYxPLCLpXUFE
wHooPDxFc/ANDQNmsYDKOgdwAFVyhx7tBwMk+C92GBc2ged05WUu9q+yKCk4FOJYF9+5kLBIN5TO
vXjhRxULStYWOoGlKZKElcelH+3oyzPcRomIlRYOOwgo1zphRQ1nvdEOSkEYQPwveEeiwtbctb9s
U3CCKf97YWSXJlT5dxfoDSPamDXc0j0mw/xnUTRVoHrjrxfsJtRY27oyavBUl64eklgUIBleSvSi
ncqnZQAXwOyJp6XysRzp5Te5V+SCX6GbZ4JMEA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
YZsQ+aaG0qix80sak1H6kixg23OQw/47gRkG5P7dS8NiMo4dQjIV+T+6NLOOVs2TXbAcHWGxiomb
rCYONM/6c1bZX6ZgDkshPrD8AqonCdHo5mDrWRh/rVc3IYB+X2TbGaLeWuCWQYrrnzsqE0xIV5cS
Uyg+rAD8/88kKJhK+B1jyKQkCY8JzouFRre/9mgE2L2KWnccm48QhXvWA3AeAd6VV7OPReVVIsIr
YWRQ3By5ySzwA+fC3E/kad5g5qTtF6T4nVuBIpgS0642tKQxyBUomEsviIv93tZco1hZwYaEnv2e
iunHwS31j1dT6pWMJNyh5jYuehaWv+ntiS01txscLeQOVA6z0QluG4rgr8/Gnbga9n7MpeWIZtdt
HFTUQnFp+tgOIVpFEvEUeYhQnYQRO1hunlRPEmd8w1xxj8Z+3YiJZ+QdL8gFSsmY1+IA/PSP/r9O
3Uo1efciu/agAml7t1VDerBFfr46ruWKIfxgQakyF9IpHqPHhqPN3NdUDgxc4cmxeMrKIGWo7qKM
2cSwPc24Ht8AeP/PL/tGcGrN9drd0N/RoYQCNGmRzZLvkCuSqyrCSePs1LbsruneVPjR4+SGeo6l
f///HEFtApdWJqsNCL38Ov1HSVv0pPhCPyy+QsJ2NvCnx3KRJTBWvAEgXxRKVALgHv8wUijok+0z
t+TMb1K59neSMGVdZwu5uP+w734WnV39dVA3D1QKTPVRvuil29+gfEjpeA7qG5fPAETJX9gch34d
V+HGoBS3ALm1XG17b53EQp98miG0drKGWniaWGvuyRK7oW3wCD5IyXM9mVuYnn97eHsSV7H0Eljc
Q1NPFdIw5IIcehaGfoit4Yu9uGr1PEef1RMoxbsKTndxv85zUcULnNabsmfvvWExlPhz3BUtcZte
oSdB8VpnxQHa3k0L6C/o6Jkoxde/k7GIeTFFkd2XlBL6X52b6X7T21D/e5XlObuT8IUsLhZtdOvT
mEivuxzmKlxV+PTrS0rBIBkfD3IKe9nlztgkJCmu9FDFOThJd+Kqge9V9GFTUmX3fKeO6miQVcb4
bpAT0bCKUIXtElMurf2jDbtCZVSaL3fLh63n12nmjhwAtD7l18/7ownEM+Anwtx5ArMq8fF9XmX6
PrO1cqnIzAjGQkcUvjBAKjcPdnRQ0058+9wEIfZD6nwv8KyFyUl+ZPzVqEmA66eiQ/aWXC9Kljgb
oyE5CkIoyPXwYo4eHScDkvHo4gEGOgT/PvA1OWk87fHw5tTmPmIgQMK6BeLkO2VLDNq4svUKVxXC
ML453wodOAEwTkz2wxqHrVhE6rLp8dSZ6RWO2ccym/lwt6hIedHO9HNT485+qH8ync0CKhqrVoC/
rvRARqRJhIl1T8oZ11oxMFv48V5Cd5rX4NeJOsJrRZVF1HJgVDCtTPaL+D0FSpP/RUUlLraIIk/2
Hy7MQ3ciZg3Fi27Mu6CUn8nb+B1V22FAND8x2s4j5Xy+Y2QrJ//HTSxl3vM/Gfn4qQFxB3w0obv6
JOge3qcN4sHMYhxyrh87Fza342qmMYLfWYUzCmjkNR40CdhoN7P92Vpbw5XisID+3OISeDLz7uCP
Tcn/CWivo8oKOLc1h+gADalLZP+U064vUYGIgYchmUK8f72HT5+hMfCGDw0Mp9tA8PtThTE6uzrn
GAEePXHe5KYhqfYO9THebTZcldG9ofmX49hm99Cu1W1hteW1ujMLfUBUgH4n3e2KhtZOOIapAhFu
jTjcCeMIoAylUeXLg5bkyBzLwD7zrK7VyFscDXcEp2RqhhCXyVy1vkvQW+WHbeIecE1AbKHBjV/1
8K3/Ze2RhglPaE2rIdIT8jpAA7qgSBXzA2l0VLPerKIfqF8uEldM/LrABwbzjUQ0zn7nuEVuZDdg
1bM1+v8knpOjiKIp4t/6imis0qxSs88ZG0nX6hXh8pYb8hLhcH7afCL8Lb/eZkS99QqndeKVT8Ug
CkRmMjDCymdM+ILRdMM+fV5y0MvlvcTbw+IHXEa+LRzBtebxYYH0pyTTpoHX63IrpBZCKGQtiQCY
7QmfS2QC6FwGj3IHcfbbpzDIGOCtTdE+BYdbLqtiXcQvm6/wZTAtO/PNZPoWMADZbAE1XrbyAtwS
2wJrD31Hl6pT1Cczk+LNIMiuq3J5g/npa3YkhpUP1XD2slbl8yOoDGSAkB79VU/XFRUZvcllNIOr
rb4V3DjRF65npWUHVNoxCk8OwUX3wUDx2awsphO40YCkC8RK4HLIymg4C903dLJDko+O6HUimfun
ybnxndLLig5QKNM3V2aAFgKR5becGbKIeGGjT6rWvG4wlnJxEmDEs8MwLUycuHXfdbd7P0N0W1QA
GYPGxgYROu20B2kH0F/TAiwshIxyz7RGBkcc1x3eLLyE6jH8tieR+AEKqt2cwhHAoh41cMpIMYgv
K4cWNtzH/wJUYFVDcqFiIeX12W9rJPZb2rJev10eCig3inOI+PBWC9XZjwT732GMEhgyE3zseu/y
NaMMzJXDNQH0s7sd10fqig4w+XQ8RP1gApKbyJ3T/gtucR5xH8knjS1h/E28YsIzhROveaYb2QsG
FgMllx8or9yrR2TlaclMjq43ANWmg02TlwFPj5ohB6EOuXjwqWrM+BoJW0kuaUTL6rahfUX1qJXl
zJqeI8rDoHT7fi90m8QJhp+tGXqO0Bdm4rkrHCVvI0AYmuL1LjuEv/ABhoh1ABF1TE52Os9uFY7g
QU0N02E1ZkXCFBO8pPINy7VRpd90jM7noOxnOJXPA5FAAfpJ5Ym9EY9CRNTFDvdjg+xXqYzOfark
7DNzy/grLS/2nC92x4Y4ADmX/Is58q3KA/i8meTPAabTzU60x5GMY/N4xq/3MXA0gaTeL8nYYbqW
LOcn1mFJZ0k21QRb6NjG1KXmXD94ZseZh9fJcGRnHoc0p9KdH3r2YbMEz4QMYHMCmmtUWTomWmWw
D7pGELHdKMmgV6mcMgIueDnqZ8ZZrdxpGZSKPNrqt/DVDJvx6dZYDqm5lV6xmmXqtffVxJ4wTL7y
tY3gdeSdkFfKVLnwMubUUtL1QM9i50pKx1gIRPfiYAKxtatv5QNv5NYydlqIGpD1urdtxgMfobC6
vmTBPImwMqsdQUJa9pnPS8l5d2Noj3m+P+uCXuiaoJNdIrF0mF2WhwQLzdRmjixi06lqsADRIsBZ
S1x/u4Pl+5CffXOVyjrU/68hTfH7nJnz/CvpqJigFIx9LgrEj9K5rgiQopmH3FSfCB+8kultAkE/
X+0x9OBucD3qkFTIWpSSnuAjgxXdMr5LdgPzuFdHPBmO+RuH0zuJ/FMHrM0o1qvYO7+ngwcUbgw1
o/tHcw49K8kOwMQhJYNPOIIbko6Xo+tOssIcVym7UWHV0f8BFRAtbsAcWpgiUYmgzVXmdBjIdaUC
2Lu1I+jQQ4vvbU+BHDChJiJ9lMfitMijwp2kOmCNRhVbWpdpf6NX/w5CJrFB+S7i58U+5FCp78hS
ngdeLZ2Tg/W2D73eMmKCoAUkYfifE/fKgBdFnqPsphrhPGSs79QTEZT6hrF36bP0M8/2sHzL1/nx
XtwO4wNJNiFcREaKLAm/0bsIAgJtLsOqIbSrPotC/8Xbcbdb3HB2l5kW/UF2ItZsWLIP9W+bBx8z
m7qMq+3fXFX9Fel8eAME9EWqVGtHzC2PjZvXizGTGx9et0D8LlD7nlwJ+VBGvQ5NAHg/g1m9m/lF
12GZbd7uV0LAfzS9YtrxxnhF5s6Yt0HTipEq/VH2hAtn7bLQk/5hpsDDsdcijl+53vkLQ/LYz/Z5
tJPD6gyf+t8kExRquWUj7SkFeWc8mhB11si6fWr5S0pk+YtxWxyKc10QlYlHW72ckR9ue/jGai1v
8+M7rFUjG6GCO4J+HGnfrER7IAiDcFePtXjOjdYwsZSRMiKDJ/+C6zCZ2qTBXZt2Pks4ez/xas4J
UeaZV9fcLZ23RZZwuJa0yyQMl3dBHxnifFqI4BSoaMNT57gqTWkujwSa7dX4yLBuD2iWCvC8bnVf
+dbfJWjWQ0EmbFupVCFlMYdQX/i+G1lqknqtAhU84nG7Lp6tO/Oz6MOzp+l6rFcCs2nhAc8Diwno
Xccobf0D2RnXB2Qkn0Z+z9CBaCozsRYHoQpHeXF3WUZ4dGnjC5v0CshVINCBWZZKDkPDqJtW4w6p
8UYs9qLMbUUASSp7P/5a6IDLNrV3/gFRuUGOP4L/I2HGp1vUA+UEPvNCefRx/4RCm+n0QeJq3Zzd
rmonD3Muxjd8gImTVI5WAuN9HYwbqXIDGWuTAABYNNr6yp/CMGtlGQc1A41UUJyJApHml8yX8LV1
gfkG3UVfo/IuesaWQaKEsdhvzV+zEMp3N4ieqYRIQh941Wee+gc61zExltOb7dRUgy5y29a9hfvA
TT1nychyae/VDWNb0xsAPryH5RyUWzpV35CRQwAorT6bYWNDN12qPpJIz3w5pjX0W0WL0WtUVp7C
LK6qkZw7XMflLluDNtJEWSYO+GmZ3cZntPeUlMnUpzMkOTVJ2yqnyMEu4M9db2/pjcTjSBHjTDd1
Foy93l4amgaZzd4kB8vqmATfMfZ10Etyp1e6vmiqIvs7apaftjV0HM8mbhUWV9M1PUMIqXvxCgba
+uC9NpMWef9+Fya5cijgyNE8ElO4KO+JoV73MxULQRPkSlcMl9C5YwCJiu2o29rZj88c+NmTbtoh
QEawh6YSZ1dL1+SDGq5v4VWZrF8sGGHHVPUk7ytroL8cyG51A2BJXPHECXCdlDZPR7tBksJheisv
FpgCO49a63/zfmmE+ft/XdpaP6n7NVv6qtt/5OTxV5vcNVBEPqjVtTcSqESIxEITKrTt5+nblVk9
fRReQ8YgzZftZRZeT7/y3jG4Cmec2Z7SReW3l1jmpjeIdKGSlsGtsm7D0qLJKsm9liQ/yfPurPLG
q98cFKnooxyS1OhMJrnAWzDIYugIfq4JdhCTPKUZ4lQnpldkMmcH1sgh5jW3Od2kiqsu1+o8+ZhN
dAJwKxv3mO03dWCw/E+YOAe5OBYwwwb0fzztti9cesY/ItMEJGvNiqdtEnWshJlKNc63h1fXeEoR
C64b5Ym3Vwb0VQYnFERLxEhDv3YG9DR3VPXOzbljlKZGTqqsXMS41l36zTVagNSI6VpQfUI8Exnb
1vuWIik86AxLgylRyMRr13Sp2rcebB0zGxjtSOZZFkPl8tSbK1TIIAfyODNy8bZoxqbCLxwMZlba
uEBgL56oQF5Ve/PETcBxwSy0rOfufR4we9KbdFJRkoUHIXUTNc+UdEvE2gR9N52IoKf6qtO4IS29
TA0+reQOTyIwIdMS6/LFacHTCyvOv13TDzaNivngarbNnlIaPaAflZb5ygA+Gxtr0q2HvYTqJo7y
x+Umu0dxI12cuVFTl3UuRpJaPU5kYUW86d3AjRMY93MjGAME8brKz+IWi0erVebuhX2ZGg36sZU2
InpGOR4Y3Txhxls612bCEQ6vlTi8l64arYjn2AD0fTKxnfhuGbpanukmyG+SHBpaln4t9Ayp7fCk
/o/Ewc+MpPEg66Cffbhb0LR9Bld11oTMCKG3FkOUnr9y/qYmm9DruKTujmYlNQoU0uN7mKZLYnZ4
zit256XI6GIW9ZFkYdsnMkfSRgOvE1G9fHsGD5oljuR31Sjs7Sla5YVoUwqvfSdytoqc7fn+gJYb
Yr4fsSRhGDy+m8TnQMl2od+B40Kv+0Ep5YsxFAAmy/lvIzhwqgiwfJDrvu8oM40BDqAroFdQ8Mlu
mq4HYIu7L+2r9c1P2kyLDRrW1FW16AwlZ8IkKLyJPkacl/LiuUNGx1yAoHLdfoMWhuJoKeMapGZP
LZr6ZGF7BmfgPVM6Pkc98tD8TaFzj4DwP1gzjiH/kcIdXybg9P3P+tV4YfOIAVB2Y8kYPo0RWZe9
3ZJgweaU27WzSRTUOhV1gNV8VwdG7iBMdfM3u8h6OH3n06tqGS2JipAjMkoUEFoCZ34G/yEJ4Dvz
lSApXAEYeLGNPc4F2+wvUAtOpabIWumK34ZousVcu2gFwQLEfz3nsbHsihhTTrCAKPYEP4Mcje6w
KsGEf5o+k2fy8oLkOp8rkvcMLAJNrBW+G+iHT+a2VBdP1EjO7ED4n2y5EmAzf9/KhD1AP8bXFMjE
M3R7mFBm+Cxm56MDwGJUoBa/rzGYBpbPrYm/AdU14dDytjxU8AMlyLp2OMOuld/W+lJPTfoSBVMe
evqZi08eun72vxAIGat8MYVllettpZBgtPstrSLHk8+yggOQC+k1vzpA1fog9C1PZ4dNDDq1K/41
el7n5pfPl63xRZjpb4P4v8ZC8nILiag3zUQ13duSrhAyrkI0pWNuQ5ZqCfQ5ugHX1ur3C+fGsZUU
NycCva3HBnEy2rzVrMHwhXd69n4MCb4pUXst4J4Aq5tYwmJroOnzk9FELPC8iPrtWjj5gGTP0f1x
dzf3hihZOiVa65TxcjrBnohg7UuCbbmOPmcClpAi9tmALPRpcl34TseJqf0fqGSxq/zjYw41VXZq
a/u8do/SgrDSPjiKidbN95PiMHcP4PgkVl0GqOFk3B7paPfIjWMBoFp15DFEcVI4dQEhtra0RFWl
myhrTgVgt+joGRdeubbADKaH3MhZlBTspdT5eRLskdJQkbQTbe5Kn41qmYeccg8qBZyY8jLZ6YWs
4WYePOj24ptsBGwEyB8UsBwvI1bQhZBMXlEeaO1HZrX+wvoDobjeoDd5MjbU2utFOClI/NATtEEI
7aecxQvmGIVK5zRnUgUAjqo70W/ZZUoiejMiPcfzNy0UknRW8BHhhalZtnubvdWptzinEomrgSAW
O+XpcHvPChlxKlP1c+YfqI3kOG5t5/tkcTbWLEJlY8SPky8IcOUvoruXbQ6d0tDTolOOsPCUHjH7
X2tgYv6uzV5G8Uwpx1W9TKelLB3zOkIuQbUh/XITIvj8Qidv91nnNuK52jFPLqR1HxKJJ50xu2ve
F6T/MGdRG1nBPLnwqCEm/mM1dHAAxagZeALlh61grLPi0Z+QlT6RKgtEQIqawWgYEzUvxgWYupxw
CaTbOeV3bJFtH8pX4PDisBCZ5+AasBPt1pY3omSJ2YiZpC6rtkoQlIZIpKpo9ux+XTFP15zvuJ8D
bV6ZA6XsNcaLwl/DkdUZo6CQQvK+kz/FcDOZqsP63+qSVkcl9fYeNTCWiYImKBjwkGuiuGGVU/X2
Ggsoofk5g35nj6MXrVPS9CiGm/8+IkHMgpxSJEcqku6WzZBYt2/PM6QdTJ2bSu/xyxrGnjUH1LrN
lp3EQlwSxglDIf+6edm23G3jJKjZgde5DjPjDTArQk7u+7Oj67VUXAi1RepmOnRTWbfENGtmMD1X
hquchlhqlO8EMPRke7yr4F2riO+ecEFlP3mnXM23v62bBUYc3aV0MRK6Wmi1In5U/3Be9O+mVuLn
DfCzQUCqi49vv8ntKjntJO6aYb88vdcvFCMzBgewKnHEqeCg4WOTxNkhu8eZYJrHYO5ceFTcB8VZ
vFrxSdG+tJ0lL9IVTaDkdx2v2oRhMS5ivTxXBnSGQ+E3xrHhdVK1JmJnO9ZzR6BpLvExOfgfWFZT
UUp0xyuifYiWEsDlpouQO3pdp3I1Gb4dFFZuAvEOsxyqRHyNS9qSxmNHpRNmRJzCsPa62eSF/77R
ISlWq8IUW0vvDW38d2WL2/YPUAy77e5o/OP1geZnHDJAatKVjzj3dXpzkAZvnqkkn+9sHDGDwdRT
iOfJfAS8CvCNA4xowRI7EC0l+zgDwPB9UgHczsSKBJymChL4l4y218wWeB16Q8OBcmpaNz5fHZub
6w3eZ7TFDUW9SYaaE8mS8C56/5KYBIaVqEzsAsRIGeSWC+JtAZyRcB0OEkVhm3ROcYOooiTqoSxg
Cq4awB8kfoljveNa4NjyJ6HEkWK+GDNCzRfxUZz+cnG3Vru9kfxefRw8aYn6q+ChUvl25/CHw+jg
6f+zZM/JGumjfHMQ4iw2sMKxD41ZMXGRjhGBUxwOlGU4xEepOa8VGfbszQAforNruWiGF5XFihMR
lN0Gw96Z09Iti+3vaDNu6vEF9saAiqJIXsBgS/bZG4chQ1fkny9jpPo8wsAaCJIeRhQXKUodoMuk
AwI4jjGCWmFsTtIjRR/McWJKBlDYIFe9/7zSLHSpRNy5OTQh2Q4wrpDW8xNxQXkDGHGqLg8Dn/8v
OI3JAJe7/Qc4K+BFO4kNLTcMyFN9MsKRQ3lZ4A0Ica69FtsQ29OGM0I3yp3S8aGv7KKSo98kHUF6
AyKV+cNABEBez1UoACmiZ5OBrNogiv0Io5QcTtDb6WCHWxZRgbJYsHdSU6qeIQ8YdMNiD11hbBiP
2hZB3PDU8E09ZlxvW7o0kayjkOhutfgD+sYFN44BOEkv9BRI289JW+hCdHYlW3wLOoBJxpCJ4q6U
I6B0FcueGzcjwDN8GkXxvdAcloHy79zmzrKli8JrTko9TqDndgaPX0ZSHgLYOFe1W0ImBD95dFOx
guF3+Xv2yJY/F6jl7nMLDcwCLJjMpOZc9xX7l5zbGKXZG3gjV88r8Pyq74kAM7hV8w7gnwJ+IlCt
0FqgBfksD8f0jkd85rELTIkpkOnpgb+nSm1VHwfZqK7FrPNorTJBEW3gMqKmVCePVih9yxJBe4O5
QU5QA84P2msLMf9TPr69ZGmZyqZrdTBfcuHE5bCzuSPxRjOFUcEhmVmGmh5LUiKpNw6AF+uyxpkE
suI2aJP7zsIlFXb71Ms3CxlxWeos4T8wQ0SmNQ98VAn7GbCg7J2NvkLHFMTznV4ejMNAfLpURz6O
R47Wvwg5yGsGFqtUQKtgnng3eM6434tVBNRRNlly6TbhKQZSc+lw1lR5leYoYve8cOcBpccjhT+B
lXL+TVTUuKMAA9wBSfLk58+7kBlAD/rWKO7qjy3BXPCbjiOaCy/NyXynA/a+ML52gfuEtYcOtJ+z
EZqYgcpHZH0cmw833zDUA7sZyFj79k4ERMrmgmjUJE7LGGG9X1LQ+Suh5iRBCQWa/HTeq8wqmviZ
yk0W1aPO4BjHjVSVMOq1gXR9GajMnKATYQeXxmHWJHOyruFGftTANTXOEB8x9y2eTedj7Mxzl2TD
q9NztKJjssL+cuOtYFng34hr/653oRGkdduapBzIVB07mfDa1YyldE3hZ/OVrn2b7PdFlzSI48qn
U5lUrQnFbbXyljpbzyOy9i9Gka/V1a8iLRrc+e8BGuSSUGrIXXMQB6PLzaiZPK5Dg4RhptqRFLpo
nRYewcePaEawFsV6EibyRgJ6VO0qTZ0z8X8Mkp1QrvfIGoCInZzHMtUIpHPYUqxZ8i6Slc48z0Ek
Jh0TqhYc9XmzIF1QZ4gnce1fXCP/aCElnePYL6zBsLugLbY+CArkKQ1YAY8seqb7MOOyWfbYydIl
a5zFOKS46tNt/efUOdTO+1eMeLgs3GTCT0skgN7/tr+Bf1C2KqwEaBif0EGRn1IDEjpY7XgbVfEn
fdg4ZNFRv12Y4zPlfWIOSZow1BqJa0wz0im/OjzxJRWTGAPsOLCx7fh7YtHGPt5QDDXXiC5P+V2K
oFVQq+aML5y2GxoYtJo4HlRWIWalCngknwslh8fzjoEJf1vAzwuYD4+szG+y+w4VsD5PGrLSoaSb
HfOJjT6ijamxUPFbse53BFprAU+GUVGKD7OvN2ZgKwrRk9FPqQYpAxNDXL+FyTnifVpZzw3tUtVa
njlCe2uHT/58Yi60g799d9drmOt04VW7RNY1yHopjXwR3zFQ71kfds4QVPGi5D4rMXXUcYfQvkDl
zggbnQk73Em4UlapGbNqBQiRoeK8bazf2OfJYHJf7IUU4Q1c+446GGLmbAi+XzztTUww7renG36x
o89CRbIQbmS8N6ByzlioGsB+nL05iqybzjXwcDYrndnlhDkUTBS0Y02ovCDXiVycm0YPP4LVv3pH
fQpeg1YxZXP55wA7BN0YeXUERdxyeIM07LIjnVGFOtO20/7wyBi9LhzUK7m4y8eyUWlLxQNRbAez
KmhMkZ88oH98yP9ohayqFCbbqEJEq4po8S2K1IU8HXGmRFwQ/Mq06eWhmt/QfSgck0Nb8RnL4Uai
S1qw5u8Njv8tGckpbWm0BZG1DvnNS9WpD2NwV0hYxeNVzR3igg+mFt/RnYbK6wAx+ror5AYYMamC
tIZsVNTe7HVjKUuflgf6k+9SyS75Dft3zXAoXOXyEu9Z1qXesimMxBUh2B5WbxokiAj/AuOotAsI
qxmrMX/KAtthw2cKjX5whZah43ktu0AaCI3gC9HP7kGi0RJX31z+8N0m2LVTaycTGWNCq1cJqHGD
KRyeuF+zZbMY16VtYkeH3l/Nur82LfDLJCYqND3tBiQi3Icl0ZwiNHUEUA2MvXaPnuQzIyD9+wNZ
HEOoPTG6d2/HTkbId6/BORGgzorzojS9kUgviv2cPAvbqFlFIdQTjWT4Dpzjg4Gt8uQXBcPiOxL3
yteAn02qhzCRsoODLFE7qxJN+OTz0hyYH8n8xi/dNDJqbs1gMdMYZU9+fQituaQ/DhNy11VObYbV
lkcwZSUcgCTgaroXiPq0ssU3YH8b+l/jIqft4Ww8Rs+P7KE/5NIPpDYHhcWCveLnr1YI+axKA13w
X1D/m2I8e5YQ1K7Bp0CIDkBhqn9VfPf9TFDm2fGajIY+THvgsB77vAdOFgAXnLCEIxa2s4Af71c4
5Kk3PWY4kSpoCi96DGEVmLNNJJWfTIb6Lv4CdeLoeEHZvGhGPcoQ/V4CflnNToXRlQe19qBlS2iy
2FsVUAxOVCgQTARf6OF8AHVS8Z6DujpleNRumAf4WSTO6BLoaBKuDF6zqCTaMPBAuR/zv4uVkKtg
M0iapUaJk2tVKXlwp1Nc8tTST57b7mwO56GhFAQR4eS2qEcmygSFIc51+9BgomN/rkRgp5e/Rjnw
RmFnEKUXBLzYppp7nnM8Fo7qmOAaYIEsqAPyPcag/VdWYWyKgwBJtNfwALf64Vves8SacI0+3iUk
SPAAaCfv9G3FDhTuGaZk0LH1iOz5COgOV+Cd86wdvoJOICBcwW86HYkygbinfGBbWv220LCpikp9
19jNNnsFDwX//DJfxilijsRpfMocxieTUvlLgbXGblNCclOOaJwjG9tMjFOpHaMEfSHUGlJQchSR
8CtxObRCk7s6FGvJbMJzdXdOwX3RnEsHO4pGMDUmAMQhipp29FaLPc64MayHmzGUIxZ0eF62hu4T
q4c9myes6+U0qB3unA21QuVtsqS6pWfS04B8Z8MbJSTj0mBsziH9lODf6aazwb1wLAck+hRokv18
tgkQHcbVRwY/qw0cPh4v1vZ7ZpTlupYBTJ/tiPXNzveHRqNL4JIoGZtxtm1xJ+yUQ7FCbqTw5CI1
VkakVt0Jx0a/meivq81Bk8sYJb3viqnimA1lSfwHAhclT1ZtkmYrqJ4qZ4PDcleGTgazvx2INVQG
rIXPG9/nkjo+oLL69wHooOpi3qpdFDVWRS6xGRtjOIpbC/QMM5lm5FUtt4+VXWWH5lSoWFG9eI55
jWQSq1zzD8/FK9/JR2AA/kOZfzaC3Yc9NVuMekP66iUAX2wlncu4Ulrv485dxX0nEHsfIB2FUqYe
K8NjS9ozJLyiSjANGYZnF0rpAOu8DFaBGYf2msrMa0h+j4jdsyzqYIwYRykvz1h/7HpTjeQlf51Y
TqHKzoPxesajrLY7SfZ7u2xdCBMsHhevOYrN9AYV1Rr8MNpzKIHFs5gOOCN1qAV7gZ3N1k/3CndK
x1x/Uw41e1BdEn7peVFZ9IUn6OfpfNUCR1PwHkltMFFLiZZ9LjM7TWBt8Fbgc2SOL5QRFFzKITLT
dj2joKeFg7l8CRtuFfvveNUZfmg+FmUXlOPlP+VUINF1zUgJYr+a8devLeFqI7FznNY4FQFEdr/0
FD1WPgM5993M1tYHgSaCpx2U2vgfIQ6V5QEGkQFHE3JrOazNoY6LkdkEebnZ89tzsJj25/v8Hn0E
HTOdANRztw+KFGNca3L+V+Qoy3hrns0MUxWbn60qoZ5WUZ+/Ixwnk2nnB3S/aVA4CVL1p88TwxXV
3XyzwrCezyV/epG+b49+qy5XfVY8qOZLDgDH/uWRWNMN5QBf1esmaV3y1vMg14CX3Y31sqWJVQek
WtAjDzCIxR28pJCNUD/P4AMS0sh/OEh4fPPnuS1Ise2VhRGPy/u9LiyGhnlst7BlZvztf9x0hloR
PFAYOTBhUsNZHoLFtuePgt0DuuuXGLliRUpznRNAa84cIbnd8+QAMLUtWfwyOijKMcVpNvvfXhIO
zXlxyvmNioWl/KBJxAM+aVflqPXWn7cs5coO/sXRHVwMrYC+CY9nXST3Vu0VZjngLb1aZO/hMNNR
SVkKZOrZ9kFnFURRKgXD5oWIvNzJIpZUfRupABBGzSZCsmg50Lpy//c/dem8h/NA6eSS37eCGD0l
twFL8TdOb+M4fbTQRmLJoLAQIQoDHDOyd6mrsjrfundkrQe5U3+3K7AF0aZNRrhB41zUfTQQDEYx
UQc9tzLGDt3qaKmIw7vKZ5ssXmL8E8o8PuVnsykR23C+xO3ckbRcyZU4+V6ZDN1gYOIG/TOr0R+O
ULWbO9YJutakG1ZZBt3Z9AFIlxZXMV9KRQtpfzVWYBig898On/5KhikzMv4pXP/nrzVedSTN/7O1
kNwXMJ+sd/IvQd+rA8bnIWf/pek13w9pQ9OewVzax5LvNMk3KAMcyONvrCrQVmjPY+ds6C9zlboz
CucIfr/IKrZ0O6z5YuX71wR6H4F8Q7zNlNwve+PneTQ+7LrIBkgX2ZlI/6+67TRHN9umChoV5r0h
ZlKhrf3j6xdor2cJf4SL2rchlyiLtcbKoaVXaadoLoiOtY/aGkgiGqOmqQt/c+wKdIiORMOjX3WW
ZTDFfHJailjAa/GFgr/g4E0vju3J80RVuG1sW9LVmTj9i3HYWDuBk6qr7BUl0q7CGYKs9cLMyv3c
EhzCmsJVulKoWVY+Rd3knBrPLC1X5rLT/25FdbSG/FpWAY6KIgbLjLxXKuPEom862wHEcuYNuSIA
lnKVS95SB4DSoEZGBsA6sdqGh0kWkCn/BNdYljVE70YYpG9AtUVp2DuHelx6Fiy5rRyCSar4NeJu
m3uOGDwQcsoWsav4gSdRs5aS2LHMv3Cjr6vGKMWmoRsrG+mNuNfPAmFtb7npmmnU+w56wOCjoRyR
U6b25YrifRep2buQ0qWG86kDfClRmlB64x8KFoq2uurFEe+ml661UTa8USA3Q3fM/GEjj2Ntl6wW
O9iDf/cCcjHhnnNdS1qlqtVplgIQgT/R1wIzWVhPYQ/8WpAdjKk3xaekucRCa4LguipqIVBNi/DM
47rcQd14W05BgnBezr3Cv9Wj5Uqxa4bWJ2bwYta+CF8MPqKkMZQ/QQhXgivCS9l3E7boG9RlEFOt
GSoMiKK06xpetBVm4GuKoXczTuYaHrbYwAq2JiWw673HLSJlJ7zT08UzCwNeUPt2l9pgHPVLfU+P
L9iq47L5iRF//3kiNs8dr4kOW7Xuqdx2mKrt+f+laMbbINkGzFUwRzwlGqb+xUZ41/Y0nrhLS85/
+bTACoA50HJUgYf/etbnnzjHRUiUVlZafzaZYP3Ymd9GueEvnGHbVP286wQjncrg8lVyxjedFeSF
QqzNpPa50zcBgkQhmv1NmtnqFcpT1q9scOVvU/j/sx3uvxurPa/YyTabp1Ro5uLYE+rpWAgQH1ic
tohryiGg6th+1ik5wAecHIxPYx9WVLbSJH9eeNKX87rvuLeBC2WnHQU3UpI2fWLhhD+nIjcRlEoC
N/WzX3K8O84XlRWY/ulJE7ftgW0VM0w0EhUJr38ELUtuXm8b/fVN9ClGUXFB2vUrSFw1rikVd2ax
r6/QjtgskmSKBkZmvmnOvd8f/bflAyEUyDSR6f4fLPn3cm/Xb2KS284sL0wRC0LH+29VdyOU6woT
PSB9vpuauJzUK+Y+u45IAam3Ypuwu13PYTMlNP8AuRIgJvEWJmutO7lEADqDa/43lS3m5oGUJUvV
QkcL5L1IUtv7Qt2iO6TxPJm2dFea+d8QCtmm2RoyH2Xf7ehhi4vz6XiEgqQKVYLojZ7RRdJWTI8v
QpDK4lukEymYqGiOpS0Yt+HVwTpcnaUr5pCzmBrcKWo+Wy1RlvgZHIu/mbLHFT8ws3SJ0ILoYIYd
8D17TL2ttmlUnYDpo4MnuS0ATu+oKUde/7fr8KZ8n3meolStxsoxy75smM5emPpoPWEERk2QxdTJ
AY63Ure3f/5Z7XGJBaDomAmShkaShwubELdt2jWjnFv1SezKFTwyCq4o5r1s7j7r/EAbrVpJK1ki
kEid8OjZyUe/iLgQ0QggpYB0C2954HsTXfKcoX8efJaKVuzb1qiNkHo+z6dKLsBsAT5M8E3KCTzE
hE6J1klgvZ0/Us6eFEoQBalF62uiiDoSgZbTGoZMT5wO2JlHE3b99rUKmxls0YTP/RbhynmKu5hd
D4TazGolJ00ReCTM8M1zWfWPD+UFjP9wBIf+D8/WnDBmaNaxYVokaAwR+n8gnaKDt/HVYt6tdfxO
Wojh424lAyOlMQYvxeIZ7lgDqsWZ3Ttt1oKA+7wnfvlZbSM4GwWAbyB/19bTV98rptqtFe1/IBIm
/C/XqJaigDt6I8vOvI42+E9I+9sYuUweWr2VIkHfsNCotsL39nvhdYqj9IKcJLJN4UTqwJ3u/XB2
VfGvIBwVd1mJJy8JXzu7fHaGFvlko6IkZjjToVXpAsUbnf9qfHRl1nNmFaE7zawqFk07xe2LzqJ9
XdRDK76bChgOQeJEY8YIZnsO2ye0r+oQkWNSP4i7CZdVN02ANHA7U4GwaJ6hD7wJO8EwgbCgd+td
4hs+K+gMOHDfdO4HZv8q4ZZDyQv+HHcigxPQGoDv431r+PgpWZSMsZisTFJva7fLnYQw+JhoVSSA
rZI6GCqgyT77Sv4zk31jT7PZb7TUBdIcPV/AzPDhO09C76tFg6YoAyIF9gwZfHKCU3KGa3uhAGHd
j3I61PxcxXuOzoWYtLZJne21u/nyg1h2otAnW9N3s4qPMvoRukIiJ+UwXwP3IHomjCcWci888sXg
JIYDvIZUGAWun5J0lLwjLgQwuxk0/P9ywRn53fTit7biP/DXdTbqvW/tfUciAZQIhZW2z5HwT/AD
jeKaPltkS8F+EaIZhPFphL2+DpKKzKY21zs2/UMwCyQm9Lttx8So3Xw8mVi9tqDjADamUhPbaRXV
TyDaxj3SyZdpoc32aN7b4yhK4OhHR4lVajj0SXfjc7oGXqabf64bUITiMUlMYNOe3vBf6lyCM/6K
FWpzNaUcw764yff52bGIkc+tHquKokOlxoi6WuOuy9WNZfh5dn3XO3O4wPkGrFQc4s5oCAhTyDoX
afSmjx8CbVAV1HOui3p9UBThMVeUAEt0sup6IqDeZFwRpu611L1g7CRDW7s0CMyuv7UXrUwUKEza
pwU1A0m7lrqQYgPldGjbcDVjhVl1lsuLknW/xa+crrqrMNz/w3eqXQXA/iPsgDbj9JCZUiwvTQN3
jCC8gzSQmFylu+OzBgl1iwnlsMhGX0KrH29ijl2nBHXjRubH6C0ICOcy5EKR45uaDf8Ftxt8im7a
5nVQ28kXtMiZ18l+9+WUIGzR6KkeBqr4xJRVoSwXXO/OFoibFBIlq+9nk8jpJvolvlhKFDTl/pk3
E6HsoZBbn7efv8brSHVLjmr+cv22Oq0kRVVMY5fFcPI5WOgBWnSDlegwZzmnfjnBrjA0fdCBw0eJ
mM3sgsO3JisLODX/NL7y7o95niSunchbtsMxfxKlvL98Bqub9vUJ2fLjHvHOHTltC31nD6jihHPD
r5VOtA8w6+Kx7ldsd+VYpHZrW1sLrrxpixOEsKTAK9vy5s2kP7idndM+Sbp0w1jDy3JLlJM6NHjf
//84loblLHHxbwZIDh8fkYjh8ef8PdDrZkIYbbE8EPgmB8U1ZHx28J85FX/bHv3mpChpQb09tvP6
K6ef7TTE59PdkGb8s5rIcETGW5kiZUBkQLByWFUnY4Jpp0gzIt6XrF/dkU00IsDz+FYfSDqsVPcG
gVhkG9MA8MYMt3kcjHN+NKeJZT4XofLDGKtP51WcipLDL18Adx3C+i67AHhEpNwrpaNsPaFSpsd+
yDQCPuWSWaouU6fxPc2sHbYoh3lMBVu9EGzKmCox0dTKxhTRamoiNcZIgYX5mlHG3FBcrKUKEBUH
BAt8DB22Yt01Ijct4N/mIOZriDpOmfpGxTU38Y0yekWtMiVFGyIYsCvC/cgTjoBWEV8q8A6Erd3j
LLP7LDTX0NcWDv/IdcEIlUGK+cGAX9JX28iCNVm9JwFI2/SjkVwPV6LlaqjbWoAEozMX4IclLsTY
TvcXTw8eh7UQFhxlNyG3zr+FJ3dT8owFnDSFCKHfExrTKQgZrfLAVPD4nDvGJes8NfyXuDOXRiD3
+pM+eOMFFiZqWhMFGYqbOEhRiVhnEQYOMUQsYTrHkl+4RUr+ngoGbE+W1DI3Zgp8kZZsjPVOf4d5
wtYabaGE1N+uK7TL0gjK5XQoMv5eeTomEkpWi94s/RJMcwqipVFT8llKNyflPMbg8tW08xbwdTN2
+jQuPtBX6Nd4ydyhlkOfMqVKIupF+WKNMfnLFR2qEfqyDh5u8n0zLOtvz8KrAlx9ByjZyAoKkKdO
wUnCddmRGHsEThBceBQc0brOQTsFxL3U5gb26X5kXvL4lnJIdeypZv/C0P+H51C4bpq2adjZ0vsU
hsjSQBJh3nGFbb4fEuwLG9Zzat8Ndp0h9ZFnUeyWMsgZswssjqjzQGstg0H6YTqzluhZMW6gy207
BGPqmL7thwFAnY0+Tp2C9RbjuqlLUAIS+5H9vJp+eijSJKEsEPJBQbHgD5XhAV+ZvWzxSadTGh+r
rg/xLdmb0ZeviRX/7OfMSk3k23BWess/JC6yzlUZyhMJSiSqJgrLpmV+Jf+Yxkcgs/gOwG2ha3CT
2nQo+3Oi/TeMjxF3QGc1RiyjEOyObTFOAS/ZvSw5tMy+0UNyUeCaRdzlmPJDk2A6lisr45ZQortr
g+Lvma6ZSM76fZkUweAdNOIZOZV+TxfhF34OX5Dmi+7cphJ09kCS5XDh1E/rFs7m+YE5BwNDatka
lKiLS+ctJxhhiNf1yEKFwlDmnl4m6HYO0qTwVIAE2+wHQhcuv4I9b31cXAnANn+EWKeJkbNbjnsX
i6S/ZhDQXeXS5p00OWtw5Bl2M4o0hCQXbuiDtNQaRSO6+ZPrYCw2mrFFYG3RtNdrPSjZSsUAd9do
69e5lk8W8XRIHUzp3vVHL4TyMq7s+BaJHlRTmbbpWerOZgXXTuegQa8Jf9qNeZTIVoQm+VXBH58x
5T9wY97ipJ3KZC4ErO1DEpdyXDzMXlu95OlPsE45CJcowWg2X80FK+DY27Jj/a8QbEYKFEegfke5
0uyza9yzxnXbEHMyopewITu/h8lhP6TVBGQaE/8l3GsQnfBzcZx8dYou/1d7H+j48oCk1LQUaKcO
lX0D+8NBhRsIVM5mX25oXitwN1nuVzXP9Lq3Xwq5BPWrcZQmBFmKQv9K3taN5g/b3zrZz95foQOn
eogpFXIUF9r09UM4fahb/TNoYWko+QFYzZ6r/HGdB4N0SG0Ldkd/GCrS0U9NTYip/ik22IA+goaK
rvXcYjnTvpAnaqCsIiUzgZwNTl87JsWEJhyzJgmvCBe05MHdgzTyTsmdmCp5yydxyoGbe9BSw9bN
nC4bE24FRcs9jpI6CINR1lbMZyVoTcES6gYvZUyXfBjqzI1JlesUerwopKLEcZnUHOdT85OOQMVZ
X4TT/lqKRE2HIGSFNnGn6gKWIFOfOQR3zQgpV13HDfeoT8ybSAQqPrZl9tgUjpGlswMXy2sYIeSS
1AB7QluTo8TfRGUsxqizCQkvdMNhjzlbQfW/UDuO95S8Iq2moIUVE3toY036wgc6QYcUxVZj1Q1P
uYoZuDMxyP2feh9QR2fsDGvolimDxebo60ClcM/DUb0zH9R9MfRRL4uovYXfgEr3YLshyCr4tzOF
P/vK3IY/0DrFPMN/O5RaL6rEi/dH/VxO8ijuUnW+fNh63Xn+E4KWFbk37gxd5JSVbW89/b1imxxV
RiSgHhl1dPyXYgp+isXnyDCWeB5dE09z3QIAQSqgVObQLo/yhmCguIZsYqmMy6PmxXJrBR9SfSWS
f+7rb4i1wMtVRZDJDXxZBVNA7/XMKJUkSXpJIDEfi6fxcquaT+PobKo8QfrVV8+SwRgi1LaqU8Ew
ziztW3gXSxTbmOHwe0coLKjajFrmaabnaKOvmkYZ3EqyhOi4qjr83IWuK6TLnA4Ga37chQV4dYpj
MqfopaL/o/TWNUYJBHw3UItGn+rYDnxUTS1AW9DuJOzILduKMhC+3/qCbYvuSOw08nar30wPOsz4
p9ucwNpf55wWxQKAmDs7/5r9i/MUNu40Q7X8Pq9Y4yskmr+DwYpjoplP6/DuM93AO9WRCyY3twbi
K2YqTFVuKEl58FnmTWVu07Jh9h5HhMVC7rIn5JJzTW5e6in/AfnTsAd/lMYm+EDqnNMmlPgIFoNs
7bFUJ4H1h9UCsk+RWpvjVxwnAPE6mDsyrZDQaLdLUGDqZ37yjbJsHT7zVJZsHou1x2m6WLMt6HUX
JCfxNgKA/OduaAL80IZp/gawF87KWL9vpLdl5fkjUb46/jERwSs/IGckn1h9/pn1XHJmiaZlvzlA
YfzxtZIU3WUIM4YXuuja+HPElmLmquMZWRQLkkc9TWa/ZL8lE3yPzsA5L6f61faLV3U7WuQ2S4HY
fex97TuDVsYGnOoWS9VCCO++wrmaZTF0TOyDewcFp3Kpvgt+XH+72p185FTlGFe7D601kjS8zHdT
LUzPdnMlaL1TzVBTnepCuUOut8auBJGoNfKIRFkOjZtJx4Fpf1MfpYP3sXM/tq1ehCA/H2jfjByd
x9LVmVP44tAGl4ENIjxdl6uUvNVBJ6POkYUQUokboONEZwLYQREjlR+PuV//VwaBudXW4Rk1C2s8
Wu3U+lIDtNyZpyUPDACYB+EYRk63BwPiDqpYSyp6W3J9P440CwSzrfyToixYq7Ay+/HyCagVTp33
9juHY8E3IqgcxzVMagCBFd2hFWXL2V9j33mTdS6ztoBKvYN1p2UA55w1aAE4cmbKQR6rFBu5ITh3
dZ67l1wVXQU/EtX/fAwDi4/fwPxVWI9wn/IYt96stYIj2uWneMJoq5Yvdinybdkr9IuKtd7q5jCg
qXHIUBelS9anNgE8BiuPqWqwQ9TM9RGF5NG6xE4Re8moiWtKVeuG/+Mohg5xvS725yvgpqoRHzCP
HFRNkyBmShb7gtaED419l9+bICszPQBhrzufs1qdeXFGrNf6pTSBEkh61+OnPecEnmC272IhGJnr
Nlw9YD0uBusheYC2et5lleNwQZyLmBWhTK3gMHgRwWKyZHWFWBXcfDq397hLjapZVUpqxvg40Uv/
3W4tVR8D/dJ8Mo5Oa2hKytdi41AbPteSX+vMh5a4/zKWEFJHh5OvJbv84L4ktIGXQUqX06/ha9mz
0teutWfJata9Q4vZhiIDE6A5RdKDtcwHjyIr2QNwK5tAGJvOPsy5u20gitYjxJ3v8oZd3zUoOBmY
uaF4M8xYsg0O0Azb/mQ26n7sMYyuI+QKVA41G2+i3MY8VSQQuoaqU2+WiledzyUbt0VeppJOixo+
L9dpwkuDdkPw+9k3q6OhYFIVHCJGUPfC5cpURYTYkgBL4mtMLONvHMVkaew7qm0D/1AHBx025imq
X3IQJ+R3xUU5+Lp0B36CDM5JjkP6nBnkMIbY58ePebywgEqWdjl3mUd7p5VwR/TS5lYNXA8nzfUF
gH4RcJlCiPPldSq++OJ18Z25gq2x4v01K/CFFY1lioggPlp0xoF3kJ6b4bNhjm48vuSYDjWl+5G5
a3KgdC1n58JBVHygFmp6XrGRX76q/v7QiPpWGpyCTg0upqqpWBoacniDYcntzLv89tO3LG4wbFDL
JWo4mmasmWgHpjByaHYg/+uX2ph/WwlglZ9xyLLbm/t+V/hcU8+UX996xc7siobAoYiMAFSnq9WB
pcTI1zotsf0z4HZ6AF64WqTgz+zpUqBzxUP3bs9Z1chh0qex67pHjRFwv6fTJbyofh2iVE1cyr5l
qKTxNf2lBbxdnmu19QpfvhlbLZMUbuuloX49K+c6Hv7lJNDkhny9fe+oRz/snJ0AVcX0dXaap90D
5RgQ198Lo/8p0uW8c+rgLJv3uDZ3hyesA3Zw/aeecsb40IgFZQtjRfLe5gHrzgQDteYcu0MOU5o0
2eNgjM4SDidE2tCHt2c1Ks24HoXn1NsjHpLixtML5A5jx49LH7WzrPcdyMhuuQPw8tEtbUjhtq+Y
FnAdPi+Iu2Aj6i2txz472cKMwafusHTs++2Mphx7616gj3ajLmL3CN8ux7yjV65+iKIij6F9GpU+
4flvY/BP8yBr4qYvEOXNI6q4g/hPIF1IOID3o2jMKh0Dk9V5AJEnJmAETPrkRJxkbTCfrjcVBoO7
sZU1dfdXTSckc2I15iTZlTXY7Qvzdl1x31A45YF/UzZiuZayps112YBfi3feie9Nmt6Wqzxvhvqz
uFQKnwEeq+HqKrJwqVwEQaa//4heUbUkn86jApu2ZNht47eDS/VAl7r0Dmx/uMd5DijvIoo3N8R+
OZjG+A6nmsp3XCQRe4JFM4LbXKEiyYEQAo6qDeRK8eOScYtOUGi/jCiumnJs55rCq8pr32f7oyj9
UENWZGqvK80aUFMLjit+SLz9BDO65cOXn9gz3e7aOzmMvtOaKaqZ9z9X6qr3t67PROuLb+HQgcaU
XfEUrIURg9MmuRcUMTsZry+1de882XLQWH/cLAvLCm458tXADuPlMi5ukX3VeZlXv+g/4eZeoMIv
CpQhD9FeUNQK2YfNZGdTeJ+zmLr+z8qaTBWdII/wWp5bwSlK/DnoWDyX+QlhcijSzpR5UIak1Yts
2NXjE7+Li0MBeQKBh0C0Yb/45mOhjRIYN2Wwr5HIPBElybdZgLwVrBGggBxBVprRaJchAYFxeb0E
023k0y7OyJLJDJ2NomHTViQlTCnifIhdedGWDp3PX7OptkCy1uzHoV+8nfDBxm2cjWh+FcT+vnaO
Cwr/cBpMfQkB1XqMNy2ZQ86yKOdQJwqmQWfUzzYPpCS+ikZC1iIy8i21dtLGisCxWMHePmYv9oQp
67Djou7AESnthBuv+yvNZ3xIsfkWyyGQS8329LyjEGqNXmKSboXZhfFlEZBOzrS16UWdgGKgMtNL
ac+/BHkpCA3Jn+MrouKM3UEk4GNsyHS+XSYlbrYAlDZfCu4XawRMt5bnllTsAetPxUO+hvpTRW8A
j/4KKg3s2hCC8dr0o8zaWmrpuT3MeTsT5ynVvrh7VuOC82PmBXlUqkEJ/qDu/qS7Aqf0lhJZLrZK
3ZKHTbnUF7EvnsgYAKDuWG1M30+lF1fEhCco32XMWZmBSXSOYifkDwhwbDqylDCm2zlbemcn3rMz
7p2aaVTOA1w0zZXK39+RRafEbrHItRD8p2uEO92/tMdWmkXrA/7BprnE3Gpd0UYH2cPZ5BUorrJ9
lUrJS79XkXIfPRuN3qbqyi7OsOkc+2Pc79vA89oXs+5f1vxazFbd/hdcn58v5ouVRNLVbLuzr/iu
e330V4kNpAYvpy5FbPUII/2v4QB0dcB+/b5kNIqERzXJshxutcAYtwdJ4Yl8hb4MAxJUeEY4J15v
9xS1dJ3lIToR53nctLmPBZ5/IATZ1/tIPLpYyyTd6fZfpaJirgqctIyA65IJIH8rPYWkLbH8Pyfb
JOoBiXkwreGZv+tC454eF49kyQNczUqoLWgAh9VqOyhJYzsIzuWf1S8FkWmDfwOjxz5TtbTfwSIX
ahAs9IVtbkfoFYkp23cAfeHp/dKE8A64SviN+/70jno8f4bPScTuhCFZEMQlBC1ezwd96UO4javR
EJUqIlfoctfnDsqa+Lod3jCg2XkjgbffzZcMxrMStKGbEIAhKXlps0a8KKwU1OlmwfrssMJD3k2P
lvzPlJ7JAZsHt3GXna4lSS18BmWzHWsA/SAUjAMf3We3riRv77DaadZlmrf0kGZvDGXodSh5QcUh
qN2pNS4mRnWnm7f/8OKfl/0JBKddH4S/N/el3ijV8mqkode9R6U4rDW2ysYcukYB+CMjhl1k+SX4
eFs6X3jxL741DRPEZNxACQqLqa8yRt2dcOSTjz8vbHge1SU4okcpmEvb9dEPNNWLP21DkBU+/y28
ms/5yrVwLeqq+PwUsQNN3X4N1QMYh0+yAwVJWktiTCehO6O2JVY7K8kHjw9KLOgF4nfdKlZxZP84
ng63b9VkJtz0B78nOsZaRpJE676ZyN6g8Y1eW/iRt/hpDtZ5Kzz9vj/uBCi6zIqEb6TX4BYavT1F
JUgJKA9KuSRCeTsU7pkZsOt5Ix7EJJXHHaFw1zd8l6osQWXTzcXxQOEr/5OnrauFp+1a4xtl8c5/
u45rDDoIQyucZDI1KZmSzA0yH+/wpjPffs6tPwoW8zfXtSaBxEo1hmulZwZ8yEJKQu08ocO9q26i
41Bik72kbFmKywUbDIsaWQm9Mds9OQQ/iCBqR8MZkFS2vH+Uj5Ny6znsW9Pd0s11APzy8hbBettF
QLvjYVpUiFwqo97yLdiKOwCRTZbMJLrPWHkewrre+pgZS5NY0kFzUIEoBgmEuTZ3fqIF6fV6SfNv
ujS8wLn6ZI4Yj8D9Xj/zA8+qJK5ZCrKlmyXtMNEW6DHhMNINkWDgpfoRdi7YpUSK7M7Q4YNOsahY
4TzZ+ngZ9sH+il4/X/Srdis8rmUKteEjNPQp1W0uBQvTtgDFcgdat37utYM4Wv8WafoPaQU1EOEz
4h6gsDUMofxj/iYmxS+83k/ClgZj3HplMX2/lSdMYytd2zt91yBcDZQb76HOwUZY4mw5tvQkWIWk
NTv35Vqwvllb2d/vgo3nfVEpULve6SkdwFn1LGXSModV7KK5TGFRqrz/7BEPct9xzOHzCssVMlje
Fg1OLpAzd6zcd4dc+DvgUhgUuLTjHsKTSWH07RgFYyRI+nvWwOSCv6Q7Zjmqb+BO2EX6hdcYFV5j
HPQyE68UbGGMRTy8Qrn6/KKedakxNX29zG0b4s/muf/pozD5WB+bK8kr1yp9rQG43XPILOeOEWgZ
E9rc7YUBRbeaPMzJnBsKqWn1Z0B8fuiDfFD7SgcqbQsYF5uFie60CHAk6q6IyFG/TqOFcMBS3dxg
e/Oa3Y69vgh1cSpQExm4Fqrc06MCbtpWbhmZbZJW9LPb2mFcRUx05QymxpQcRbpIs9ceJe+24HoU
T/r3q1GDtZnlY7Dk8QUvSJOB6zwbwKbKJfyshaYfJW1weTrpys7ix7uLdZOHKRdZgCAJprotrIlp
7/x8SOjK4R9kV+9O5kzWEe7wOdIVO3gdo88Xvf283snFhVuenpBrEGSKXrqNzw0FPEuIv7jmTaNc
taXcpWzC5kMt2nIMgzW1DHW+jmGrdLZcT/15HSQ2NS+8CekPJdsFLm2BjVB+biYAPLAZ7LN/X1bu
kPwNzKD6mqgNjcvGt/PUPhJbC6IW0N3zHciEMPUzVOb/Qu4u3bokF+zcTMmkzc35gaKeyTjtHxKQ
y0LLJdyG7dnvEpDWTBbcIwbpKdvlRxZ9eFotHC2J6o7oFXTjHFAl/9j9xhs1d/QOTUn2lLHTZGeC
uVLjKCmuPtG1deU6IQfZaIDsSSj7n4jc1oZZOB/uCnfw6AzDav1/EKEqn2t4thjsbTc3ApHgvNa/
7KfaNvCVaaFmfdXK+err2i0Uriz+wGy4umVhmolA1lIddDWIBIL/2rIKQ2SKMQcOzyzMKJy4hwcy
maMjPqqermOPQ72k73Yrmby371zO+Wo+GkO+zuwzGmu7WqeYURY7VHwojvTBbE6pFv+DU/k3y12K
9C/mi+dZVoxjwdmaHzlY02SxEQCZq6n7dCMlp37U8hBpWGwI6zYbvFkfzXVGqq7djlCOakyc1MNe
BfoOlIFEEi35JFn5naRjNCSDZPwojfsR3PhM+mkdfaPD8zxMdpseJyfBSqbgh78X6c7Xu/fP0/OL
HXtQimYlbpu6pUF/NgOnfONL+huB577DFWH/B6dVWzJS2FtVcJgHJEgVblu3rGdPDr9rfR9mcYie
pWpJbHbZzx1G2CswCTPTBcQUy/P974nGEjZdY6x2podNIfy28OZEDkVnAZQVHBUhAe+BkySPVvzx
n5zxrqONcdVl6qp//r0ulGB43qEL/NvJFblUno3u6GK6T0BtIX5IbfhvUa+p/uP4nMDvF3TzfbYJ
7eMBKXu3wvY8zzyVToZhLeuY3bE4r71h4Y+lUubLMyZH+sJadX3B9pD1WZ/xLTEY4wzW4JP6Fy6z
G/pU6mCw8toIUY2caLjImZx4cKmOISujMkP1/5ZPxQ/EPaD5wzQj91TSI9pvXfLxCJrF2bH3GHxh
WTBIl6WfcvjlkoAeCe97Q/Nr9z+GymNKBKYK7F5HZpKSPdPLr9QEkY5TtOMtd19ywDLWiWwKcLOm
EtmfnE18YGsS3vZxddvzFP21Jo32Wi377Iaeic8By9guMNWHY+H9LPdxyKD1fm9BFWQi5W6eK8XB
PJCQTsQmnUaDd1AvU0CGJae9+4coSixMAjHkVqfL9o0ppI16ELGabhG8UNGo3v4Gbq95+Bg1HBum
qxS3wdtQteuM/zO90lv2K+oVZ4O7F2NU08pKn8uht//asY7Y0iVjNi7wwsjxgcisa1+JK0O48lh7
9kx0phkq6Mtcd5OylGbzcbcJf1m8WSxwDmUkJCdSWJGgsCo8wH9syRSfnlimdrO17X3OTyfwjyAA
WpmuY2xKhxMy70kEDXzRFjUy2Q9zB0XsVt4JfdPySfkUmK4bGAz6KjPmCuQxoE5glDOaUjc98rpa
HtVQ2qmsKJB7YxmHRE5uXATkedZ5+68lil7hlosDHVlPxE6WhX6xTQ3BBnJhBqdb0BTaiCwMCEGG
kedEii9DthtGuS+mY2X2jOia+a9VwRCHIsZnXGneT7ofQ71BydYj6rrMIlbA+hQrb4utvlMiRH7/
9qjdEnCrXkAaSYHfFse+HLByg1wptEbmpBUHFIV2Ho0Szv0hwN75+ozZmNQXx/ppvRlPcyR9Q25R
Liu2X5TOEAS/rD2Odhhty9MSWVLmxPliXHMrHBzfC4kfIAycOQJFLzJw51klRldLLVJ5rmpbJv7H
RdrVi65cYEhFtiRJlR+GBLJbjOo+CYVetbOEYEePxjQB/XE1Q+OMJ9KdPYMfv4KmpSpYRbbX25DW
Hitu/MzA42LSLH2iQJ1GqBLTg8Kh9HzfHbIwQ0FALT/BsAV+sOHRiwV/8Zzq5+91bxR7cMo0YyZ4
w+QZJERzuT6Sgt9xJtXDJtkUYxDFzspSeLIWq1RDxNtE4jFXrf88EEl5tp2swSWUpKFGQdWZy3dT
beIVUaBJWULkrV66bWOshbB3olu0LYPPU5IYi5m4irCnCHbM6TJ88cx2mF8pnrDrQuvPnqPCsL7Z
VoOAJIFrSF4lKE7H5MIus9xNRETgt4BxdtqwxoseOr3OmTQ+0CPfseMtayBbn5Pa1kXD9OX90xGX
Wwrh1kct6UXSlSjlaoN8ZrlEqVOGVMg6ONsL+zctbQcJfq05rLFseu1OdL4J7q4T7H2nfAKMzOkq
sT66YeEHExoOrLnP9NK4ltmTmr2WqtKodY7B+q8MaQr//kCFRQadyLSLttGwEvMQlx7Ddb667nwz
htJp8mA0OojVNBdO/MMgNZGbhnlTv5JcoGBJXMseUmCBQf4NHGQosgl24T5i6+3t0577STzyl5uo
QaQe+uQbzG+7nSXzzCLw42bklzBzT6lzN96Zp6/jOus9oyDlAsi4Vv/ffcsExrYShZide2LV2uUd
3K0AXBfgRvwETt0pnfa4akbAmzZyf3vid/WsCqufPEcX37admd9Zgub8Igh9UrWn8U2/twVshhUI
53b1F9a2ZkfO3c9hZYbsySlhb9LvVvQjYcFWfEPYvcym+ke2Bxnjz0vM2kmHFBWoUy5or2i4SVZA
EIGzun4T8XJYt00RvlaN5dsVrq6R5jVRY477wEF8wwfjVC/AdzA5PB+nNUfa7X+0VOEtVxiulL02
sF0WrEVE8wniE+i71TncsbLEYdSjF6X1AKVnGgC8AyKb5j6RlyRlGiHVbevnqvbXomFQ3gt9iuwC
WZa+lihTYvPyf64gS9gZY5lcWMI4skQfa5lvr+tXfU2PwefoRffOQdqfkAKNXUK+5rfS1N8Ph4H2
B6dDaIeM8EkZZPDWb+bdYW6+YpPPhjhTJ9XYgGqYdJPXn86kJxZIpkLImjPfTffNVucfr5ozWIkL
Gc2Hjm/oi+/G8TOMbkKpP/s99BydhmzrrAQuQAhipjhMx7aKrB2+ibJuN0DPLs0hDidseTwn9kbq
Y8Pj1kXhG5N9aG5OyL6rNwNKdOgDaKTobMDldjKEdhxdov4LVK04QZYyN3oroYiUnXfk+cX6R52q
/X/toTAQJZLLAiUDoKQoaJJyW+oCd6HXI3sp3hvZv64+xpRHRt5NBN1Ddx1tKhLbhqCeQA7AHu97
MeGEfk3B+7CU93jTyXuGJPkFsmuKnkwMTBkoRegCZ/dsGPSH04pR0rOKZBzxSSNAAxo6YQjHNhCQ
COyneNqYujJQVmShAYVMQ/IAs7Bg0hnQyHOnFzszKb8EmAN08J4F2F9hI+233+H6ST6TPptSwJth
M/NXiXqT046t/72v7GcjNgri/qk6zFfUKBUpY2F5RLnf6y7p78jjYdoAE3pBTGBLd7EyieS/r74t
M7PXkof5y9iS9SOPkMa7gndZYfDTd1ofFiPKyTae0hryGf9IISeV5OIWP9qYXmPoNtlsOi7x0Uhf
XHPB/TaFNo+kDQappTO5HFuplC9KL7c+497boNo/6XgAz3SpkqOhCGPx+jDG4BXoxCfYyMfr8BK6
tD5iR8ByYr3Dw0lsLUpUHqgwcuJuxcdodyRy3V9gfILAitIs0RlcKBNYkA9/vn6ZqWkX9kttFu5d
uAgBjIBm7hqQG0FSY6cF7Vy56QQqVoc3qZ0RP8YHUl92ltHaRqcSVP97cmNzf5/ulR+Q83pZAWfW
P0X1V8VRZ5ouWxdU0KwuTxmu2bQXNHzNTmK0d8gme6PrytUufNb2U1O8Z7JQHszt+sQIaFYDf6+P
ltQCj4AF2XQOsEaWz6ezJkWiS+EVbmSrAbkgZIWv+Zens+BDCClHnFvpF3PDkUZStN1ewAjtXfw0
5qbCVc1YEowXojU4qC52xnmP5WGNFMhpN8GFkDp59+KYg988jyR003QDCRXGzLxrQPdj2p6IjfrH
SzdMpHE+HsTtZyfo2v37PEhqsit9Nsk/J4PZMOKRGyEGNVpy/d7tkUSKp0iLjo9av/xEFDuzRUsw
ng9xe4UIQvQjgJyC+2GIQheunkmVLBCdgikJTakXOflPFGd+N92KY8qz/hrdk3saNscZF6JeWGO5
lhLNYZux3dEcPOfOX8MEAP7mxch7Cr/XrRiY9t+ZadFx1pi5uqVKaimxb+SDmAbxci1ivri/szxO
UXBrtbXrFF0p/WM9LHM8UXXEnImWuYahEwPj8s/hqqvj9RhI+XYptvSZLhXzfTo6vRX6RsxypjUa
RifNDL65U8DaGtOsbrpzutaS8QMItXH7DMflJ9pBr/PJoEK7SlOqSEViREXb+PCQuKfxrFl1piPx
h4+pNiIpbq55tJo5S91LvMjovL65UGFfRieakuBu8ErhMqyBCNM2GonNH42jOu7C28ttPzzWMS3l
9i4mZdZv4luTmpnPxBePyiqzOoqSIH4LVmI5AaTw/N0N3X3O1lmP25BHRTgNS/5RSox/bdOLJx9q
yU0r+mfz4mJ+breDXYbVPB21xpLt2sz0pVQZJ2d7Me2OhMuvvhM4f2B/A7/0jqJksEWdhP0a01YH
lgQlwYJLBZYu+jBGyz4AznJTJy2/PxjceoS7iVlpAINCcuzmTmJRtS4hXzGZFNqwF6yBD9Vof23c
svTZw2RUzdVZyM+6T8q/xsqVnl/l2stZlLIwbKjL8+KECNtqGjiYlkoT8VMDqBehTlOhZJ+5pYPo
jhdR3gID8A9NDlWhQU+fZYnTlaoROCTGMNZ71n6NEMOvQWRl0ARcoGBOolc+tiwXRFdDkt5H90X+
1Qzi3RkKqSeGAtytNIWoRYUIx5/PR/Rjqhqx3jj7BX+nHWouQ5hphWKGdXvED1/gnYH4c5uJjU+h
Jify9myGro6zQbXVpRBY5jD9Q+KmWixnj0IJDuVg/HKC0JvPe42K9EFWOMQDfpl7ri/C+hVWEu6V
EXSLTQi1lwJ22Kd0bNS06UNET9X+Y3ZqX762Wk2uTIY66hEWwDjkbsNVUEOxFzq73MnPvfTVsQiN
OCEZRF/zPXyzk4p3pW+E5j94jkd6I83w7qUhj2kHrKEeEliXmf6ur/+L5wievNxid7+neiFjLPpc
hzIGgy9sukJw7/Y5tUp6VQ0pPruvyYtAZRNlhmml2qvAAiCPVvTU6VguAhPQwGhDHeY2qINeiyPi
WJxGKL4zZW6eIF/8XLDw1as869VKk5Vq+197DiY/pnThMHhGzKCVUnZIppDxR9FEzQdymZNWAMe4
kV9s6v7x/N+neMpuPEuvIAa2fFf6faUAjJW2R9pcpQ3ISJYVfKBD1VBVOJrhyjDky+YVTRD7MKg3
4l/fXL6ftVDSUl9IkbGY+0L6S88BKKpO6TOzO2tp2iDdhlqkD89GnN9reMYn/86FTt8yBMUydkQz
ntSfoelQVWxIihX3dF3MpUh1pWuuDP+JDKlXbbvHxjh1y4cTIl1acf9r6e5RK7+PgQQ9a6ER/L/T
NOwp6ue6Hyyv6l8ZeK0tFWiBF9Ek3bqPHCVLh2oHN+FuquVAQa3OEHsvuHhi0dOkDoz32gcFGG/i
jhkJVijlGZnl7cz/mRTNjS4agZO5G2TI8l7l+niznMwYKb/hK8WfWqCntXPfUg7l1tCGzsEIITCq
T9WbzkhpHinvrG3VGQJVi7AWv4C6hIcIc0GHn/8QOAMiwDh6c5YeAFKmiMGbyDcXc/Xw0sT7yubK
pOskAGSKQVWaRtVp7gq/w4Ru0jwlRO8sSd848juNcRDNnZucZaSB8NHEAErfPBpGFpkmuT+M5ZTG
TwLXEG9XRqOW8eeiL5xd0g/btuuBWjD4v/PvrgN4YeTwTS/GiQXaUE4eVkzw6NHXqdrxKb7tJMr2
XRhfsdosp+ejuBRCxRvDLNCEOmoZwxil+vdloqvtGSkOlD3X5t9+xLJco1SqJEgeoNwyhfsNLGGc
pakKAHUp33ymU2ZRDRzD/gXUFQOELnsY688D8yTJ9E0DvrzRyskxp+sPUH6NlOmUb6UzB1cmhBKD
IiPqeZOPAws9zdWIiz6ipvsiS57/8nmocsCBOAPfR4KQPxtww/f5iq7mpOZBii6I7OoHx7KbMfsN
URo3Gqrznz5phdhbxm1AvfmzSzftDnPafISBTJQDlStHGes+UGx+94hdSB/15B9F/Rkr64w0XyQ1
+M3R3N372yKDfvbZxmZuQiGLQP2TPU04zpTE7rkJ/ze93BNzURCX+7vyM6m8xDk+6bdRCt1u4i+u
fBOU44QJw4vgTfR3B0uuPg6GVRQwP0fjeNfdZRTW4w8NHErvsGNChsf/jd4Rh9c+0/8ucB45XNWk
rUxyMtJ/QFlJAHdRgMKQR7dVeV/dpkeiAoGTx8j/E7eXxnzPpIob77CggWZTLSEGdnOf1vX+uEJc
bWkAfUtKZIx/v6QKLhWQgnYkBe0sXPq2u3VSbA3vT3g8RIq9DNU4iPNxRfkJ9wCAL3+nrbHDu0TA
Jvmc/8n6VaU+WgLwDu6TPiwzrazo0T9ina2m6/eMvBlY8d3Yh613dZDW1NJ91MtUzYwAtz9Y+zTK
LIdIivgvOPpyVog2dRz/xRCkO2NVxXeaKlgxY9Zvajco2V8finE5nUZzdHEtjOX8sAZXzRCPihre
6Yb12MzLUhgIyR05I4i4Q8tBeH6TMRXOZQHl4U/tdM2I0Pq+SklC6pUwDFOce9gXnTBWdxi8VG6i
fwK3zNnfaKrhF5u2f3IZmTRvJQH4KGY23ttItOcj9A7iKZKw+bsoWcKo46zeUm+0KhMbQZ/vB41s
TImy6JIQl+iDx9dlbgGWcopwima2ZSqky1EAJByB1uaB46ItUJ8ViAwY942D8AmgwhBbAkVWQo5f
LLSpc9jQf86aToNkP7X614AYF5Ylj9rNmk+xsWtAy8uP9EdEao1HOgggE/GbZIUOHZMiA4xEymCj
SxQiK2fjnYQUEj6OIVGoJ5lrrYbJpeLpXgk+pbKKIZfA3TKHRGmBHIl98yO1TSzbX8h5tiTg1xU0
qlRxqg82lqXvLi6rcHr41IyHz2beGWZQHyoZe1gdK1Cf1u9+VbsKOip/oYEtNVySW0WbA7rp94Q2
0EPZFsPsHuwpBMNIPgoFx+vXhSfFi6HWUaW7nUMHHH+BGgCh9yDctCd21Tag7mA5jpzVWWA4dHpD
jrUhK1kQZO+oCjEgKDp/9KW0OQ2rfjo/qtbhWmg9ggnOrdzSpojK3h9X4OOd8UP9VUyMNa3GYEjz
0pL4XpcYWtuP2bHLHtRB5EyhhizrqayCgxeZsbSfv7dVrlXAy+/R+9GlMHqlKdMG1v9/a6d6DGxf
3ypkOaLEor1RrGIdIMhOJPmI6QG65cffwlipxTTnVmXa9KiICrL3Hr7npow8ekP60367vnKAqNoZ
JzhmBkAQfALtdFYkkJqdCgrf7eHB9otQPYbiK/FDBTjfalXaUwbeS4uIcM97+7h7SJiRAHgY+Gap
Ep3gphNMpOTXvRkN1759+g4XjB20XaaymdtYXvuGlZiZ0QlXN1sW8m8jQnxFodScOg==
`protect end_protected
