-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
stxbvAVAr7H7P1mrflbkUGG3vNq+HnOxaeIzINw73YVYFafDeLB/u7lePCZm83b6VlvxMbUSQt7l
RLSs7Ly5mIFXPp5wbhfHiGXdTSjtnCMEyZLv+wySquHsM7o51OCZo0MlKRPVW8nefrGgj/asMG1M
wflZtmH2l/C+Pbz8emeFi1PRBQITEkV2KFNMAnnf+t2dp10RxQkqcVllkiQbB66oxissaguQjgGZ
8T1BBqrqZqo0KLI6CwFkwtzpw6CfTW8/h2w8GOvYTmaUNPE2VBHY9fEVPG/I8S2Uwj0TH37AcuIC
QdJVmJ17Py00ETm3u5MjClaK5F+H/z4dQJ6/fQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3040)
`protect data_block
B6CVmmby0WTu2azHEmPFV4YzkGjvAyE+uuSzEtpbH+jb0Yvwz+tdaBonTv+cSPEGo4dDKabtcUtS
DcNxwEn75OkXFn1+frBJABELOk2N2Kc3O2eYhTpD/ubtV4S9ITqCaD5QH0eaYujDorDH6Pr/z/SA
3v8a2cYORMuP7/Y7V9aHip7h64Z4ep6fl0xe+PtZHhBvXuoDwVdtaOMKvdY+l6ZY9nd0pm6JhbgF
P8ue76LLWftgjNHp7oIfKT8jCANGC0zP159zWebBFS5ZEjOGWNFViWJ/3Te4veqGTiERSjbMZcKq
hYCyq/qBWgAoPCkgatd3EUjKcb/RqfwX5/A6k4PlC2tsoLuUIIpOibJuh1ycVEcB4qhm/S2fN7ca
Il8/hv8YDeU6ZqJB4yJLlzC5kOjBw4PffUlmO1EFzTLs65j/i7pSWqnQD4HjKziagnablGOZsUbQ
NIfk6gG7rginGv63/scM96xFG4EdjDqhDiyck5dfWhtgZMrX/2e450snEDDc7EhUevbxQI1sPz3A
rfpFwzMvQmqeDPsfReKT+ZvEXyhTiHNpS0OfMUg9E0mZ2EPyQCyNgavDEWnnyOnOoht9d7h7EKpY
mE0YsBoqY0fezNgkTxV/63s53NxHugxZtgwrvVAoXjqrSjuzIMA9qomJtCuT72hRFxwiVmA7sIQH
QO8epcsW0h0QvRnhPoq4zJ/0smDk7g3aMiHAdTjpoOEeSmMAeOLOrnqj3OuofHDtHlpIJJnEA0eT
xhzoYmnduDv7VeiGAtcmenbEJfGqoWIS9EDu8LalROeoaCXo9Nyq+CIkOyONx+ycHJ/NFZBRWBLN
6zt4dz9gvg70DzZQeE9DnRtNdOAPMircQSG9X2iAFAo2v5w70NpalxQN/wgLCofy8bvZq5HqmFEn
N3BpMAFCV3fDTsQp1t3cdp9gJM8SrsCPM2dwwm17XxNBpMTY3HppIRabbTozgGD3drxMzLMqNeq/
npWYf32aRa1hTPVrSIYF9VuA2e2Scr+SzZesbkrjip97b8yLN3+MTYeHFy/EOFsD8mYcdCTdWs9T
dZ7bj+VyMFb39WzovngouPa48C6ANFGDYuoXFLswUAthnrzHT3HCj5PXZbX1TqRtICs4x3IABhYS
bZFA4OmsoUU36PoAUkrOaRbYfrAYY8mME8isUB3ZsO52L+JzYpEwMEGj8s7BG3+3XhY5HcEbNle+
7qIRlb/KT1vzMqQUe2LpWFZlU7b3pHHOeFH3jzGWLjS/Fs/OtDEcbYxxdrs2O6UW709k1rW40S6r
JgeqXr1y+MJqk0WxW4nXHoHGO2aFf23ClmHMo6Bqt+u8ic1ikxoIFlqxWle0thEQFCOqYX722VOC
0upiee61Dw5s0DlfX90U6C+LH1iqeRHALNaDYqUUkUTASgRU8zmtLeTxGqmmvscy0R0H8/FO0OPM
20D6bnJY07sNmH5Qs6ACvBpNTYyRyrefGPeOAHccp9TueWI6RwDVUIiO3y0ZhOjzlLZknOHIdrYe
m2O4vHaTs894QG7CamsjjpuekObAZlFhymZSfwKhjBCufHugY0QQqysqE3bSXxjTNGucH8+H/vd1
b35oaPLnXbbNeI+i3/9BSmAD6ZDqbjz0u2kR3rA4ezgeYtiBJeDB/jbi9ib9PoS0pR66Fy+9z1ej
Ff+ckjuj3oD6FX9HNC9XkJKIAPtaBYNx2QymaRUYz+Zc6Hyi74oK8bQzU9Boe4mWodQd124pHNIV
CD1qdMzeFzqWTK8FQUhMsVF98jUUGuRPJ0Pt3cGYL/1Y9xQDePWRQDqzBblw4UfBufvVSwd2Z/dS
eWY5d7Q82X1X+mNVox3xNQU4CnGL6429AuEo/gzUGPoJQQ7ReErsduC5uS5BXx8B7F9GMqxXk8eq
QUcz0w1uXkFJPWukTYkPacMkZjDoULgvy8tiSzl/iFmuM//bQckemthCnqgy+2kVQ0Svdn2WzkKG
fBuTR5jcGSAoI8d9ZHYe3mylYe46QL6zCdtUOE002jPO/mVcK/8g0gx+1tGipUNO0wY7jbrG9UFu
DwQQpHYDqhhmFEBuRNlZQSrvO0lyIz+SdCeOZIfPSXZf7Ohei1lFjIM0+6mjq2KYLSJZtFRVepU4
6L7sowoou9f/5E4B1rzPJ9O18josf9sO57+RiPvjFZPF3Qz5YIG5A4Qzldh1/jLaqBtZNp6b11oc
dW0SDT0/tEbqWgVrozZbNmYHZTYygySfm3Q7k39l8yH5rNhwy1zcxhKlaqcpnPEIudkTfuylRFGI
QHfQmPtTrO/MZt/J6XYJM6Lh9FfO2g+wHwDMhfPajMRF2xA2T/XCeXQuox3vDBnt4S1rO7nycVhD
jwPh3A/JjqYVcQDGIOYhZnn6PgepbqJoyfZO6m8/dUVXRSp7jbvZkZfbZ5sROu2Kl4xpZ/5Aq3xf
MriWJDWpitCFPfq2Uf+2tAs1qjSYNuBeIYYhD5Z2ZKSDayvFa2oFp9YOTRkj7nTJHYflGpwzWEHO
Erscvt4rATrK3meJk7vgFPey+4m41b1wXta2tOEa3m/1GU87jViI9NcNod5qS8SOK/lE891PlK0p
BK4Qmo9hqzPOCyhqzghi2G2RfFaPLEX37UBa0raIHGCiNttksnW374dgTcUvoBYR0CtTNIndEZcu
pG9MkB4/OeCjE5MD46WZdET93Pa9EtreKoMJZ31AMXGOrTNGgDCCmfO++cKC9XjkTRYqbcQZ/JCe
vNv0y5VK9ay0GYFMKB+KRsFyUx9PAk+WD+poeeG8D2ykD2HC4iPU5o7hN8vcSc7AQf/mdzrHLuMX
PIsBLL9Nfwd/NX39myqJsCkPZP5HEGLTHZqXSVM8oKiuWiHGfRBTXxDGEHlTKp5LWGLqOrcVDVk9
0Q//Jpt/DkqGsTVJm5r7nvfR1AMyRZ5aRCio8kg+rCkDQk+H9+2HHPG2Fi6VlWuaxd5lU7BvSHV2
alvrCebyH668L3Qpy0bIfX7Gxg1G+bVDnvhwYJugv4//PfZjYfDGvsNBAZctktoTyJLJB5WGHJfg
fDQHNI0B3NE7yrEEvD226ulSVFFR2L2bB/imoyagc2jvqksZQiFOD5ribtHL1IAbrdWNSdFnA5cV
YTTeLrpMGZnllKIAT8i+UivWvOMh4wir2hGV1xBqV/4C+ScxHyE5XD7gZRE8JDm6jpF3jNa1quia
j0Nhgsk6ueu3OPYUryC8Y4sS+TG8EOzYIm9MN9f0PLyqgr6iLzsX+dsn489tnmUI7i1kA8VmiKSA
M5VbFnCVki/sXwY0I4A8tdUj/plxHhSJ3c1XSrfZl4//NDWE3ZmfVOAc+XZ5040JY3yKruFLhlF4
h4rfkSKbB4wr1qE8p4m7t5f5vQ7Mv8M8Cace3dcL6fnLKCLIH3LPmFIsmLtsNR/VbKG8+ZkIzpNc
ZBEKFAFwApe6tf5MO+9z2Fpb4atgqsqSl9fkr5hqKyE7PB3BFwojC6ZBtQHn69aH2M/UMz3DvDE/
ucIOdPOZt68pRC1X+XOILR2iQAKEWEw+N/vvOqx5FmjyrJtfGHS1Zo37YZcSV2EXrtPV/8tsgJu8
Lxc2QTXIoMF4g9PsBSWBBMkXl0aukGrgVoZwHbhXUcnLTSG5xqcX3mbXKjteO53rXArJaBGnlYNo
eLfKz+XNsJOYVOrW38cytDeQOUksns9Jj+/LtQveaZ8dy9HkU6zbe3WYDeQ2XXpWIzQv55huyHY8
+W9qr83/hrEj9k5gti+4duYyt1Qw65UUc4At2a1R6Zk4aB6PefaCy4aNckQCS2WUwPXHm180YGex
ESTGRa4puPZQLzxVr41lxVlv8UmNMGgn3vLU139hZBf0XeiF9EiZ7m2qw+H/aDpIh1EgZklJ+InR
mWbb+0QNzNfLCr7pugwZqs9GY+x1068G/QLWV22x1d2JCIUicX7Yt/JgnVgUnkW+5hVI6WKwgamb
9C/v6o50eoOS2NSP0oY1FBRD6XWgOvKx4r8FnYjsMe8ytqeQ8CgO8zGVkTgRgMooiltCM6WXWKpy
yuU1FmeQAbLPzjrU75GjV2oKNg==
`protect end_protected
