-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
F52i+lR9Kp6aoKAdoZFIGQkuifdMRvs8yGZFY8frz8BZkh/oCXl0PMy8SvhYrI23M9Q2NIcSxZ31
29G/jvr1gOjHxl/uBO/dJOHauq/a3FW8cCeie3ZYLFmHBarqf0eZpYy7PYeNUkwx7ztdfwf78deS
11MSvIwuwECNjYn+A+4BdWgCrfjHZX0aogvuK8PIHxvh8G4Eq0vA82CGhxTnEMCSIj57F4v5FKk9
pnBqJGYkDViOAIbQKDr6E5xFQQUmBTWXzCInDpSNXTv/E2TtFcKDUNfHE7l7VWreEl75mphieHRz
axHj5nM/fMcBfeNZwakW/qTrOfTaiMABlu1CjQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
8hVIkad4aAIGmD/AODom3km4dtNNHkyWjtuFvFt0m/vxPJCw18X0PrAiUmLnIGa6nqGfVQ7aRg0G
WkDWtsC5QwxhGusZEQCGaQfhSyoyELiMZQs728OL2u/alnlZy7uY3WXDQ+cfrooZ76dpe+g4deke
/+fRt7gY1s2g631DDGyeBbB9DUdBkE1jza6L1PEg/BarFY4h8n2xMYCKutcSG4b2queqUGsmU8HS
oMcxUHLKr+4dUwMOTkN5F22m5nWTRcjchSRiDIDO5/9Q7PSfDs4ce+K5d0bwr0TpMpQGMz7LtDu5
9gvBGctXFdR0hUrrsvbpsHT8iKtmuNpIYXQGoJw8iBkkzr9Gs1vagktpyOAxPATDDWPLvbfaiz9/
3yrNXk34xe+9zHFUn5MZRMRKj50FfJHtDAyJV9hI53WOcVH6UYvgtXN0/u6i/G0P1MueiVe+ZgU7
pO+flJTQM9J1oUnqppBcS/s/wx1IkeoG1dufxjJFU6YVKkt8pXTOoilV86VOBFX4KUykzJNklLff
Mep+xiagzKpjRlPKGJjjPUuTRiLFagl+vC71CJsF93sjf5H6shdYajVrHRbgCbU9BowfkXaA6eAh
8hrFnwuIEONLCEaawFKko9sb/1K74eR43vsR/dvxQpnaev317JEkv5kAhaGdlcPw2idX/TJGWoGm
YKXgrZt/t91JXLadTzSprqi5qitcUhlAzriPrgowQwf7qbAb5K2hQkE+zLaSmru18u1a6c8wO6D1
2IsC3eRo/CBRaG3TFSjpz2usOpBbOVh0Z5IJVMDkyuFV6FgT1Zw9HI2TuOGyuHII1cEMLXNvVg/J
GGcHFdBNcHE6BamJfc4zv7YSIDvzgoe06/QSSf5lpZXWIHXabs8urbBvDQZjQTPjVSbrFexyESDW
lFIsCBRs6/Xbxwnc6Xgf6ZUJY7OFv5mid/jZRbT52YeWJYXOLq4qrRdcVyzyboIdSY2TD0LHGBkU
ozL/w5rWHsJfUFwbOVAsUyYDaE+bxO4xD9n5eLPHNgiz2WkFM2O9xUQ20vLENewxsnv5Ro/0N0mN
NMNTs6HIhxGfFEGI1zpoVzhJ/QRr8N1UyIbmkKCEuhy34ZJ348Uk4Y4vsO+VkLEW//Fnz9a69+cb
m9/RdRf4wgAYS2oiWE64ybyb98cFyyEKGAElzRz56TzHRoLPSQlQPvBHgldHre1cpsPe++37TTKK
6Z6PEqccAbaIPb0iZAAOasb3jkqTZkfPCR9VZ52uFigoYOkZIbXpeiRZLpQGkInEiiJcmF1FKh1X
2vH9v6jbeKiJ3PhwaQi5pX8n3AsROGqmfDax67uLTWSYdJv+LQbKgIzaHCmjS3HRI7cPiD+rL+N5
ttzmO9pXcGjUVKrswdqk2rI/EYucwYcGKwVnnOR5rwvb+aW5Rly1PAS/KGJD8SxxIL8JgHynuZsY
hEzjnHR4aea9FBXRmfRAVhMr8+NDw7sBHQj9F+r07r90iIDrLfPIWIRr7tndbY+PEANzpnBqZ5oU
8CrMzpnlk17lQ1O3d3m9kevYSPRhhlWsRWFDWrjaOz8EYmDwOiCghDZnck1yB5saQ5j9qfoUgfeO
aJU6xA7VCO5MWpgzpMN2C/MSLl5kpSKjwRXPvcwtPqbbujBRAH0vhZf90IRxji0Xkd8aHmHUZbzk
joJ/DTKECMVOaRSXC7gI+uCGQjTrRw3P6qI1lnPTUyImCLrgkRY/hisgTA8hLZOUFfloegmua1QD
8tR/otMIt+GjowFbwQRhGL1s21NqoppAtNM5rTNUkBTb48gpiK+PKYqtfo1Ea4H73AQ5DI1wb6F5
o8BHtcfbbwXFm/E3LNo4Dw9vBk+Q+1JTvja5wdhr6HQpeMk29lwWzvd5mP4930Ji1AMvQ3ts6fbF
ejo+WX901E7vwNV8cJ8c5WGkPFJ3R3y+BrqYDT+2Wj0SytAb4EOz1YlQAzhTdGIzA36e0qgEQsST
4xemTaxo0vTQheA9LS23NyJBUZ2ExzF9Ty7qP+GLojWoZuPkLc6rK9ckvi6075yCQcsX1jTgvNd7
xDhw2xuRZwadAFS1lbpjD9IYHrYvS9LASNKedlvBU7Q8uX5Xz9UWzvYs/pjUlNpBbGo25WU/1mK/
TFR/63EJIfD9b8SwxAxkZntHE3w2m4WJAkugPlBYpD3oDgndA9P9ZKEDfFoR8Jke9w0M4G/+uLVO
TL78xtCpU5oQb+/ZHRcMaJPUke9Qcpe3W5TMQEGMxN9jIwcMg1knvbTZh+/UdHSmTPlAXQNcmFa/
+j/pL2mzvM3wN7aG6dqWxUzIMNXKtDUS93NfyGyG096ObOtcPXMXWTWTcdzlfRNAyjFD7tppar/g
hEmPBCWD7n/B8oPMXTB7G5zfy7yiEflEwlb8YfoMoH1PlXt9stDSDL6C9RyxbteiteZcz2rKRSgf
AWnCzQbJz7ABvQi3j+4qfEmy6LGeCyKUql7V6AmmjBql0VduPS9P+VH3pmQ/SZOMMGGfwExFH0MU
GPXBSqYP0bg1ObL7exkP9hav78N4IVeb+69nugjmXIJ8rygI5LQC8QQapKCY/B20FTft6HxUE2QK
PaC7XYO1/T+5nLZq7ZfLU/5bFbR7V1E861ZW5kflGzTuKt78HqtxrSQqHQov2NMk9+lSKuYKWPmv
7uySZU9n5wz7ckET7LcypKJpuplBcAG+iPsAL4MPhwDQzWwdGpksH25QiMhqNSMLoE28wbq95Mhb
4iDDef1A0XUy/w74tTbqnPsLqzgYxNTmAZaQPabHpIHDjFFJj89gYbrffuOdUhvJnBRASeza10Dx
GXFGvE25cFFmuL06FK5dAhmFMwZ1qPx5dA46y2+XAhibhSm7TYGAecytSj2T4W9JA9EkWg6TPcMq
huom3+JvYmokBfYmHdJhcvDgcGRadpAF8D99kD2e3w4UCUhjkdfgqvYPRrIysJx1u9xMETvvqY61
kd8CFgi2vu+0/TU7OK96WcgxIkY6K1wY+urBgOlPxc90QfdvdTvDpC6QQHd87+lH9iEhtBg2dhJv
FdfD6fkdXgGKEl224x/PmX0EvskSI0WTx0pmpxGFyfoxEweW6i+YKg2xex/PjQbkHWIOk8whVICI
Y6NUPhfbhPjyySQwSo9cIQd5seTX57a/f6LMKdrnsPvlSfbBwssUKtJPv/hM9wHMmKrjqXr1RQfM
ymotdX2RdQts7KCyTR8OChiLjiLtN7DWSPZF8c4pl1aSsHPJLwL/xAqqpo+q1NOYYcSEUeZZ+P/b
T31kCki5kt1VafEtMbigSieljJgiOiiG2y/+5SQVoyB3/Kb1GylDah25jRjTHul4J8+A1gNy/JE9
fpucpBexd+l1gQlYqfo7yNXfkUq2Vz+kcZtjiyMKLvh9XjnXW2jEWffmlOuO5L1GJ03ihggRIxkb
KUBEfzuWP7ATPdOVVi9o9LsKNc5ol41h2h+Luv80gCvrxPGESxErOWdxCtZLHhpd+yypoFV1MjO7
IBxNSnC2ApgTHj8lvSf77Sa4Jf8BBvOInIdtHEy/ymWwnzsF2KLwxQYhD6/jY11SN24jb1NH+1HN
bLowk14o4hFmbKhzJmLxItRBU+nL0iGRYVhK0sstbkbji6YLvOOq5yEwgse6yq+JAoB79jsB144j
xj+4E2NAnW1IXgz+AVqQVSuIhFTP5lCp+/4K0vVWsjo0L8dTEK+6Q8JPi8kHX09JN9oyQqBEp7B4
i9EWrOhDJslIf25VCYwe3D57VsKnZt3bytfVLtE3knjJOopHZ3tK74Ovg7Tm7kWWIhLSTFmzxsHk
lt14RXq3fgFietDp4c6HRswzeZm/ytbaF7uirHGO0IfTyke/c1CSGBFNKp5kxrTcy7RlzXmoH7S8
HQrdF3E9spBtqpgcifa4fEPaVyiPPL0U2QqqCTTSwiab145+ESGQ5BTz9Y/bo4XDQTMSGWx/ecDE
7NGeBQZfN6z+HellCKQw6slFOPlSE3poTP3TZ2qlb+VT8zG2BBDV5830/nXaQqiB+WqYwoTR6EwC
hrBrf33MeE7qfUM+2I1PzG7/J8dfQAf4/Um0D+O5bXTdYJzDosCfufb7fi8xk7rok7IHgywZDlpI
ZzkvqLoVk1w7wwRxxq5zh4e25yyAEUxVvLqixvVV2EhF80FYcaqz9DM6U6LCDjXb8wPc4DurjtSC
tAK2R1Z6Cp7k7xAJqjnxvfLu1djW2mGQnc8ZI3ntzWU6jnPMLhZsH5h2CWkt4crceSOBOYTb4rI8
7RiUitUaJdb0pCkFlCSp+u/IWBQ2wM1DUGEIwqpUomQbLj1+Kty/XNlMzgkdOO0X46i7zCvq/hcr
1wyvXQxXPokCw0QeKd9tpnKW/CTrcuWW2AE0B3CJCHL70HpdEmHFfnIoENBo6GJdY/RyjDxeQ29b
NcYwmJMKvF6RK4kAt6aRPpU8wIcWoUAQgzbzHDEfJY410tkUsQjBZLEnKGbmn0hiyl+DQ1ysUi+i
Nuq5iH+oOEeHPTwYQOYfAdAM0W83tRof3ebXktKxqzAMZHByylzTuI1zpoRhfpMa8PoFhC0oCAdv
4PMowND0HU0F+TS+oOYSx8aqqmSV99AXGKkDdkM5bN8S6CVPRl3iKJPWqSHhYp6B9GZIkQS+1n1e
Sf6aGW86gPTupvdxUpc8MTGcp5LsGWCTaBuIO3vVYpMahFFOgaK/dEeYwm67rwPsnSABwTAl3hs/
v4FzShLHW/ySUEIOxqwLb3dbyq/QJLvyIwcvRzvkGB1ljJSCtAusEAKdWV3cPHptpfm28vFD9Cs3
34OtcwUfK7Z1e08DGXlsD7CkFah/Ljb6wsCl66UMw2cAMJMd/EEW5l4rWu6G5/NXRseit5w0Mv9U
faKv4oj3dJrUPtPdM8akZME3Z2Mi3XmWhAhWQgqISqlZEHju8jT8slxs3CPRZNO9vMYezFL8MZuf
+EXYIS5/54QX7mOIveETywao7jYeRQUETukjWR0fGQaZv6/OrmAeli15NdPV2xJiA68PB9Ofkc+S
lahr1dqQnlrmTQy1oNqdNZ6xbO+BIsgngON7bYuHIJ8l01wneBeA/lMwngJzDiocj1+yztd074r6
jqmEfHChrffH8BwJxwx2aDokU4hoGtNfRSpd9uyD4AVSaGwU7D6yjSbofx0bA+ZlPS1tH6YDGyvG
KliotosXWJPhqSvGRDgw6paF5DkdyqzeONrBfJIMHbxQ0HLeD9wlWn0tT+i7EraFZ7MsRvrF553B
Hwk7J72AgoMbyW1h5cRRO/4/K8/tCKqqwlwhAqG+YAR4l3kLXROnQsArKRYvROyyXJcfuENGIynN
RCbMFBfuPRgHOJrgdgIB8rFL34j/W0ij0+Q4M6fkqV3ILzqSpcCZAsj+0yGc4WKJY7Euzl4CDx+z
aVxzr7Ac8nAnrvxpqa/Mpr070pGu08PqmpKPhVKtdhm7osfEwbJXaYZtEG8WbjMcqzss0lL78TZd
qQT6VmN7QAoHI4jFMEYq9xaGYep7Vh8Tgkrcl7+++YS19R/rNWL3CFrvtuhy9sn4HZkqbdD01kGY
zX3hQSFvZ7mmoBgiJZiAeEF81o9wUCjgaO3NskwKd1jdMAN/FNwMKxUh03DHflZdE92vu/yvO8c5
zRH5Uuzb+IxziwxE5rgrse3wjq83NAWcqqHEkiqc4ls8k0RltXwhRF4dHPTk0Q6CFRsFWzzfwEel
0EDjcGmWTK1fJeSbqIWg9VcAZ2Gc79NaZwNo+iywe0RxfpE5s1hDzBg4H2k27kWU+xOjO7efglWk
eVknb7+bsSNXQFI9lghiZ2iNTyGZlxSJZxfrApA2KF8MWUh6m6V99Mo+DO5hR/C0KHVFDkJ8GMtp
jZx2Q1o7Xf1i5IijVi4vhKNPLwAJTHrhdTjz6afn6A6OxNxo854d6ojWpLOaSdL3OLoIfGlSYu1a
31yZggHeVseGxf/2LqtOQC8UPm/ftF5kZq+ncZYrSimrm9sh4GdIWeI66pPkKd76OWZMA7kzNTVq
ZMPKZMAU3wiQGLzunOtB6GERVHTmF3reSWPIUxpNz1Esx3ktBHcpetEWAnAsif1J+9bOCk3/n2jL
U7fxxLrA8mVRlZSXDlFu1ZStGudEwlD03AhyLhGdiUfAHSpNSQkEjXvs4kXBOS3Zhwr5fFpFhil5
EgEZyrPxkWvpn9UmNxwuEbMkF7yBdnQ5a20feZIY5TxeHFeAbXyg1/Ar5PL67TzkSrN0c3IteRrL
nAi98dSFZpQCefn0kEoGglAmVqyIw6WwG0Svcrc1mLBkJoo+7dF0VTrbPxCjA5qLAJ0EYASoNchZ
BycRVoAT8dmhQGvybdZvrL63VHuy8xew1swzz2kH9IEsj1mp2UnHcM6ML9k8EqrrIgfOFTZ9xxaX
SUayYE9zRsVE8scNBUvGtScV1moL1M6nKnNYUlCukCrfR2X/Q2X3QNgJl3CNTd4Y34ASzIb2QdFA
tePu2qwbEuJgSB1ER5Yy9MyDO255aeItsojFrDBLQVMhcKUcvGdU0QQHIOFe9XYnVJr9krzx4vRu
m7SJwGraXmt75FtbHnF/dRB2ICKjAqrNIYvreDGXShx3Ba7Fi5D/70TIHRvqokJJmznCUnA5LL7I
FWj2z4Y/9pFKosO+OCMhW/FRLbeXN3W+fD3BnK0kLPnxmn2LseBjGmvPSAoYHuQjC0i2surIFfBH
pl8aXaDVmlaYG+PZik9J6ZnJHLDiCecTRN1Z2O3F6FvxwjfODj3e8KvIYE8cbF6RcOsziC3mku9V
zJT6wHIg/nLSXnOYkJP0iPMzd/YsCElkuRYMAP6sBAN05Dp+u7PcCWUFlSYnE8pvv8+k2xKI63dC
TWG1r7RhfMSbxA/pmsjiFegZBetudV6vARTqg1RFyIG7swdGXtUUGFRATx2IjOhPQtsC5kLYHPAh
LXZIMA+s9Sp0XN8GmBlJ0wyfMdQAujPg+rHBaFzLRT8RBhjJs2BjWgKeuMoJ+bqP9fGghDFbyKaS
MwtElBHfF6p3fAcERWOMGRspI4GcIJZLmbq9vgNgslhBELt13H/LKNDtmLnVE30sDP/nF9QDaW/8
CzV/v5hN1Bt01YS46FwqyF7DmHhvkunC7xV6javCNGoOWNjwOocl2xAxsr7qOgPNv9rufZHp2knX
PvOES7KOnoLKQyi0VEa3hRL5F6dX7wlZqr+3aHQRtAIZ4E+5MrwHM07L5WjU7eiVX6QX3OwtI8zd
wY8VVdw2qeGNIiniZ6pJXo5ZgoNSnTSgSKa3sX8hXFNFqpqu3rQNBVUi3Lc712+eR+LB+jJFopN6
h7F10XvXZpI4ksyCBGelvcQ0u4ab2x/Q4ovV4MGD2ShjjgO7TcXasMVTFrZPYpWFgQGLjtshawZc
hDjK3/Kn/1tfdRU8yWHh9A4txWYMaaxHhn7/tPZc3ge+f4mzcqH8XGKxfRYQeW1pmRE58PjPuxeh
PO3ckKO2Lbiy2iepqT7b4KSyEtOBCulJbXBRrrWVNZeSIZ+vuwJ/bgHYV3iIuaYOX5/bRY9O2yTb
OS3HgjOtH1bHmXm/RRRY2ILNhEiMsVcyCrVRRtJBu0wju84CQuDLTQNeF+uZJuRYn0qKVwD0HMrx
hvm+64Qwvvh79QU+lzuaJkIDEzzo+19+DYYXd0oxQLR77Dq9mUGkBEWvoxhs1/Qkk1EYR+2LR+Rm
H8cK4LLC5g32Lg5qmjLxapDVsicrB0rMub3y1E9+WcluGGqbMwb997XdmMxMdp5ZUjbTPVO8L4tS
2FCKQPuT71GYSarVm7QxvGO2UHK/LZ8TBzFSpoxeucL/5RcZ54/CKnH8dPkyrY9rrmADByIZ+KDH
Q5QpR6QlAm2H6j0aHX7HQqX76i+7Ywrgn+J4Kwx8RVEOUDo2fcUY+I/NVEa6QJlPbTFse3rYYjiN
C9R9i/GhoqHcENo1M064zWGli2r3+nDfhItvFWYcSKb5sfSMw31zFai1C2zcEzWKFHn56/Y0lUmy
6unzHcB2JoNNaYEyZ++5IOzvKxCX6ex/nhvWLRIny2mki60yh0KxbfAttZ2fYkJaBdiLIONr5gMg
rfshVymQgyzkrHE2NKSO6NjT6xo9rWz8STZJlr2slRUTN4u73smHmOc6BnWdhZHpEIS0+geKD0Yn
QPvF+SXjOnoMg6l+s8pPnPsMCEv3VpAqSiqEiT1wrwYzhQaPSuUnQaAxrrhOBIh/raZLw1Ft6VIe
KaTolQifa2e1gVHdR1dDIHdGxX9DG5R2wHwjXgwOAMxjAyjaIp5T4noE1EvanZq4+bineTOckRei
JGC7rdGEbDYkkepZVCwWHV1lIO3dh0I2SIP4YbBRMQgau6vU8zStvAmpO8ds3zkA1Hv1CsoxYnE2
w1iaAJWOXSxCkVc41tXs6nbxm4B9/MWBKWlQn6fMt4oJ5WLngARkWisDmP6tp9WMy/WwaRyL+nGk
nMm+JIEEMdjzG3dtVDgU+kCGFeTXK1v/K6EN+patetU2kdOeSzSylIU4IP+6pulLBu1XCwYpBtNC
VN1JaEIZCfE4mFCRcaIrZ9Z+sIlRLhhILQrm/YoH/rviM7MiZ5kGZnJ3hbTnW6jsJzCsq4+zou1B
2VjBivq9GyJKdbM/mkXPaDOHe037tYdRoIV1DBf1Jh3U/rykX5KPm4+DWU8LbduivmvNB5PhIRAW
q7h78OWg55s/A+iwDQg=
`protect end_protected
