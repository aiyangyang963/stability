-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IaFLpEXF4X+MN83upuI8OLVm3Q4SBwjvoWKhehubEw7+JD3dExI5qjmhEWJHNAGvXSraUnjrUDm4
NeeiK043JXYIUAogcgRmJQirZmnPikuOcsw9r0/5awgrtRgFdZlV1i8oAOexsojjChRtQ+glzoaa
b3M0TvOsPh2NR2hRc+JjIS03191viYUyb8reJ5JF5CGSXBrybg5O4h/nrkRip6bbBznUIxZkhbaG
LAmX1rNy+aBKDwoY/4ixCnyJ1yJ9QgnWi8YuHcF9hJvLi4pIpYtt49hFCbiroFLigpyRRsowptRn
AhqXVKvK518DCBl90lvCSLJ7fEajbS1trBZEOQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
FL1I5fE5js2JjOeDDGQCjcBwHbqB8gx0LyX9A6qVso9HmzhorX2HNCq7dWXROz+GlyYnnEhLpkt1
G3b53GT4DwTiWbHYrbCXIozpJqDp2rbL8u5r5p0VuDSqjFMeJePB1jZYfi0oiE7uXoFeZ8P/qvXl
bIt69V24hagdCYxKh61AtmfDGwybPc6VDag+goGA3GzU2K5wpWaWXD5LGghXeyN9tCzPB531A8Uv
CEEkOcyyIkjF7QgeIQbDRftPcNXfOURQcQCefMh0MK6iQfeUoqoRk8cw4dMr0uIKba1S7wpsoQ5e
eYXoxwEqGmgOu7jV1Ol+kkCvmIqn3mfiM1w8ivWt9RwMLSst1N/BH6xerzAoXg62mjnTy+TBYrSw
4OREaVA409HBFFPRHBftxMep+0/ZyqXC0Ak80YDZZBjhB/NdCaAYr/0JpCzzz2AdXTl6Em/Nn6GE
evfl1acASFFNfIeBMCgvgyI2dOrGuX1NSrjqxDWPZafymKjbyx4dJXoRhbNaNZ93MQCH4VbNLIKn
seBv01Q2anqfwxUfEYXxIe+fWtkZ+vdIImXW3MDOcSACtDs87HNIa/LzSdJr2X8qOFpZY+oF3sO/
9tRlHrtW+BqpcnNkVk4w7heGDRXoCEUQ5w6orFKx7qgNywFu3aMId98TAy4E53dzaRxitfAXAz6t
IQ9Z1q1clsK62NXeZu20bMJfqNqSFAyJZIRu1BHG4p/Bvv9Gpge1YJA/+nL7fIyrdqUNhsCSkWRp
fYj6hJjYtWroSRm9WC0ajxkpSkfJnlZAtCw9ydPbekB5ZBm+AXGymtfLFnEIIo8Z+HMfz6EesoQY
YWrZBZBNz/KbPU+gjWrdEsZu57Abr1u0QeZhHrbh7cQjheOUGHxqOjJBl/ibvWOr4y1gDrjBYPvV
+C2JSRqcmyg56kMrG+fApoc/Go0777vkAySXO0BhdbWwiqGsh2PdLSNiMvBoc7LOdd94Y2OV98rB
ibC0o2hNDlt6KQkSb0g2Q98siKnfhHc48aSoN5LAdB/jDOoNS5GFY8brA+EuWnjrdSsD6fZAy2Ex
LupohuZPMFT3CDQ6VXAttwIZpZw4nqolxhKGUsYcgvw9EdHnWM5azK4wIthl9I7472PToEY8GQIH
WE1OhIIuiagBMkq8O5K7jzLG4z+ARvjoPKygZkSYVOPQKLHEABYrLROYBzN155kKYcI7kAYUpEK4
yrYCEbdJ77C/XqqLIM2sTMbKY5jKkp5h8LuYhAgNPXIEQaFZNE/NekYkCSiS2py7PVbTesYsjbNU
fpx2T30fvAxBWasTKh1Zpt1V3H2UWDVsJrSEAv5KeuugZvXMCJvEukDwKpuLqUwu6IIcp6UMTCqQ
wG1qaHmprQo1hMq8hYNbeD5Xenls4GbcGfsfn4gIId4xqvosBHgLXQWsmuL9vTzumpL6ld5RZOqG
Rjse5PVhRENXXquFPZrE+l8vGeuQfNacN2CuYNEsCNPqGWNQ5x5o0oiAIX8xCcNQzcUbYKMA8Svr
Mi7ZXbI3KucBzzppmzsfW3SHjSRKqV5SQbQVzwG7ZwmyI0qaWEpzh0J2Uhyf1/JuMaEp+d5l7usf
8S3A8r+er/gtQD99tuqpaRjpTRV/bq1a5OSfUjzJA3Q9ALEtIqyAA2jNB6noh2Oge+9UxdU2L8TW
8R2bA/hDQ2lHuec/2jECW8UE4aOJ+24UFgXyI62cPRGS0yUWPEqAhQzwx+ckOSX0k8ExXE+GaG8X
sRMymeEztUAE7YMJg+pSgxl2KTxFKLQrWlA+Un7S4p5v0IEKCASK+kkOP7uMBCJx7gkFpZ7eLlvX
FDeVRFACBCWiJfDxXsLFkVYQvzpNY/AMT0Vrs3EA6fve79z2t5qhVG7JFxkIPdJvZPc7TyX/UmOp
ypSKnlEJKfGBhaYLhJNiAlwZT8j5hk3c72Y2sJqGoRRrEAEvL8/U1t5CYlwahgclhmqNtboecRGF
tsPkQeZoBNOp5wu2WA7KfrpHLkqgdveH1b83AEkaiHxeA+alWqmHgqXR6pH2wxLsW7dqjOyBN5xk
m7xj9Fc5VRPECSDxFZ7kufz4L4VTIgUI75ihtoe9SxtLqrwyVnMVxTwMA2iSI0wEtIan9UJKjSoj
ORDym0Ag98pZXeRHYVksHdMLjx3Mj9tMxh0MtSdWbu457dDr58LXodyVwaffeXVE+8gHfEu5p3la
lgcoz2QmsTmhz3AeLepokSrUCVZxYPwhAOnjdz+gHaI3B7bJMN4J+R+hWmk1NCWXq/Lui9VHaLRk
W6UuiEMcKXlF0LkzRNmU584xJfCXzOa46WYu1xfaBc7QWthuiTLNgzh6hYc6Dk1J7ajzZOPWcHAa
cp6jA60q7P+jXrs6j3kGuH2YYdji8H2+BGjtNQBDDpRX0DljXJG/1htyx4qilMjAm2eXOZUG9WsN
5OwkJ5YO6hAp2Yx1vTa3/7Gjm+POyhu3dFfvEj1xY6Ee/z3Toevdn+iyULzlPfEgZwRKyK1P2/pR
t64z3MHyINcQ5MmvBYg3DAioWxcW5174p+k7hELSb/emVgc1okLLR3sGwcAoz8gCPFKNPkTRbR9F
2Dq6KiG9hP1FySbSZ76/P25n6iZhTVScxGV6n5xqheUO1aUpxhqFM++H/YuaCcSuZYZqFQjBgG8+
3fJsPi3liZoQm/QOtHcroQPZZhh2kyME7ogjO67fvpXJ/AvVu4ezcR0QdNTLLD/z6UGNAEoqHUUj
FHnDEzd1q/tGxAuA9flinADPxz37KJ8J6rShQkirV2SNwpCqxmmCapJyuSa2BYF/yKHMGRgQF3NS
VOtpFs+KPSMCo0bgs3mHUjXMmCUsfQD0n+fCHR4rYQ2yfGnn+6LknS3PmM/FB6mrEgDIVwl4VqQU
GwQo998Y9C8tzEg38+kLxCecMW30vtzXkXv34COu3eTcCc0u/VaiKN8UmVJFCveKolHaZ7G4FJAu
TcauvxUClYHr6fKAYRFdWaIR1o8nFUcB06CzucpxiLE4FTH20plqRys0ziR9O7v+MA8Ipj98ubGP
Nik8LzW/A2mQ7/GpchmtRU3vv+BDKykjQA883zXGYHPhphpTj1qnGA248GuBrVEc9j0h/+FTgKEd
s+29hulOIFTv40+ATer8bRt/2+vrHkFsYBzC/KrkINedxWk9hHWkC66gWg6pFr03rYldSPRRrP35
i4lBVDlm6FsKRV9L4UDpjjFEndPR9VF6iC2cO83A2giqFDzQmtG5iJPssQ29Y915csJ0kEcbMY3I
jOTn1Pc/3oruc3/BvxyOscLe5AKHBuPdK1ITTlSB7OCP1AWbsD/bLymqsxvVjSf5G4eHqI71iiX4
Fzt/beWL1ac+F59G0whBEcHXEuh0vkRLtJOYSCgB4DgCSHoludprxZWevm3LZT5zyzPepMRej73B
FiTPqEy1Rz/z6p4X27LTt1vDheNn15A3G9gXohM7qKF4iyBy1h++eNZNdQ6CKcWvv3/s/+7FhdVe
Fj3funkp8zC82cPfjLzS3aXwApyUrlecH7/WpSlhOWvGcwLBIXsdDhXd5rM+fZxgwYh3pCi0TcK2
az0tETD8YrcZHAHTSFoSae2ZmZ/s3Qd0+yaptLSBtMZ1T3a/NvHA2X4BKo30/BrGiMWzIPIuHljK
Fj+8LEQZIdnmGcAHwolAiKMiWkkU8j8cmPbP+O5kOUlQ8K0gii9ZXrrWIJFpK0yp7KG6dhFGs4t5
3YBxY9YTyJuDXyyARYbpzflPZXp2TZj0QyWBfx7FD3K8a778GCQeWTAxDe+uZ3jkw6C3Bn4WBZEU
4pGTdTvTJi0hVgvHGzsLYFcyfevTAGWjmG8teAsd0JWqZTAmbGf+wFysf6KX5IaYqG9q3rdtBzZC
L5DUwppF5GCeE5TB24Ur7g1w5hk414tWl6q5WL7Fclp6wtKZbHcDMqekEXdI5ixHtGbPH1QLbQiG
wjLjigv2saEtd3ccwzOCd+on9pNsWvpTKLur18lVtyjkS3P03ARlYr1pxVpga1GFirEm3f9NJAqq
GB1D4UxiETl9m90m9lIIZJUPKcB2xnUkbbOPML8oZSp/EgxP0HZXdae3G4sV/OBLcbUeJZoMna4u
cWoc1pqBtZdCCwwNWtMOwz4TnayzkccZcPirHd4M8EktpULc82D8yW8wg2qIW8RzvL8827MXO2Ad
KAKQodF60saDqJBvsIJ7SrhLqy6WJSKJWO/UxOQYWt/plx9ei0caD+cQf9XCIOmcGDJmAtHaSSbA
Eq+aOhNRCTLzMKgegMxHbxwzC7qknncCW/404merZ/ZJd2QHvf0wXsosphT2qOWR8jO7NT6j8+jR
0phk5MKrCk0G+FfZ/rgYcpWKBRaaD/cp4P1jHTIzkD6C8eyFJ3BYCsgJZ6vx986jGO6rEl/i7Wzx
lidFoNik18T0Pqfp5HmbHD6z9oxw1BUvIP+536hVJn4EO9+ws5rXaQREbnqpnzaVlJlLcBmN6OCq
OYMMgmt9OFF42vNxv/RD4zSeIaDDSSKaX0I2HYQpp99Ig2gZ+ahGE+TYvrzIGcbvTnyROkISVje8
qikrM9TQO1gD1A84Wuy4/i88kvK2FuFIZJKpfdrPPgaGZ7sszOlQaIRtYopIeF8fS2RNRKIftHk7
kHOdDFVKplzt3kelkLbUJD6W07sjX8k+QX1fVJtveY6vYZe5v0O61lpzAKdLAghKEkfI9ORAazDY
CblIsYidDKWUu/X20IlnivWHXxoowtVnrntiNcjUleOGc/9z7ClYZFei7R81lDfc3upD7dGkawsw
GLcm9e1/clrmwJ8rjzC5dQfsyzPBiv/XPJeCyMFiMel1txtxBNHjfo5xuJT0eOgzqEDgh9CeMUeE
brzAbeYYDYc/wQ7EofF9drSrMIW28VFlvooT52w2GuT8DxY8BPWM+aKBAOzcDKWfHfXQ6DR+fK3I
LyjpTTplvnclchAbVawvulY2Ihykk2xxr9Ppuy8ida7KZA2E0gH2l5vcGxELsmgajRCwDp6XqYP+
61nYDuEtMFCyefHvYH1dfvKdbDtv4b3ZwqoRBtGAJUjayC4fDXxi/V62TTj/PDFv76YJPiiIIBfn
TbZXt5YLhusL9gB74++AlNedoyaXzEWi3oTBuAGmIJiT2Xyf+ogVEAKAgeWcNqFojXEXYfu7Y7uv
adW3gXh/EAZXBcV88ZQkb/atmGi8Iftx6you4ia1APhoEDIT3kVPm2VtthY9GK/cy+IEZLLoiaSX
ELzA7ydBlc8JbH3cRQyl/xZDoeZmRGLn+FcKHCKTcyqK776s9b7ZE5EQg8+Wv7at4QnEEZoznY6H
WkuaNEykJjH1klhHPhydfzAsQApthp58nNWpDpisNcEQeA6kn5AJr0b5qttImyT8BarQJA/Va1fO
PF4ZKABi7fBwz665fp8+FTEU9jRjFl9o9eNcknUAANPUZ3dbswR7Pwuj8ZFq5ghfSPMHh29ugjr3
RiPcIloVmWD1EupMks7r1+0rNbhpn+7fQRxr3N8CWauV9icoPRVaceM8VzVGQ72yfEKIdbBgeD2/
+v3ZdZGvGMZoZ2Ay7b0nYC6WxF8iR9tX3P1ABx9RTkyYwebbJEicTXudr+ekgCrdHjMS+JEH3wmz
eS3tOnJSo8iXS8Y66ldip1e5auJO5gqdTERygp2J6LgZLl/heQnvOF3+6f12vYvmTOzHxMyFk23g
Fj2fIxLcIjPEKrM6MNfCIqeU8LP0RGN2pVoluDQthsqpfHxf7K5U7a8cV69aG7JXX/Xv4t2ln5R6
LcIl1mz6FyqM1XIPCKGwEU45kDLsbU6IZ/pH2wduAJRqPfum0SLJCU+dTLamVM4uABGFR4dPDfCO
mRtoJh5VCllcI0trsq4Mm3OS47Athm0+sf5yumVnWfS0/z81G97sQwuXvULURjBOWogmt7L+nXdd
IDuniASvAzBvBuOHfEXzjB+N0sD2MatYGLHYsJjw0Td9wGQh1D+AE5WyC6+GlfCrjg0BxZL8BuVD
QoBwJXiNTRF9mz3OFLOvT1xZ/rj3Uu34aiglJySaBeR2HCC4mmVHpYjwUul4ngfF5K3nbKt9mu9s
cZmTdsA10Krgy2GG55jF3qPsV/2Cwbs+Omy1ZvMN0b1dim2wqvt0UnBw+7cdiLX/UMnaxwr3LYFl
1xJmYlfgCtSLBNOIInPe80rR2Qwq4hZz/lOEoQzpKwF2+E9lf4gD2zqKOG8+KkX9Q0SCtypZ0fwU
J2KvgeNg7Y8V2A6aVAY/quAedGKed0sVPxiLnTvKJsENcXKxgYtitH5UNTxpAF5kd1lZ0ckHK3OR
Deie6yO5FiN/ebYhduJWAmMSXmJqip0JkGgZWWUFppKVSgzR9jfnsYO+uAVJZ5/9VYblUfF8VE/a
HZq5zGIGX1qW7uva5D2HZpMptLFA0TvGHNJzliSncSP8Td+LEMFuGv/vlR7ZDPBm01k2bFWpqp38
P4rz6wp8BaQ8SJW+VTlD9ZpWWLI19pUDd6G/uLq3Ey7nsJeAl7ALuci7CD6TU/XTKD8vkO1oKSB9
wNHaeH5+90rEwsl3xleqZjSyr3nfJ5D3n9eBb4rG6Biuono9o370Abp28TwcOQSSm8KNPmy7/M8f
dWtRpKYEwLBDTzKoOrJEre0WdWZnPaynuNhBRiYCt8bGoumNB9Jei5aTdsIm9pRaDl00AAkM0at0
BopZwDNeMJy8m4AxIuJ4GBw3qYxGsFFd2uY+yyuL08WRLSO8Q0A4SbbrAhaZZUUClf1Ao2JPsVxP
LazGN4wYiu63Ykurce+8grbyvSymhPwUo3QAM3S55/uu7QEsMMN88AFoItyR20C6so0jI1oT3Lrh
tp2RwlQDHdhMTcOzsDFo5WpdXe9CwW3aqYcwxDePDoM6bsTOaSqOp0JoT2ou979PkVOmIWc11Tdn
7+xskiUkMVaskITfMTiKBLU9QFAgLqjBEKU8aEWYYFu8GaJthoJKc18FpWM6aw9hf9EPPeOQvtdi
KJrCzF5vdDJ8HmLPuryAP7PUHoR8slybbqEL9eHnqTlEqT0NAg+UI914v7W1pmWUNx/Kpoxtb/B8
cNDx9sK2m6BNJLyrq8mM/YK6XJeFu1N26LNx6Ig8OLHuulPTR4EduALZcR7vdZBdOC577mTUCNWl
3bYTu/MOpiIpHUJWg7wTS6l9SjwTd5iJOi86BM8hfbulkos4Cm3SnYKAmdp8KTvSDNCd+A+L2xGw
4CpWSXguVVsmbDUBgh5+de4EBVJBWdDg+XKF3nyjPZ1Z+oyMubohF0XBz+/y2NEskCzwiwj6j/nl
oxGK9gxvpKOFksQ6zGel99XWqCcTvzYOnugy/cyAP/Agvx0Lz6FRmxNpjobJLpQi2pleXQfDgD8L
colTCYBDvKs/exxQTOYKNWcZPE02Pi2z1wIJwANnFC8u2RdhiLw0q/040Pcdko9pF3woOu4WWb/5
hIxaHfnvTc8AL+EfQ9ajI8/sc6EOWV4A9Z18hiTzV6dMIR9TI+ODypFTKIz2tiJTnPo+MgaANaue
aoU9/nUzi6pUlGTyqT+rnSn9xVhmhUxyBabzlkkFl6xydX7ygwU3G+loAzv7mUjWK/hEiWMd6PAK
rNzNY6Piq/+JVGWCVK8Vgb5LxR1UXvami4khM/brqfYATNlhqT2Lz8NZvDB8az2Npkz05dcd+AO2
J2x51u4E4mM0ys1dIUAxG0bbyeMco1HGnFnT2WCwwWMjl80xcYUC34AzpcOahxU9CaHvh1kLzUCK
QvHjKKjxJgFKl/JEBgxb6Xrm1erDBPnaMj4li6AXh2+r9D9sMWx/imrx+cz7Ti5DS5/LwENI3hz6
LK/RoMlYlmx64k4nT8FdyihyrbFs5o0J52p3ZYBEToV+2ksVzGK0X1haT2CMzggbx12iV3ogaqoB
PkwpzWqP5Hv6RS9Ups+MKh3FSoLtEQWkMIsVzC6mroRGHBcMaDZQwXoQ+l65tLziyz8Z6y3kabGY
8UPLQ2T4AQo0xD6kJyG4y8NQYOyn1e6ETHWkZXCFe0/6MZntUg82z/nSa0+JtttTRuG+xHWYdR30
kHxksBfGPxA7MZv0Clm05vy6rdSYYk5qtdw95LvaW+LtsGdYj1XW0I6UnhO91wPK6sLQb9XEX/Yx
M1lB62Cl6iJSKjYbH+vwUw0xM+mb4dFeJPasWiWM2i4j69hVXPJcge9IRW2aM/4Rj7j9BUEulLdS
Fuw0ER4FRA/b65j4Op3CnIPs2KeJ1Ks7Q3PaFkeKMSOqYE3uUZlGI/CCbXtYmtilHRE1AjV8IT35
+VGMgGhXMwVMbu2tCo4MBZGxObfx9K0+hq5qBeE8Cnq/ii1nJNfZYQdu/4/iKNx1SAZfuUc4Y4+E
DeLdXbil+Wcoi7FnjnFwbCYKxLROuH6xPCRUHhKqkjNObALJlg5GJ6/qbwsoa/W1pMYVpFDfzuxZ
JiXpkfhU4D7QdRD4nf7vdLUXEoENecv2FwM+nQtjSS/ORuQp7cGzefFCjnEhWCprcD7sFmG0LZoQ
y1Q7xQ1EiqsGnQeNcBtyDSfCRNlozvYCAm4TbA7YpZqAhmVq7e9szGZ5tVLj+ShF/XwJWPXwGslb
WdFanAPYvAIFTHq1GOBHUENA6jxs0rXI89QJYyLpf+yy+dZ/8Pl8FyMrfvmlsmCeYAz+FHUXeHIr
9k3zCchsVGOfgTdyVZEgxf4Z+PfJSaEPCkLntCJpfMhQC5FvumXfrzSjKJ957Jzy306DJvjnVt7x
gIGKWw8FYbAN9G15jIMbY6LkcO4vlUptSUgM1DY+7UoCKJmzWhItoNYW7x7a4VsaQnOGqvopI9Nl
BuVgKtKL17njhXOJevOhbH/CuwwkGuXIMuCmAVYpap7zPw2Ff9t3tjOc/tUUzyr9vzIvkc73f4wM
lJfXzqtJoSsvII9U7etb5WTmD4X3oTNpHwBBbPtgXQXDbtevlpKzNrEnuomIbLnvkcw5xjo9n7f2
1e6dDB4oSHVe30RSLkJzE25Le86466pqXEGXQvpLyMJeLbqmAex1/2QF0ctLNyFO3mBiVqrT9S+V
Aa0zeW/WT5GP+lKj5Wh8LRJ0jrdmpEQxWrhY3NdsAGQLIvHujHIMvY9sW+795zVv0qOBTF6Y0OBR
jsEFt94ceVAytzJfmwswQKfAfCI/VORRQ+NbaGsPhW5IwlzTemYg2eScpGvue0ACZ+PXekem9Q+J
gzez+m/287Cxcn5DMKOFz/IIDg5beTc5wzH/OdeQb7gsTP5mvgWdtDiyooTFN9ztpIRO4lmyxdcj
EhVcpNZHUUVPvTp8Mkn4uf0MqlgzdXE61HABdaD6AaZUFSLMDaDX+CjgzTwVkuUBL0fGkIMQsNSU
SrIcTZL/XWx4IUMSTAyydwTODw/50zWsTcSdHe5+LwstKDV2P7lX0sQOhqGMI+KukVek5WhOfEfl
BTl3tFLFvJ5vReLznJLVL1Mt8j0AZRAvzbND6JkkfY/BluGVuDd8gCgvfOp4i5rxrnQ/UyP7oLE+
KuncgxGdMTLr4TLiXkP8GbH3acVjFO6mwBrvD1iWlk8mjaDrWCpIh3On/B03mDYAIhNxDLqyrtsR
EGHHmRV6I/5+nQ1E2enTTcf7i0xVjcK43PRrsmCKOyF3DvA1ldlxEa8BqsSlpG0UoF7jZ7DZtoHT
FEgrIzH8kuXUvCOFqBKa/SDDZFjGZfsoYWKNFeRxVPrLwt1rYGUlPNY3ZCI+ohbeNLvjRMfA2zva
ziVX6gBdXlOpUGIwETYOPHabICZBDSP2+XBWlqfva1zpbHtpzMu7qAHmh3tGaDdyP8bxvNAeKYBq
qySQ05Hs5fTBhn/Cz4PpcV8xD9S/PLlblhPRJur5N5ZIrIyOtQ3Q+7hOjZcWIXgv4c3tkQWpMfYz
FDCl/urq3sV3EfgqLHNUIb8yqYQsH0LSd9b+5hjub5gjdm0fYmnIh4n8rsePsU7Q4eAjkEqje/Pr
ORW9O8OWV3dMLEWbJAfDzqWZCmB5ApTcDxxj0H84BpREoiGNnKH3AulsQEimK8pzyaUQYTo8iB2L
9bwYzoHnV1g/kzdRFfMH8wICZw8wSmOYhQ62lczEXJtUfZmHGQjH82iCozNxr8lIE3elGpBdWKMQ
8S/TnrjZRStxqfMzL+N0EOW3/yrVmpdekDRkZSHriwUl39MypR/Ayap1qkjUBrdsyeLV672/0cw7
k+4IoYc72vkBd3A9+ZKf/E8deFLncoCukL+008Z0szsq5pDFRq5kVSo0sEgRxWUK5pUT2gfaWsxS
kiQ0qgQgRo6BE5qBxcTbAeZMO/YGzX3x6CNZHWQD3dbcsO9fHQSTR9B4cNZ4X+vOKl8H0Tc76IOp
cooMWxAsAZzvE0mZcWLctQ5I0pR+ndJ3AJbZ/NbzX1eK6N82VcidjjeDkYMUJJWEIOpvorqCPjUH
2RYsPDGCAIwSLwYEXESHT+/F3wLY5pPKL0TZAmFlhUVkPeowzK+R4udA0n1Qy7Lm9IMXZenWzZV+
E+qbAFDFJtSEpyFAouf3rdRkQHNYE6Ywg0CusiEXdmVXipJW5qBbm+qfwCYqfCouMvELldO5P/mb
Cj79MKaYXhw4Sm32C1Oe4ImCKjnsRjEig/BHswnxclUlZ5NS0yrID3E7v6po3AS2F0o0ZimxQHyt
X7CTeVYagHpNSSBQXReH1DA0kO9OWHGpXf77KP2FSuQZ0R7ChVyH7LlUym6eM1yeOg5hT+zyEg1d
0OueU/AVBE3AnkmHD+/QE0PDSPk6e0cbqCPL6+nZoWk3L0k/fWZh8xIM7Hq5NZrKrbBx2G0ZBFtf
+NR76gwV1f+6A719HoJH+IkIom2DVSgOWIwFDh6Mzqf/pKaYuiXomlMukHFclBTseJhBZNu3PB9e
VXFay4BmZqd2veSKoYMiwgFsVrb55lF0N7TSozV7iSnC9TlFFPwlhGisyX7ITuWwSmD1Mi+vqy2Z
YbhV9QPYAg9lSjucnJZKyP60UCYqstkIAWRI4/oAXqdoBVuQ/jDQs3McE9/CXpo/BmLtAma/OBWN
nuYZyYOcrd1eQn/3KXc0WxlW0JPEMdhoDHQE055Kh6Ccl2WvQPsKcz7LW88TDe86Lw8ZcQydDRFF
plrh6nQmQUP86Lh0Gszy2lMlUMzNBHSsPDHimC8ZMKod5uU6NiAIW8Iqc1whz5/l0PJ21HiXi4Lb
xEmYTnjO7BW7HItNRwH4rLMkT80dpR9VEqXGOZE2fgi0W38C0kPZzAwW6jNbNTF287rg3l4AGnQF
o6YpHCIfr3j6/3N5xjavuOcaFTOEkLDp02YmwSXWEQdt3l2u7epXNpnou0DIj9/2DpkXEto06DdF
GAzVQvGIbgDKBuy1H1UrhSvmPubKzlSPah2v5a7sEBXhuyqRIE8f2UWS3oXtjsoEbADUp+mtRafA
OJNgbnKZr9a7RNBmGu8C5GDIfZIP8iAul33aXA7qc5XaJci73AF0pQ6NwS8P9ryuxpdjz+ciBgib
PPtSGNmKluugqdeCcMId52SNja4+CWRARHIj3r/NOOal4Uo730yy1Z7ohTeUv9jY8KCiDN13tqUS
tXEWMJO76wUFOUlwXXExM48HUReSosIiaf3EiEz3JO0EiWnRndhtlg/gAlatSzkEGWLGyla1Yjr7
wuglexyyhJsGJpK+WFPxQNlBYXLv/wiKWN6AxMmH3F9OXqD1SqxnCV9bX5jaKNfBizuMjYBM/m2G
aTx2/TN2BT9ErHSaxFjnV48/hKy3AYwQZJst8KuKf3Q98uWVxX0U3gGC+sTyZN6GdGElQyHRVKcD
Q0OyLGQVk6Rbkd94SwdaCLoP7wTbDylHhWHRqCkVkEBBc/aTKhuU6EughPmC
`protect end_protected
