-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vlOydmzJgHsIIhqO2SjmKEDhZTmrCSSDLnHdcdaSIq2JdvS+7mZUaddhtwX8iqiRjtV07CS1kMvL
0F5D5kpXzfKu9iGFR5e0F3AJqNythVDP7UybrKHSOhvYv38x2D8mKHA8sUXlnOgFWj/NARp5NWcq
wjR1DX+nJOfxkGdBaprrnRyAoXQ7Qc2DAUTCXHxSdmbrGyTwZTpaO1c80p93f8+hR19M6vyt2QbE
x2T9Q2LCqJPtNMSo7Tl592SHBmpXdrHXG4xAlAKHWdx3dSU/l+gkLyQa06iSMAKgI2gPVS0FyOt7
PAkVhfn7q32sPC+FcqC+y2df4hHhkRbtfPUk2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
8fvC8QsRG6UGeu13vZQlvtJZFxnCWlxYKC220n+DNWXDchBHlDJE/b5LJlyuKAjgJz2Wj0jzWg/V
ccy3TDaAIkZ8eFFLjinUpmM9/Hyn3/0BuZTq/4sM7MvggrviTYB3k/+2vc4glmyrLC2O114ZcPMh
r+vS/rwp3XxLPkHHqsFjCRQYgA2pLGgTpzfipnkE+YN0QpEva4iLnkMekPEWY3hr+Q4bCWgwznyn
Y20fvzJhgv7elxmNsc50OtmPgx5B3sPuw1nEPUcCL17XGPoW4WQHdNCSf826R5ec1FdLgtpC2NSp
HU9frCZW+gjKJtzQebrQoAKEzaRX4GUIcWX2Q9p/DX9da75teXwWxWugHR2H6R5wx4PnlVg49QdP
rWQ2aebvVkx5OhsPHr3XtTvVjzfUHW9mcToVLS5+pVv61ffkXPFfNwmbfqRrfuxx782Nh8oe/peV
QVDfereq7z7JoSuxCFuh4j5zrkNnQxSvh1dInwKbLtGbOf9qfgMXUbazW1wBOty1Aa2g9GwFEpA3
cnFE3QZKamPG6IXfBThPUB563rh0SmU3+oaWVL7tctZ9FAwv0X6E7mGewugiTa0oXl+N1U4OKSCY
DtPzHHDGJcgKH+7Y7bO+XN4O1AAdKiZ/ElJSaaQ965a4DZTVpb51GsPWCSVSA153o6qZMW+iznn6
JWI4+MhLzCCGP163amaqf0j0XvlXJydYY4K2fBxQObJJOnEV7bPjMY+LWwiRBexGsfptjqbC4ePq
xtW9YsELXAqWIy2KEMpPDIKM/we0cnbjUaQrdZEoEQrE7Mt3bUkVjADi2uQkgRpfGjIww3q90mkJ
DZV0pCc70xaveiD2IfFT/r6Ieb9Rqm8o9scqsryEYO7SpO6maKhacdTIklXaC1I8eaBdQ8nEW9ap
bbRJ3+JfDrVbJSQH4nyJ3xChQvittoyX0TP52nd0p90Ohmer9NBNsyLuTEVd83BVJdKC++rUvD32
mr1xSbh2fQQb+eKGx3UmzTbM3agdB8sPynplR2+YhpaR9fd2O0Dkvc6ndtPp1HKwSxuP7HPevPyr
DjWYSxZS/Uw4DCgvu9dnQCLruWGD/UmyaB5a38Uf/mxfteUTE63BgSBr9al9Bj94d74WVdWU3/95
4i19mc5Ze63Lj38v0tnQHgqDV8+MJ+vL7jXdLVHqNVy3IIyQ35aa59n44iBsDHdV+Bzj5Mp1Jd/q
ZMjEF7WEF5RcuKN0auKp6byHpRZx8LjGn6EZehZbdfD/b5VtZYsyruNi5qP87gFG2+bmUmghFheX
pwXNe15RJ7+2R3njbNf53iIImLwbJIeoSczNBlpQFbqhqIubzGSR5zV4IRu9scfkhBUDkIzIqIAw
w5SCd+0j+hjBhlI9eqggQHExFyzHGfOxW2s/elG3SNne179u8nSZyjv3kCU/Em/xqnXNP/k3aUMW
freI9NCjg6vjweNyW7Mb4NHt3MgBczXgaG0eh3XbC49LKCmDMwU40RZm0SzmTW5DchQnGZBxYHgf
GKo4+pr/cCj2I2dOyKpH3fKOICT8G/0A6aCYMyXRbNhyw+PWTc3ECTHEX/VppkarXv1NrK6m04yc
LHziXU+hEmBgyidyKeM932id0pY4wtu7xzHnKgyMkHWwcaqMW96Z6rwL0ByePGkUSjkAmZoVFVuZ
waHo7nlnCbzZCrdZBu78gFH3cs+X5XXZAM6Mp6stF5CSJe+E+hQvNCs0INRCBSWaibkI6a3BMoZk
0QAdHIzJxYdlqPLjdfzXdwJKHPE3wpV72f65f5JQtH2EMNqDdPI4q5TlvA21CRjt8pqw01vC2pQr
QFx4YHpEakht4T6QwYI0GrD3p6OCSXyvVVDbxH9rG20vPuVz+P8sRGDnLF8fCeVd/vCR5yEhw91U
CmS84/atJuOEI/d+60AkQIblt+CQ+BlhgWH0yaI+7HdngPEpnya+bKflNqlklkpTO6yMnulMb3ht
YHXyvq5YKFu4xFHlhsOVdkbxU2iOzpccmxehO9jr/KZWsWLcKw+GMHKoN+vr/UkMHpLpFUNRR7B7
sZULClghwxDri6upnIr0hXWA/n6ygg9QUIA+UuAvWsmtEdqpboeNhG/KGuWxJ1F3MDcJKcinTSte
m44RD1sXgIZVfTxwg3ra6JNM1UtPgqfWJRqkXXw766OToM12omlg28RDcIvHZNNpwlAub3ZJGySk
nrvi2wxz9CGdW5EcgyIFpxE8nlUPNpqjKft+sTiQLivB1sAWT1wbelb/nWOsEwJ2TaTXGXChmyYr
uII9qr9dBswsl57iDEeLSf3w0pp9VwY4KqsxQmHHHdO+MmU3zsIgU8PTXfPh0nI25+3WVU4ntZxb
zDNQajiL3S3Vk+h8xLez0DCHTGBLRaXNWeena4hBsED633GQMin4zR/wzhX7rXDA5YiItJN53Jrn
bxuil/IRwSh9kYjrzSUw3EGpsMvfbPZKQS1mIW0OmpwaiQXh3lnaYNxzD03OoHjwzBd37q04f1Q/
ssRYuKGB2GrF2wZwR+Kg4+sHe7B1nM2tDr6bOM7+WImVSVDCbaMBjjZlaFk+whrz0gp6XyqgQu1C
V2OE1hQpylBwgpaKex4crn4myfajrGE2OpM1Rl8Nd+OvRMILOqiOwkcAfgaEDdeKK//zsaL614/Z
bEtzqAv8cpDU7aBV6nz6/6PPe0+crc0E6O+K5gmHRcNY4S+wQRIQxjcCOfC42zwGRM0A6YjSp+8t
pVAZLH7JlJZAWlZn4nsuM9KlSkO+zRA1XEjq47MBaoxFrVhJ2TEp8Cw1DLjFEkmFLIlRADWTejg4
PXp9kdIRi+8FCxXimh2NSpefTq6gPbhlzPv7BCUgjpxKoRuPyn6GnJYId9FsHHbj7wYB3wo3ckqV
ILT5MQWuMk14KBsalglksW6+E+5mUpRGFl50eJVnjB7LnkXj97NaI2TMzQ6otw805lGXNHpOwLGa
pw4KEFjXD6CXUJrHg2i0p9VfGkFtRe0XNA/m2GZF0b260K9+lHDYy6ntOjPSBnSlxJYONzF6t//I
rjcJm6qGvYlQxYspglEL5lr5jW+jMLXUZdQ+qTXccHWXsNIg8+DW/V1xRuYfwHyjMhM2JNOjBLJg
ca7/tCrJ4Ak6UClbtf95Wx2hEeMU8OHgVTUc5d4Zi5fNieTn8XhUiEktwPG8YH9Pa1HZoNWIwRTe
Olwg5jYG3crgu/vbIfX974RzC9TdQbm/7jh7Np/lGeEBB0o7EoPUUKv+G80cR4Bz67FBNpYEIVtQ
l/ndmQ9Xqb72Be+ZQd+u9ciWoWaQZizSUVbNAQe94t3g3UYT4TjI1QUfqgkT8KeDwNQ+tZce+ILa
fEXjUPaiswAK1t2IAUt5RFmRbKnhpCnkVu5wqYnJB6fbzlH3BRVARz0ekhKGQi0TuLlrbyr155Y3
Coc1T+xVGIAG3lYymr8fu/8th3PO/lR0Yf9wl4/b2oszWrswQUp1VVCvl0gYmHeVUNiyF9mCi49s
+ApC6V7q3pjoL+tD6BrXZVlqS6piK/6UhyKCbu6qcGn+N0Q5i2m+Jmh/cm8B3nukPR/24mb24Hgd
ptVRDqpN9V/zYocArsUiIgDD4EexJU/r5yXfYR8mhnNOHJJvcIYJ1jGYdJuRrP1LzikKf9LtHVgD
P6AzEudNa3M+BoRj3nQ3dNh8OJvzsR+hPvDDaQki4vb/xBZkoiV1+kLyxUa9O1s3PLiZtuPloH8d
PQdW5FuPmchTO/Yjlo2U9Z1hlh3Uz7+XGF3MARN+Rox7f4BVJ7JAFBZQC7NYxXWekRfrY9MdnZrp
QlsOloK/+7Qe/+GnI8qVTSOvAKTlfw3hTG+fjnq9X7mdjWduKvzLtueXPZzFrj0BWke8K/Z2C7dE
Au+COcA24bvGkvkoXsIkBFtf8vSBU0VvPfxy32euwRGdIK725wpeG1CYsxpsZE1aGmqkvtfOfkcS
NnG4eu3LShWE4BuDGnKRui9TmPfpFXKGd8UIpkpotqwovvlbYz6dwP7+mDX0Lb0HRjtIBDiD+LNR
25H4+srFmIr5UCURXkA0zbjdhz2xB9eNZ5dXPM+R3phbakNBGBMCUAPm5LYNNO5/21Afm3Mzr153
Ws5QYTp2H1qW1XtLchH2Ay+Byz/TZbY/FTJnqB9vgyCKU47zg0tNX7PqvTd00vbh3WqWr7YKuU7u
skZ+6gWlCITCV4Q8fpz5imPzAolGa5IuIvjJbbU+q//lFXpGrhu4OqOh9TotwrztKaP1039nIAaV
JcRTui2LqExHFt57FCUtD4pGzmZDznNtbEfS64MNdEHtwvW85qlTXmkuFzsYYkFsoDLIOu2cKJ8S
qLBTKvnnM8mQggIteJKCt42kUQESLT7w2ZR28O5SNDlC3zj3xZ8TmY0vJ7wqMN2vRL6ABPVRIdIJ
eht31ju84vULknMAipYRcD8J6epAJtGVttJt8Fy8e2HTRBTfwgNsbNxCckSy/1Z7LFW27NfOwszj
/3NgxFeU4GY8aGR57359v10fsMEPyKNAIJAq0wP94G59vpQdgMp5jmgS4YUoaqZdoBsbatKOb4I7
+L+1nQQ1bF8lZeXrA3xBIkSTGfqB+q+UAtXYe75f6zzaOMZYwtv8eepsMhYt7n0djVvwRpO2SloG
84BrGKc+2PrwqyngmxcwRBDTK58fA4LTOc8N9w0VOiPEomgracPA4ZnMQ099PRUTQiOseK90GoBp
odXMZZWXUMhBze3XE8DdKGr/1Qv9ulwzSaSaS80D7tPggrBo/toh6YsTslObD8/bd96ZaPbIMuw9
qpUb3l9/UWjAYp98CT8uRIZ5NlC4J9G9EaTtyAG8Qxga4JQWQTug4lvWyvoi0RkroW6e+kh7qZwM
fYgl3C/KMXyeINLpypgTY2fAYwJBdEq+nqx2/LaB5yyx3ES1RFp80lyW0CZ2M+VmK/LkOIAEHLtE
7yKtFnE6eExBq14f4Z/vhJic7P9HL/jhRfj3Krn5gtphqVuPplmMdILb+S33xx+UrpdIIbkJa72e
Z24I7txmTKpLu4sdnn3HLGFPfA05oOmUKfGkOKLP1shACPWT88W2BHwrKaRuYK8XMANFQHZpJLZl
y1FIpvTnvqauibT18VljczUM9YPQx4o4s2fRo3gx+H9xjfxYcw6tJvqB+lzl4PxnmIhWwJ3cwXH8
uJGh+/w4RbHKFjTDvC8PvlH4io+hsQzKitCwnkaVkdQybph7X+QsSmhCngfGflRJDMGLJFCGIea4
vkaYxlEHS7+5JQUmcfWJ1IrvyCGuesA8rMTZ4fdvKjw/xyPsDufiT2g4Xj7V4w+652S9ckamWWBc
bhJYrIELT8f/+aXKeBzR7pPXi9wObKPmF8/bS1YkIgKZAlViaL/lVrJKMxyL5w3VVUyVtNINGYrm
NpBDJDfIMzrNC/cBPLLiximHir9xEcdw2PAkjhFj3lYDicxkaoW12LrGL/90vyPCoBrd2vVvrJxi
woOvVGawVhpkhG5CJneqUM8YkDF+QFgcsU0RvcYWJLY20YtgYd8WaWVHociknA0PqWhzU0OEnnSe
tEtfHYNmRVcUgsdsrU6Clzf5xxiTv9N/SJuHuWyg6HIsX/egKKRx5TsMZ+wzVa8tdr0WqUQxkCWj
BRyNIUV872VlhZJAsAyPPTwgC9CtKHi2belwW2xmIz1p/UCKFaVJc9T6gPqfVRvaYjzFdkyod9Am
9B8jL2oR3Fu/JND1gHSiTg7TVaHay5djCNq5Y7EzKG/OYrUb9ApjkgxSRF1D8qFPTTIBSSvSY5M+
KEUXzSrkWcVuf14/pyzXZUBKgpfV6jeQXAhlzHLDIthexky9zWieX6OCFwyeGrsLt76YiO9piwIG
IbbsG8c3YBbk2tqd0XmBhwGsph+2vtjBMhcFKTbENHaneOupuvtp1CpLXsLTJmMX1S7Dg+NEOJKL
wZQXPp1SO10Fxx4OXRw/z/fVRIiabdhcB2OOQpW4yZECm8axc81LA8YLp8dEdUMj7BJ9UMWkqcVC
aFZUxTZ9j5gPh8TUkjlyRL3v3wCK9P0JoL0avEGvdEVnQ1+QGMkb6Z5Muwzs2+H5i1um0WrEUyUH
aE7bSPu5D17rXGrhUQbchVWRIs8BaKxSC+ZW3X7xAqKNJ1nslu1RYUEZc/0JhFBjerdrio9OJPNA
a3Z06PLZ8AT5jEC8ijG6lIx5xMpLi8jGuZK2z0Ee78hSmXKONQCx11pFZnlWX+ov3KBerlsXQTeg
ZQVKtHsK5ZGMT1Aot19kVHaOrbM09tnXChvjmBsRGVPRwZ68uhuYk2E+p5Gx2CJXyRDtod6htKN3
220W+Kd0YH/+vFg7WvPtr5hT1InWEzEJyygTCr78WlyEkuFIKEdbIskA8cpoEpiooLQm71Q1GCXh
g+XK8zOZPLzSOyE6DGuz4zrKuH7ZP0WAV9cti3Fb3vobQARPsbkIz02GX2Xql4//xlunv0Gd0HBz
SYqUp2jJD/MFa3qRNMTkESAoxALWfRPJrX6thkHQCmItwD9WFDN0Yigx2dSwwQ0klZS50YHpUe/r
5VeTvy0ayxLnVZGVjpgMlZc1XXewAXDvp/tVz4WnNnBQYudJbadOS+1jSeHjq839bitTx3gCvWIE
ZJ/961ADKMAGiB3fb8MOgegSqTkML55CAQMAeAMafWGS0oz0BtB/TdUyRfSpjt4NWniiAP9WH7Uk
OAkSnfxq47Wq8HX0HYPGc+xj9LRPZuEPXH7Oh8+I0b3kcFlWRYApmaFe5LoKYjq8Wc5TiCi7Pk0R
c1GUEo11pX0LSb3iEMK3X2RGNEL3teDtcZW8bqGbEuYqKZVfOVOL4WkTgAe7VddAqXKyyzJ+Yf2k
BDkdWveAWvL386ShbkOsOzPG/hHoBWaHI0c0hWfR8KliBP4r2GtUl6hyNB3u5LLjg7Vo53nkoB+p
8N5CzvT2KEj3lbUSq/+IWnEVrcUroyMMvOdB2frb3cu5RZemPpy9wuW6VKVJ+w1fA2sbWrvIks2f
9+poxlHyY5tUTcmxc9C0ZXy7EgV3rcjAJv6ffrL0HVjDoxC7HcEOGbC62Zy65aOmoVkSlL/mLYyz
g0ihT0xcefwdLtJ0fE/RZJtEeXoUI5P5/2JIA8cF1kthiKmwKKhcVhZPOUrxsQKtHXkS4vHnxEfh
LsydmYed2b1XuAQjWypIgk7GT8B847xMqcBE1pdKP12amjDLfQetIn3dVnqJeRm6boy/FV8g28cB
OICUPqjrMw2dUy61w+QOMMRNzLIOwmOHzgZwS8SYdzuUIvVw2c+uz2XCQrYxHzPJcVNzKIlD8rLt
SrQnqfo5zHxO5TxNHHYzkG08eWE4OmiVXDQKFuNvWxaC9Ee+loo1fYjzmxK6b40CbsrWKDNz5a2E
JktLV4ugo+qwXSf1DaOlDxXjxyeKyMbUL8+VIBKfOYMrEGLTMPAI96yNhBSfTeuZf0jINp8JngTW
4nq6wfkI1uF+zf9VAm9EgxjJ04e8cwm/HtdcvqCrX4YdhyfpkB94+9Xkv7jwzrQI6IwPfd4sHzmP
YI+OJ/HWd6Cdw1LCBUC8D8Xradpvox9hZex+2oeQ7o0B9Xkn+VFrRzQI9qyCW275OrYc9BQTJ+RC
uFECv0onNUzRu3HVb9zhnK7aYzEeKf4AtTTz1RRIaLUlsQMTkivt5fQo6jJRnIJAN+zfVzlRwMh6
1sk1QJ10aWb2vaLk9l5eYzmTnKvulSr14NZQHPJQIwf0WrM/z9Qxu+l+mP/L4txDMRplItRqqBmS
aZ2IKc9ZDPaigIEE7V48610sEhmVYuUKiCCo4ECSySx7RVITYC6s0oa2C2ohLyhVQNjI3fS/BnEV
psR31Lu0U2pHL55KLIe5Lw+E6/hPKrg6YkBSlVAloek58WFz3eFrqBmpnFGTujrjZ9JbWu4EecVH
TZug38SGKUUtLTNEhtrc42cA1SETA/p960db2nrAQLTDMU2GROZPTX6KsKDTFO1PzsA9lCifiBgI
98eC+ogBNOlb9BXsNwvyjWtUn2mrrnVS/+jCedPJW7VBrhw4onMkCbK7S4vCPZIFIg/AFD4jyRVP
uhhstC9EGMjZQfeuRWpssHAjDpq7iNMp+mY04ZAdgMC2MU0Q4wI+bPIxocn7cUC5hYtwWCsq1vhO
zfmWmiLTqDsF+elMKa3/SxcT+3GOQaOB3IcIQUG0WLYlEKurdTtWT+3Y2//GC6iNpMsmI/YKhiM9
sW4g+kRdHvD4f+Xdwc65qN6mcj2/VQYgWBMMCGMLutn3oQFE1jbdVxx1+eVxyl2zZJUpwWIbA8Pe
zF1hMUPZ4XFayN09YbTEUJLyybljrl3gexvztsKDEqOR9vlhvNziDpOe8zlkTG2U5qhDMTivAG4W
BcIIBWjxvVsgCoMuLDSzssxE2BKx60lxyAhW6m7qwespz+wR14SQjFNOBSZQgJ4gwstPLh9gz/MM
N0DmAwC5lBal+e2uW7A0vOEr2VRxD18dd8cimbAX/il0isHHdUCosrJGfwtxe5h7kIiVk/mcv1o6
rj1vnKbSEc6Mw3LZL5qfDQSu/dOOxIkE/y4i+H+pKKrIDKmoYlLAAuYE3i4HrvjCRzOG6AX+3DgX
4KBJRzDozxgbjD+FrTiOilPXKToHkGy2zxLaxuqElBgWfBmSp9xEwad13nHbMDaOcl1Wwn6GcMib
pajBEfuVlZDLddGS3s1+ua7Q2lLKsxbBD0KQpnfoJwWXSGwjg3dcYCc8sMgIdE5B0fQePFpJb2tf
szFu0Yq8pkQIy2Zg60rcLde7qloVcp5CMh1knOvkQZARVDKkQuwSzbDSygTdTh6RoMnokGtPfjzU
2KJDraoScjEsHFzlQSSFuLwTeMag6wKnUTzd/bwiUylPdHPDxODYmqKzAE0khMHYKSCLku+dwoB2
XRetINYwF74EUQ56MpjgZz0hyb1qooMaAzvST2W7MKhviFdIm3AcQ+j4NvoyUFl3Slxn9b4sXvFk
TIO3vf6DCHReH6kIoNQBE1KjTz8NIfM/jF6X7xl6aTHX5Ogm4w+WEauoD5tdJ5JQEUbOAyI+A212
89IpmZVPKCQ/3a+NmgsKGhi7iB8boMnez8Ek0fefhJIwAlCbryOSnSEwUWK+l7mVscTDgQXLzLCB
5as/E8rKEq2TEbYbDrqH6PtDaeWp+5t1nvCr1XgfLg2av1R0EkregYKeQVSmpLTA3FxUKgtmqCLT
VjgUrMzZTfQEzW+YsL6FtPQCgpi+n6nESTXtEd5kdHbuUcY0HJNt/EhiMwPWKX4Q54P7AHdO8qJV
e4Ie3MD4J9WPL6kpcfoRJSKA6CK4kBPVFqlLoDR1GaySBTxN8UaUvBY45XKa/pENQkioAPJ5tORI
VG8Oc0+KnWync5q6NqPk0oTDs17rQPB4ORkSL+yDl8+wRyB5/oRV4jbk5BTrHvAHrwwS7ULkthSH
02nRlgEdYnnf559tEZvbH59rA6YflqgiebpOIoX61K8F2K2R1BQbWQLpZ5XL/t2sSUFQWMqEhgaT
hs7Eak7xI4UnSNXpJX6zV2K2s+b3d200jGH7RLgjv7I3fbonceCTWCWI5iqE88/3Avlz+IbU12KA
/qyv19x4a0ZphdK9+ADgb4NO/Sp99HhTy/IiHZREnrdbCM35iXtn4hYt3gSATtMFG/ryivihrCpM
EimKuDX2e8faXd1EpduGA2AZ0459hjv/g9jH+8vOTCHUblSQyrWn+Tr+KoIJi4KRgrpSw5s/ACt0
U75np3w+SuIDyesNDmZvxd2zj9B2Jdf4EthC3htmRyVuOd2wcuRvlt89QxA034qBJMJUxmlXqH1y
E9kOBQPXomgHlsuQPaK0MymxfB0PKGUsVEMmyg0JTsvtuKlXlqyp1sOvLnn2LKM44Lh5TVAQaX+C
ej+Bwa7NJnVuaz4o3K7gZsOfa+Q36uEBuvVpirM7hzjGEOVJ6a2ZZ1dzlytn8w3Ud5/f3CKBK+3w
GGsJnpAIymIJ6KKqqVEpzd0yTHY0amnz0BMHhnpaoLsr174AGpe6rffSYFmJtggbqWUeDDbPL1gz
LblXalL9KP5EENtnUoI/UK2v2KlTpXJ/s4YmuNZLF+6tliUwFta1KMI9lpVetjcTeAJMp5TFxoWy
6z3q17pK9xA7D1Lix8uWp0bdn5LH9WYqmzAmNC9jYL8YK3pqRsLZYm0oCg4/87zd35R7RXIGw2A5
74SPSMaszKZuRz2Dc587VG9Ksno3E2mS/jRY6R6ndTlaBjbfh/cvjhj70khBZxRD9LiH5yI6neMI
xwp8ASZfs71JdhrRv94zfdhOW4t/Vn86Eruc4yjwcl3mejVzAan/VKHuSxNFsoHpiihLgpRQ1mS1
MVlRFn+VPUWVG7TBPSPJqfPxiYPvmEf7BpemGya9j/fpCVT4h4+M8nD1Fy7RNOaiAWCB/50S0Kyh
Wj8sFBsDzE4OvVPkUhfdO9kwNrJnIx+KjtZM4x/zsFusJ66J5BCEDwd5/mLOooAp0kgeaZ4M0019
7IAsbgx4Ze0EqN4DCGLQQpFa96gIiCQYKykf6mjMIZ3GTMeRRqlLSWXdWtzEK0SzufS3RV4Ps/EB
KxHidYa2t5zDy3PqFYf2G4GQt9Ki5CeHdCtMiPWWDHLfQSigtpDEXjvlBYI4DLBkvixD485nJmp/
lmFwQhYncnIItfW4NwEw15W0Z0sleX1HgoXt4EQNFysbbbh6jplpj/lkNqN6tleuSKWXOq/xIaSC
HBo3RGqUahFn0DvnlJP+8611FMiEbhFNJjquUpu9PxDKofwgN2MUdlOXcxhwVBR6mU0XpUanB+HZ
uwer4aOLjfIKGnuq6D5XQ3znM5+02ryTfa6bZUHM+kGeV44kENjcJKpWVUMeTuIrZTdC7uhFEaMZ
AIW+PpzCKQK+aLngQMms/GYgXopnCIwvQWRQkyZNJ12KfwATNzlEOdpcRjfipEkB+m8a47JB5yt9
PcmBtp0snnxPVIKUrEz0oAgOHKAeJ1x0BU8Y2gVEsfdumJXwJKIAW8jFNatOIh9T6Q6oXm99/uvP
CPlYtM+kgzX3EoHMUu2Eg6krjh+1xNYa7TwWw8x2htg2tM40ZsfsPxFwDqUK8KmXMuwps6N9vuls
GHYNYkgvAvkUZVGp+Y76wyPgQwUROB18N+HOxvSJZZpz19IaXNxt0q3IXb+FMjgdsfHCg2EAtxCf
UfmqYsV72/4WGbv6Glcl8y0M/agRLPKZFyPTf9rEJqkWzdsV/gRUrgjSMoc7u5pgGkg7eWv6783x
L0NtpmVCCQEONWDmQ403ciOsSKXymK0HauklTFAwS/qjIdFhsNi/kpSWs0L9JfHAXOh5Xk1WwEuS
JeQgSu29nsb0ancOi6g2R6WwMLPRniDiQHUKYA2yPxhSfiRfYtnyEWihasPA1OfabieNR+LI2ec/
4eb+l5i+zsKknavMA4WdxsPoHEnYBGIKXacbawJlKDhs0UrRA+jBqb98WL8YIGX4RXzRNcJGH9/D
CGoWTLaKJLUU3XM/SdgnV1055SfwjHRwZxaSQvbzGFkKSpSaI5a87NYEOjy1IPITPYEgGVsIL/+7
NUs1sYp6tla7hP/4FjF+MnGrrItDa4CXwC+xwq6OIEQk3POerQXUTiDkKoq507Gc64vr/4hPISZ4
5esgxokutl2fntjE7vZ/Ns9KslJfat2OO3y401fGxSKJN+j7ii6zbRiCDrKYuuyldyaHzNoIybwI
I0oFC2aJzsDYCpSsX2Hnx63gEvCQB+ucZ8bQvKUve2VuFmzkSN6LCuraOWfnT3hwl3YMIkFlp+mP
hfN2kN1CyphR/0ElxrFcpWgCAd+v3YtCT7YcyA91ET2T0ozIzX2YXHBSpTgWSkDkB9WoUewsuxMW
OioFzsfh2RTNanf1BJ/8uwVJB5wO6gF+I5mTPCfxkBlnoBy73cMD+qyOMYPXrBrp5F5iS2fwoFsT
fueQxc59eOmRJ6MVAWaG/V8qCX3xxkU0uYmsKDEnAtpmnHZVF5weEf1Xk5AA69Uwe71GRmsc8CmI
9W9T8jK75rh4urdn/aGeMY2YRaAelP68tfN1XsHBiGP2i1rzBYzH8AWC7vs2Z0UtI0eS9aGkG+Ij
akFyyj3WppB6FXmLoSMCL15D6J4eu7YXAIg+jd3B9UxxI2Qq7tNePbrSzbf8xwjHoMYab5OyGx3c
/ANd0CMbwU8pL1YANGi884IofzRcPdDgeitNfQiAQ/1nSZGQb1fDeR362i6nz6TJjEHBOD7wZxYa
xafMKxvBoX6wuKOCjnhPE1tBvl1g+bzPI3kvrLNpXz66I6TCgGQnZ0Wv8SF0nxZz7nfckjBt+bMT
TgcgHHaf+ykDaVMqKXppTeCCHSvKG+IxJR/mqCLIqC4CGwS1tbOYi2TzeezcZ+Zm5oeHZh2BTUdu
SFKTcFALxQK1VPTvPcRzGDbOUOd7wRzXPFb1lHiTfN+1yZnUJ63ha8/B1SbFdm8tzNiww5ZMcVxf
xRvpvOSXEynZ98L8cMzB/tTsmTiqt3P6OUVjsEJtwGYv/n7M0DPr1aQxZO8UC+ak3tS+nsuBhq83
NdzeJoVJ1mBMNafUZ1i0Z9DVJqfH48hvxMIlkj2bfRAPbaODv/lLLLNbRe7NAJ8+b1eGF1Crlv8L
9ONOCtGKiBgrilSC9VqV01IeyvAxyGGgyXMimgPCEjwRbC7T+fVP/GMT2mleaCRTmyS5oxDlgguR
b+36B93SKUQL6M05uJCfM4HFJWnbws44O17M4PFck63bG5WTAfYpDO66vbU9Ki3tAd+bu27O7zoE
tJRxOynByKHA2m5Fm2otcp+3eAno8eE7KSei/YKJW8Ig8unRwa9HgXl4p1tHxxa+0Onthq9rttnV
5xR7tGDCDMeUQ1VDdIeE6dFdfF8TmkB5CwdLxWX7Y/cAGTAvq3zdwE9R01Jk2XzwF3iQJ7Nm3qIZ
kqcA/cL6/1EYzolm8IErQdIYUYxKSWXfYwKAJkUfecjwMvovXVQgxkg6URD1BSGHag6lqeXSfKU4
nQp0GnpdosjrDW5lpe9KOuZx2yC/g5mPK3jxFq1BETI6XHSf6lsYkPfPTs6UGbxtSDeHcacvmWka
SwspnJU0wGg2o4j5tyY/E1wKUDT3gsTSV5f6KlHz6CLJHb46QCwm1D2sQRbZlHPzT3heDRYYxS2X
B8eAWTZqZEIY8D254LpE4WKejeQvTVKMcVo5g/q0LvClbJYUJMH1GAcDOQ+vs/+ahhd/BnlgZvJ1
MDny7/QHQE05aVIBb3zEF51ih2pV3xR8nGTP89cXt9BgUfkUTp1/LbCsTDowN+EStei80UU7ekGl
Gv2IF5RSfZLETmjMSIMIp1AREfD3LYYBj/kT5GxbCcqM8aDahq1z1YQW/vN7vf18uD16MR0uG1nc
V5rK8OzprV4MKKsYyzfAsc4idOD+exKoV6BqZAtDOsFYKX1Pn3SYqxxzbfPPBKWI6tJaJYsapufy
vtMjFYH1vipa6ZdS9WVW9F5x+xEwB9jIBdmhYSMTDhiUuWOXDay4Au1E8/FJaFT73GMNSsO88+Ib
6GiQJ6ZeCKEiycNjF3IetYobdFtKOe2pFAnBA/m9piwjb5LstvN3Gr06vxWzzxgZK82op9hOF1X1
/vwVDTFWkGs59p24OXhYScQJnzkdGmIegahFoVUuSzJYBYgGuK99s5rqWKQ77Yoe8T+daNLK7F6S
Q4ZcocZwsj200XiTaDlyPH6pGxATNz+/EvucgsUw2WIuajAJBPZHxkDXOxHZvdRwIRDncJggZ7q6
JuCuIgLqUqWQKb4E6wwXO+6BGfMToHLyaYjvQkOxthUQTY5W9fP1PBnu0bPwpAAcEa0PS0PE/KZc
bEQpNB0wfs0RGgi1pvonG94h7tLWh2l8LKFiOn2kdZ/O1a3Obf+lI9Gd0oQKjuR73DzsJUncAmxh
B5/ORt3Bl5vVCyWUCvC2ot/XtwQom75p3Yp4cTMtbStnhCZmTxvtLLDExdueIZHdXCV4lUM6vIcu
kdXCVjV73AXMfFpDyZ/sVtvCkQrzDmRumJ6NzweHBi3ICAJPy4kXYzr2z02E9hFjf59oorTGk8+n
Cfi3Qi05pDVk/eJU+LTl8l79Y2hypbB2rxGU7pVn8uResN68DRXr4PDKonaS+AuPsNIyIlxy7QHP
vy67kbVoPKIFfyRNCoZylmEuycwKRyvY1iI2BNgpyXqV89hfRA+yXF1fNQ3vIOwppbwJ//nvbkVf
7pq6xrV0TEvKDFi7lXZpcBgP80/d2z+3ThEZDSv4xSkUoNVEN4wBQJEcg5TjLBSCBKV7pI0U6Vl2
a+qPpWGCO4IVrAAs3pEqmxRxsKzgdXOTnr6fUGkQM8a9byBe/vZv+lPeUsy58z8LkO+wkCs5+wzQ
htuAQtAtGtBbyxiYOiJy9/cvnE4SdSbKug2IkjihOAarnkOmlD7yHmEEaRIl51B3kBj/SKatFgOL
dHmAOKWyASZBksZ+QdcWCBzyJemz2saWpeXN8IOnvFrwVvXSAiawe1O/teSdgZwsD1+D4APCkBgn
+GNchYlYsc7spd8OEZgu2ajFuFOxwAfQ73SMHLsh7s5Fi/LTPC87/3jPIGrfcnfomiNUShOHdEXh
lzRhGLjwPQa4Al10mppE6FOltGf7L4cIIzzaNCVdaAMR777otb/CDDzcsZs9+glpsrNx31XSKMeF
jPZwOb2fLdcSiiIob9ijN6mIroj095/vazFPmct4JSmH6Ys5sAR4WfL6CYK3IMfu3GTc2p34tZKj
iVbpJf1x2glRiruWgHJRiHZ8A/XxzG5wO0MbHMgAl0UVGirzN+HJSGBvCW+PZX4cT7YwaqzyfAtD
bVmuiA0adIi4M8r9QQ8a390xEyKhhpbkOF7Fc11xdh7FBGCoVwDuMgUf45ehFAoLYrSw+dphIYP3
lkqAPR8q0pOsks+PLEv8Ysf5mqT+e5yOGjtnBMi6VKrA/Tjf0GkKy5w5bs9dJpmsHNJ4y+HkfgfI
G4pckZg7pJOHFVec80n64JvHJwvwM50LCOKl0hpV/GH8ij1RnFm3yC8nbVl00LdTz79WjA5Bey+5
xMiOiIRUUz+SzVLcv4Dv6hlnTp0E6hqdHymjUrPUJ7TQaveYtuqQR6yHvcz2xchsdNH9iUKzX28J
VY4iK2/ohpZxayaLyDfgDdvOgwKchaXWXSpodB2T0LVY4Iq7YPz9NgL0LAhIpgxkGOdtppfqFsVr
p6EkHkbWi0ZL5IzN2JH4wXz756xmUjyRE8T/xFDlLrYXXvhDcAzwgiYWHPK+uodv2pNlNEantZ1n
hmx4jUF4UG2LsSBXlhYxMEN2GufUGdDrw8YHFYWVLLNnYzDY6dUZ03HLj23vTvGTuKp5Wp2TQ+tP
YmyiU9akfTvSfr5bMtE+mgFp79rkCFTkUzhjPQN5y1DCfr9yFIKqHueTQxIpaXCtANXb6/t26LQ8
1+5T2jbSRjxrvtSgOw4Bv7rDSMDlMtdseKsZ72Yza3/X80ax7yctutetpZEDU8kRab/yco0fdIA4
fHVOCDN5eKWSJTknK0nxI4bx0tbcIxaHgecGPPNOxxATQ63+i44QUtOKSkgCqPyCniSk9LhSGzrO
WPwPcLCNtRWsiSQpMaDO6Uu7AwwgRo+V0SKK+DZeiQK5s7FQcRTauo/jI0OwwJceqMOPOvRfD011
SxnpxsF//2KTMAxJ6Jw6vYpK0kNI3U8aCXamqvMROpehd5tRvDWnFZK4WjsduvjSHU31qom9y/9+
It3yOxPVvfF0C4RGWIRnUk+CTJXpOnsC5G6dYWJqT28w7rgP9OYZK2ITv7NxBcQcjOtHHzxfu3GG
UK7eh0GYk7pAYMdzz/KQlH7myj/HQsHSUkHIaOS061QKCBYDXenI9GAYC61zIhQHo3Me+JMVj86p
wKrRuaATrn2mhwKpOBldV1R4r2bY+YnK6kdThcXAwkb/5GGfeMyxZylKavcJniJJzdIxgF3b366B
4oa5yc1lIWR2KD6Sqy3huHVrnXjbOz44lflhKDym90Hku81bftaNUNaZzjLMvAd75KQZCPNUimpV
Da8npxXjPAxBWowpwQcw6ONe+EsN4fuUDkCICogFf+t+M7vV4/kWNTl9EjZxGdwIfdK/3MaHQvzj
mpgBZfPha0G6sXQgRbuKDDCQ+kEoDqPrOECgYtyL7JfIvvEn7s64A6frYWHVtS19fHkxtEKizVsi
699f0ueJepTdGWwplXdiAqLug0IkS3v9g1E4Uk7c6pTTniSjxSn3DpbX8j/OPogjUPzMDOafKiHw
vb8HcisqcSImkZ47OkaSjW5fsrWOnSXcY/ucqqy50LiUv1M2KEWBWIMoUV+fyn1rhWsgXQP70Pl7
r1ihM15nNRkvRKAmGuawG7AKqf8j7JNL5b3WVowiQxeZMc7HYEdc2xcYRQAhcfVaPeap8uaAZyKR
1S6n48zTh2DuXmA02muYVClI3DRUH/pk22D+hG3qd+o7rIFxca2RDR9On3hkKLFjtu4rKoUSbp94
i9yIH9oNKAp122dytfqaz0qIej4jzoWavLQF+BK3IQcmjjNag9gTpo9RrbOCN5oOElP6Y0/7XT0N
Keskgv+NU9i0iCGVR1Aj6GixEIi3w/kJJ1wGje0RgQhMCIM/HlWP4TP2woHRlkVX6bVaOHK/spy9
s3U2VlxsMv1/u7xIgcHPkGgFixBXRo6d3OQYiynSsAqK8CRwks9hzgFYusGrrYHrLELZ6k6jfdBa
kh7MtRIE3X3YigGnqvdn2bQUPB8RvmrxMSL3b5OC9uojqI2cFUD+qqNW39ymz3dm7MXAKba8jq6R
evQc52lRFslVf/1GXCFpUfAu+6Ry/jYaGS5Ej+oUkN6l9Mxb+Y24V7KvEIu/BTDsYKwMDcwSkQ2Q
1cCm6qmtNKcH/X3Cym/seLiD/qMiZMHZk5FuLSUfBBLa5GQhFUSDcm5qaw6JqNyO/kWANLDB/5d4
K1/IDRjNroqLihz0Q6HQUGsUABzByhg6lH4L8lUhYXV/FbUGjtxbGgwSIAcB0drC9bVRFKWlb0nr
KeWIi06ZOO4eKIR2EYBgRnLEvOLxSvX61jFAeJjppohOLIlFcddKK/eFo8mL0j8LASqwZLVxoLZW
uOPc/lJFPxXPEAZrB8FOowX7DrdchQ5i+PTgRwBiJyzycghDOcV+d6jQgkxMv2NyH/An98ip+VqU
9qtEWKGR0faw7wjfFz831lkvkxEHx7BjLJg5fyA9a0XWydvi17WT+tqFy3lhludB6bIDBf4Kz9VY
sUG7OoV9zW5a8ZWABWJKAAShiXTeP8huMnaJ++P/IL8dO/WQDBjL+KVXBvj317lsfHPCgmUwL/5S
+6dfTUp3nxqF6qrzrzBksOV8xgWy15PWmiRCEDH4i2FSQWvZpRWylCeVDu6nicDAcSLEg3rb9Dl6
/nKm8XPRj2Y+h1KPD0yWasHTmX+ws4ECLaSrDzc91ZsngzFioZvOCq+HjWvZsKzq0lf865dcKPdl
BnJ02qziIZzNypg26vdNlz9x7iBK8AitIlThIvoljs3Kziqe19TAY1YXGoPkaVbdAhnPMr/Eh/kB
dd+Vyqr8GdZeIlM9+YUqBaWEIyuOpWp1YvzYj1U6lT3fCSfnoEaHSYAnNzRvFAC4B8PmdK2LzAth
rxcH4o9mbMvCuKzouYCpEoyRJP7cHLSk4d+fv6/MhvQUNt5v1a4URGMSxHWA/OJhFQiegVT3YEz1
c8GsclJtcmjcuOKfrODcqSMasG6nPsoR6kTn9k4pffH51sV4HE5ztiCIsRGYE697nnVg/y6vS5Yc
WrGNBGrKlNrjifuKYXfPaoNlyO+aoX7vRKTUSHjgaembuT9oVTqga6SGI3YlWEkERAdI5sfIn57f
I8d7v3TavxrhIng4N/t6OUedpF5S1CeJqzzD942rIubQz66dXarTxD7G9eYRzvio8kMnTgTZAn7f
C986q2F8KM0bflqeaq6TIqwdw2D1gg8RMGJkpuvNWk/X1hcWJ74UOy/tLP+1GHdDtc0h6VfpWPmh
KgJnfCA4hrb1D4tDGzKOToNWaP8daci9f1qH03K7a3cPenE5ngKRmD9Ipy+ZmFjUOgTj8GqaI3B8
XtreuKA9F4zf3+SYrKE4lGOzZURD7QEOF5V2CcXkq4swJZnHTQdV1nM7IHo2N9ikYOB9bug4O7ko
nC652dmp3u+QzzN2/q7g8mmtRJM+i/sc60LRjpA+wve6Jyv/6kpPJmWdSZQotrvUa+wgk8XjXDXV
FIWvABdSuPZc5ReM8rb7rJCSO1cPAwMIqSExbMLoxxtC+UZYqnvK5Ws2tMy4Iu8EZxB+69vzNFy1
ZmzqeDTbjm3to9QLd9wgyHo3yvqgojZXF6NQ4PjJvnquTsKmm2cxOec+Jf+4jNhWofgJV4BJ+Q9Q
u8mymVbGqrRbc4NDHaROOLfBFNN+a4oHjjuStm3af2Y+U+wtCiL1pu4zql685vnLAFU81QG8kmDc
fzM2QCLtD/0/JG1ITB7bznCjxS2ox7TrgrXsnZ0I3OdbpZFnpyVG+N2D6L/EeK1ysJugvDA0V68U
8OwMK+kMrP77GkIYHM5pOrM92PXa1/XhoDC3rfCsO060zMNZnVgaRRGlx0vWi6vuI3Fg+gK1Th2o
NT86SkiZcPyFbfJ7TqXKCO3HZhtKuwDzyq3U2MckAI0MDcva5GIKb+87rIJergqwi1Q7cLce5HU5
aTtMZb/6nN3B+kuvBZcg1dNPwRauZAXtZHUhv4Q/RSIJGzRFjHu5ipVMecnWB0TVHN/g3VTviDyK
mldlyv6U//757YTs5yIARYWOHsg3Y1sCDbC61QfkamaNm/aCis3mJQWXITkupuZ0QIdttmWDR/p4
kyQA2j3Srq2LOZRGHQMVTQgr2FPH+5nneM2mSvelmUc12qlOXdLPH3lhR+8eTBml42iveGROeJH8
U1lQhWlL+4ZE25aFxBPfKS3mzA9VD0oMdimWapzIsAm7eq6E10vJNsci9f2G0P0QrlsyQXz0o/7s
pcg78IXunXF517OrdikJT2ViZi9T07xpXaLMrV6WJ8Jf/s5s84YUXmaVhUNiL7LTH61AlYzwc7sl
2OF2GyiDDzZrAp4z43qOz4KI5oBxiAUpxasoElgKVePmOyMtLgZn+KlRPaHyR9GYPrHJIZ+K0m6U
+Ey6n1BPPqTZpRMQm1gGwfc7ET15NlUYqAqjnL86Y0UI147pw5mfqt5AW7SkVkfLseBFGRBvVaWD
FL1pjwCgwBvHMUgLwEQtVNKNk37WfWeTuPzECF82ovaUPV0qsaeHGbEZev7Dda0ERjte8bFQzWXj
fqmUKoT92wgipKyeX0pEaAMB1UMjYpIPCnmOYRTyN8pZupVvcwB3cLz5jXwFxqWH8Rxe6YdACMZH
NhCsUAmD/HkHgPj8xjPW5VW9CI/fKbmAw3lJGyIL+/3/U/gsDhBWF8T2Y7GrYo6OQ+Qeb/w/+Tu/
wBw4vavMo9/fGq2y0Sb7dheVq3i2nd5O+sL3/DxOKkyiUE+odXqQPwwGBo2HTIFCGdv7n248r4PF
tq7vC00BNwOfWsOtfa0T0p1WMewHqQ49RwdjMd8mSmcXNw+B2F34/JVgA27ErWVzTaBzrGkFdagk
9GpiTOjSmbasA5MTfyZv79xCsf/NRWaVr3AIg2UwTyScU01XIAof0qZ5rdEqGbNwqD1JiZAmxPqj
YtrM9Nyd4qDpXTou7AHpN5QJDRM4F9tcjazC13JlDznb5p8vCkT1l4mFevKX0MQSQGs+83KF/xv4
9Kv8naHskRihS+XRX3osM16hyVQq2AHXAFqfuI34tY3NrXEl2IkDo13BfB75fy9BnHPZAD1Plwy4
AvSWqP25DMObKiVnxQ6JtIrvuwRjkGPQ9JjubGOxb6U9+/5XC2MT8vvmY9TCjysteuNOP+zRQ5d4
HZfDQHQdgX9dtJHA9AjH9qeCjReyCUDiLPJzpElIoCsB7HHlBtP9Sko8HAP/GOrD4T7b6VoW8laN
QidBWyZEZ3LmR5+cUgpJcQRy74HWD37yEnS29/PaAI9JXkLaFTCylsUfVDs/jsoaUuE7XGpIsITC
04d8Lbkx68XeeR3I1nK5VapZLxH9/St2dAk9IZNmTchuhtl8zn8uqcT5iPLIHAAshsb49pS8z3yd
fH+ToKfClJE7/48AuO4lrzkriim9jzF+Tjq2GFGd3pOHtx9wn+CafEKFG8/V8kLlv74nHHtsVuJF
0zs6mjSv3D0L/JwfKqyQD3fN4iAAiHkWUDyRjfC7o82M5pM9PhmQMXhceTupuEM0wtGNdXy2sOGG
IDUwx0FuiCXVlOIzdHJpMDs4Kied2FjBOdPchJBCHibWo8wRwkUyCSz7+W/8PeY9/NoQvPTuXDEF
4PjU7E0S6D4pXeyhdQR6mkcuFvL1/ekO1zqiczh8VViRYmil135Z8CfouY1HiBa7tMarXxDpVLss
G6x++3I2KmFWcGD/Qd4ToN1Hws0CIKBPfe875WXZhwrAqnMfEp9TKNsNOtb/fxlJeewg4LMMvSC/
YH6bzLgOzIUrpYuPNsx4V1vB7EUYyAVFIWYzQsv/Gh4gGpKX0mkaiwkJAkV9CVC70h1zBghTsHWe
78knubm4KSEOfTlYwUJKBBYjeeoC4PjawQOSkyopQUNdu+2DxgHPyexg/qGh2RIMDV3IISWVIk56
qzWaAKrwD3ZGF9nKofjHYbLlGfUiZ50Kw9NKh6vfQbaRxbGiV+fcfLmlTLtm44QpAn2fKGBbbLl9
JukrFvEcc9rcwDP52RVro1CovFbcP/aoFPwFkusFhzbNn00AHr3PVVa7vtVhQ0xlloEKgmrrr4H7
sg15aNWgrd8AgHjp7JHrxXHpxt124cgTBZpWe9jbdyRXbot03ymk5bNl84Bzywux4uKHag1FNaXd
/g0MfL+xBxe+jQu3wy1/pXk1paB1mTV5eei/rge2ZGXkx7Bwe4irmgwWw/cSaWIBLvsJeZ1BUL03
OfZuhTUEiS24B418k4kur/flgasIbwWJNqqhu1sSAzZWb6lSD/ptmknFSLij1ErVoAWaaJb16GCZ
0olRbCPtJ9scMP6c3NswqeyBK/jFS4iYHWK93AtCqy/2mEHttrZkIj7pqRfzh3Ub8FcudjJbDAeZ
oy3QJuUtwsMXVd9UCsQUnHvlrSkji122yV0Clql4HPhO3OsQHv6QgIXRoEz4+zM15j4OS8emOZiW
isFuiNGwCDE9bf1uezeChCBCHKxEdUDRFexqLPFaw0Z/MfGUceCspwWOYVbyV3C2v4+DpKqKNIYH
GLUPUzhF1ZzNr/p6iRyxTqZrn1C/MQ2cvBKXI3iqCpGWX1BW6PUpG6Qg/HZjyb7l7VvD3CGB9Gqo
C5AhfaLhquOosNeALt/daoy4962ohdyGEK65TulLb+x1trNTzCfQ+fky4LZ+d0wwudBSCB2B72wt
fEkUFmZZ6plZsfDFa9J3IYWgQQx09/Had3jH/961ZSC17Liaj3Wj/eka2HXdedzyDd3nRX2oJkDW
yzeQKjaoDNxlYUJ35OnCqr/KYq3IVp2OYvZoOqjBYJXEnRyaJTvFRlrjsRpLE7uFkJAI0YVuaKX9
PdFa1k6e6b2cRRUXUodqwSwZPYai2PJOXZB0GJm2J8Ak5sfYbxmOWSMT2CyiCJFQH7WZ6jhAEypY
S855ur9bq0+NFdmbyqXzu1UArRsiCFZ9z7NajXgtzha6V3S9NIdpdbFNtRkaTDronipG+1daR/YN
Z0ArP6jDYhpUM10R32scFUZGjsGxK/qi+TJIKx3HLVlHV9yeEqJBOE9CrM3YJbzW52Imwu+vTsVI
tPleTz/UnzFiJWo89qfZobDldIBJpmc5Kvrc30nR+z+vHF1u4xPqQw62cxOjwgPWuXZujs/KS8Yy
Wvw9TlhI7YR0YQEJNcLMuIiYtY/PKb8tg3jsvJ7fcTA4cF0P5eNYF9Z/TiIafXc0NB/U0ccnbO0W
vHDCS0xhlRUxbZxzkfMlJMltqjzOtFlkk+kwEY49R9U53kf9bPbYpBsnO7+e9BnG257ZGAGyR4id
p5GUMTMWFVlc43pi8HFcmXgZx0W6s6yYfNsaSSLs5JyoVK5b7oH8H9XfTYMDrdbHYREkej1MGTBR
Y9ZoHHC/y4TncpO8ZZPdiUByThcgtL6uO7A+cjsIezgdiqZTWkS6o1xki5LDZ26QW5DWLi4tWVpF
CuNIk7Ts6VcGlez/QGRCnewT8SxG+3TP7/DIX+ADxkVlytfF8BI/W1nXCs5yBK4HeFznEGW40uEz
RoYP1Pud68PbFenxTWmOVhd1aK6Yrz5z9nBxy0SetuPemZp1OJk42SAWmg4l1xfuGApLLMWZXbO5
uSSvUWICiNebespWRGLxaV1QehG8Uyun9KCeDkWfILe9XodZ1U2UYpAja7CAW46VbRzopzBQCd/M
76OXw4HryI0NcliAO8xhmJJCZNDJZtAc7J41ovvjVwoD/cCi2J4js7rnJblz9/k+meXOMIlkElPR
AaJjEpbsZDuYKKYF5lwchEzOnCDtU4vLy83G2ct3K5oMDzwAH3BkMMGrgMKa8vY3UJiqy51YU/AS
6CzynvwC48GtX0SVjw/y2Whq7DUJFkJoVNUYvn+U72vU0Y5Mn+5RtbRCxR3kUPNeUbU0c/8Uvp6R
Ek2o3dvb/CbMOzZctAqgG1IgCK6Fr+vM0e7F126BTw8Txo88KGmWxbtIoACh3dvcHePfm5hMW9zn
LkGVSXGPU116pB7BcHAUxpj85kZ3HzoGW3oqeDPrTkYAzBcyY6qGOcEkpcZ4ZwOyzHj4dtohrnJz
515o3IKYanbBmwg+sqIxophurJlfcHchjrdlMdFAGZE10/e1Q+NIgw0A5kJ6N/6DKo1B9f6Vpess
J5ktIiYS6yv0CH39/nhatlfVEYt+u3pnGwgx1GxkhtrLO5QPtwCoSIwvuzHUI59Al8BCvgZIub9V
vREOiSg7Wv8Ldfmh154fe+bq9zQMMJU8THRes56YGyeA168t97MiJyD5d2MhbZKKgW88KVB4ddId
rqk2ncdx/tKjmuja7kqN1HD7XdcQt4ZoJslQnzMxdGxOWWlvyX258NPXQ9ZpKWy7HkfwJ+WAVfAR
jcn7ZjGhJ3Ona+gWRscEJxbhOAnJ7oxJtCrtu7F2O0nsb72OOZcddzLg7M2TVPsr4TltVdBN/0+I
1oIPlcT9aebqamSuWK333A97/emRUcSqgJzmCkka5gPBisLDl5wrp8WTIMZDbSPUaW+B0AowMOve
peDK69Vv8kMSh3VaVPvEZfXESyTrO8UPLysh/t1iawGBnYV7lExvgDkSEUbp7SAP2sTD+gixyKZ6
JPB1ECT+z7MYB9QPxVXkzLG1EAOzcbAAxm7w5CejrZpa7df2pp+6GLxVNJ1dCsj+IM4739bNT2Ns
Qd4WxCnit+zkLVqJiCTntv407oULwrsypGKWI91tWfSEdXhURo5GyJua/h9pK4AlniCsLOvAgtYr
KNaWIoVAZGEFioVA//goSoDdfclVc7og+hUkuBCtkbLIV9WlGoRQpQQcIoo3UqJPcHa07pctIzam
dfSLDt5c4omPKDihdm2Yldo04Aivn6SqLlRJO414Z/zFI4frhGUQFZA/JABN7lMXNZ1QK2l5X1eU
+DPC9SvqjYYMPM56lSsbf2GOfLwutbKx9FYeAzFtM8s4s+zHZ695wsFHXE3WfR8W1Pp2/ILduFDj
CmQV8YwSnHYddkiwiTLZIBttIjLMB0zfT+GcsFdACgzThQCo/4vPC0YiY7hiHQBOWRZaaF7g+l+x
tdYLr2q+awiQUfApFcRJQSkvkvYyvGnMo9+qAYo9TD+h0mpi/GNJTv7CJcpBb3yB4YcnHgdnUwtp
PF9g5CT7EaZxHiFPgAETf3qbahBI3lY2S1uc3CLV25z97QtSIjJVe2dN9TEVdzYX6cw6wSh7A865
uZgtDJ344CnkoEiNiiaNF6LugOIDfNZv6vxB+xvN9rw8IAO/057sKlAid2Rij4Sn2so5UA6ubFcH
8sSV9NbYltyvG7UrXkrQo8qWuv9QXo+6afo+QTa13tBnk03OvCZiJgNRI2FTBqfoO2sCTzSInirb
5MZmhW3DShNi9Yb5P105IfKTHDoUsVAZQzWB8HNSdWm/xxJmBeuoTHg17/AXK9+hvueJUlJJ7P1s
FWVolKCO/O87Sf1mE+bPjh4F0/we8dG06DPDU3Mesph4AQwQKprt+RVXutSlECog8rMAMZdh1VM5
BKdfZcjLgkscdfDS5j4zkj/2cEkkSd9GjKp5M8WOti+pO5A3/4b7IgrI4GXWi1r7zUJOQ8j53alz
BWX0iNQpBiuqAnL+XcgWiVylJF04tWCdJnjFbHCmzLCRiKAHg2ZVJq4CwCRRRPOLtpV5FfezOq4z
qJq0R6Vi5mkRgyC9WHoFzez/zSDe02tJMhyPHeRzlcNNKZh4+wEr50cC5A1x2Ngo8SyJLssYIjwf
OBkYNWO0ZZckQkb7fzuylIJtzmlZIzL+JEBrJ+S/wbGjgCKXjjodbsfW3r6iKWqaTzXnrWQmIU+z
s+CNL5Wr9BUtg3jaJ29nHIeQ4gB8JV2IsQdYaJTRaRbk1OTjghEM+6ZClF1gz1eIozAiyG0dE1Tn
7G2Y6Njdbsk0j+b/Nvbv7UvUT8uEhRTuzJ5EDeuV9Y7rmM94wULz+tEHRlOK2d1Gdq+JeDPGhKBM
GtJj9nFpsi74HvG8ElncdWGLenjtg3L0T5luwI43YSgcMfGSU3wu6vWiUqDY9dskrJnrw1vdVlkf
c847d8VH7703aVf7V+My99KN663LPaHea0nZlLpOAykAhrMgEHY2ltySf0Qs8xMwPy8JiFOxlAIK
J9V3IfW0//tBFNbAbN76ZIlbd7NT9NrAGWtK7ygMmD8EbbA86kcHDtEK48+VQqT4V7fDsMf5/3Qr
E2HoU6KIVctKvyMl2VUtRR1wTfy58jsFHwbqcuGzdaPpPRbyplS+aU9Gkcqd1ZAby2EYUKTnNUas
h50pYAV0I2YCzQ6QsuM//qiMtUruGXmF6B7mISMX8ZlQ58yNmFp1x5sb6eYP3XO5QHPKgrb5I5rP
WUhHOZ8+voad+FyQQdC9Q6E2b8dvB0OMF2JgQLvjg/xZGQUC/4FFZ8GxRG93H1v+R3mYE4vGQtPb
FwDauugpJ4zNT6CELnI8TbfWj6L+n7tt5K3oertx3mNUTfAfO/p9sxVu4L7vnLVo81ZqJppL+ZkI
vN6iavGT5xSjTe41ne0A7cAMqRApQzp9ZFvxxihWcqZIR6hsNnmignPOucJGe+c+NfGGYGvhRr9V
mw5dik4wXTy+L9i6nCjZtZKOKUxVdc+hfvca9s51l/UH40IwVzENjcEFEGJmb2Pazm27a+Puz+Ni
gHTcxv3iUepQS1Z+23Azcr7L+qfPGKCdbeV/59aQInMBW8MRPjFp8wTj9JJn+whQpXIYZT4f2WcF
tn+xat0Vosgc7N8NeX4PpRVo52HZehKpKGEy/VzEavb0PG5v7qv8GB9c9iylbedXdksuOjgbxNGY
BG7qir8IrW8/86ff7DDuC8QcCkSh0CepVeO14CywolVsZVUr7UOUW7R5Sqc9s8ysSsBPDvJkEedU
8lfOj+a4LxKj6CqBJG9gnA6UfjdEFJy7W6cBddrk9Q2OAOY5OGm0rMP28LgdvLqyP+nsRpQjLutF
AtEB8oFsRq+1Au+OhU7zX4aa8o9WTLs12cktD/jLBfp290CkA2qgT/zxRZSbOHpW0Toiido3kWqo
DaO/NfQYW1arUrye71G+F0wI/FTBAKqzI/rc34Yk95Tr5o6dJLkRF90HZx4l5c4ZYTGf6DmzUuCQ
+iHJZU2UaseOpZ8rdnuxMrnsQjojdi2cA7zT81MQNZHD9TnFx1ZzsQMFJ3g0tRZuIOEbLIX5EAH4
lUF0Ym3j9rbSs+qm3KOjdNqU3yRZ0+nfLScSl03AQFHKSoBGsMLpJh5EsmzouhQlGVDYMmQ5cAg7
e5ffL7IiXOzvFlhXPBUNy72FH9ltqlti3wF2PL453kkms0g+ehQjDt8MVhekrOAtgNwYqI0gBQ6j
1bHTUPVaYfWktqu5uCKCXcoHorhxshqoOx/HPhBW5PuFbCVa1g3etBCQhaz8JG1DwRrLOx/m2nYG
WmdjrO3ErMinAT6ZuqFjWxKZA+iVT83caHLAbQTxpETQazUDnPE2cbiC+aFpoOUL8ghziebcD16q
j/6acXn3uZ1PWH6PQq/r5hk0vci+oP+uPpDmCI1olbktpxjwhXYmgwlTa6bohVOmkd60DM+DLIZP
CugxCQHQiz+9sZPlhZdIyP+v/iNXgvUYoAtHWWxUCQAdmCJEhMzA1wBqpZWRpDpEkq5D50BlcRL4
JN36zjg7MUYtsBic7FwuQ5jBOWjL+Yxnrb/Icnq0jSdyCYU7a74O7P3mj3uVmHz8XcX5hSgndnTQ
8g/uZFpGdk9fu8E70qnoI4DdBqo4vr0/a2qy69oL9ikgJUKEnA/fF9qQENMHw1t5KOfoFosBvmED
OlM7ZrGnsrnouC6frTWhQrKMNk4mMsA+2W2UUEwutDzp46mkRair996AjIWFVNlcyp+2BJDFAiv/
nsjYHKm71GLkbYlGBhGCRvH9n+03NjwhCZVxaCGVwZspUECSfgxU9qHazFP2toCo12P7wozKDxe9
h1KjV/Gg2+SYjFulJIQosZqO7PqEQjNId57mLzXMMPHQzWnYBGag0kl4NwR1pHAYlf2EV1vzxRvn
ZNF5Z2gHM98Rnt20uS5fOoB+N0h2lFxNKZ1sdq3lv2C/Z2KRH9sOQapjZX4RMCIfzQC/quV4vsoQ
nneXvlPageyULnZfpy1yhznrHyIbWK7zvh0YGWOXTW/vxAlv98m0Bx87NnGlggQwrKoxLvg6SUh+
WXTc2U9CNE4qhlIsp+hM8hyuILa4+62cmsGPYXuz2/wgL4tuyvjTJKQFKOBshsCoylAlQTIVsiZG
6aIWQGLpCG17ZUsyqZ8h51qhi7JB5X/nFAkTE69MHpowkUL0gNxsNsGpT1g6mU3HiJ1K2Nqv3CP0
SrXqBFY5c+vXhWcShRCI/BNY5hybRX0HjyaYDjWthp1Zq3A1cSJuHz2xw0jOv6J50bcuLEj723kv
JjtynkfnofEIoCi9T4ZgNsafqMyVbPYAdJqwCWpvmH+CYjPArysdBU8oNsieaVy9muZSiJkG8SM6
aMcE4rxvN/uRx6IXagUD2ubU7aZnXIfSoxsxGzZY9ayoPylQ1PFgu+xiUb5vc/7StaAR3Sqe6UvU
ASX6I6Tjk8S953knrUZAq5dvYAN5C2GKsquzIyQf+m6kX/1XS0DxqJ1H6QJ9lqBkmnKjlRONZB/Y
CjlyqyP2irpBvLuOC95lJS9OpynYlCZS48L3ZQAkLjktLoyhTBMrkGVEqvlXpjoOTb3YoQWU63hL
UASd3xITG+zWaNUm8V/TuHZe1nRgSv5lJeYlBrIVWoqDlo3vNNs7eo6prnQ1/mJnl51LMH/tW8eC
VkX7Rnzz4nmYKQ+30c5mvo/cPkT+ztMgHomBMOYgfywraJzMEIT6FrHw4+8OEvTQ6DQcAGV8+kGF
BR9fb/jCnGpp8HEirlNz5aa8wcMpWv1q5RvK0TvbvexP35lxCi/VVj1hkSXCQj8KOhh5wI15t5BM
WVlEXm29NFelpV4G1GpRIB3YwSVCHzBCtEOLYXtiJnW6gqrXQmOod1ywe4I0MMwypHIeHf61/eSc
ItOYIK88W+xt+Ug+XbHmuntyJQ4yR1MlyLoBQgronYySUam5fGNoETrPk1g5IoJGR4nIFxfUrSpO
saWMUjYxMtubIMNiXdw69rW9Wn6hDWa9VUknZrjThpjgQrnzecFfnUrINbmHRHd3xlwHGwssH2UQ
+yqNb8X4RKIDLPwqpH6Vn6fTdAoA7iS200lP83bNnFbfmZdIg5pxYDiB8TLh+jmH3uNHGNuG+H7t
HwtsO+lXKzUIjnQeXSSEFZFlXAUN377TAzKmiY+vx2Tfk7p2N7RWKLdnAuiBVnprkTOhJgym6qvK
UHRJF4+zTRtrm0tHHyiGrXiZPWkmn42ftgIcVuGDvFXlSUgUNYEF3LzTAx4iQPl8vMSowzqytnz3
4JBE5R0YUYsK/N6QTIePqyt08HJVx7TZEhsqMc0qrZ8kNRzu6lG//xvUhLsrmc5JYKGm8qtT7ICJ
wPqQb8zoKBUO7FXkVcswtmrz8/krctUAvdsqEbGFp+ic+AT1cj1hUE1a6pfhEBYtNI6LxmmMtnYm
EW7Me0DVPjOFZzi1tV8Nr+nr1eAO15XMfS/8ykzJcQNMbqnLtfxnkcoXJEk0WWjgwghTDrmWxZUZ
aqw0a5DJ04D+BbsFCSh74SCXaNYMYAiJrcHxmTqLCtU5TvQBxyP9YZYDscuXUxJRCiwmm083x00M
lG8cHCQ4NTWkeRrURPEZjPgYlvTPF19j2oAMXaDA3CHasRrazPMnuqH7Posl6mefiSEZB3IxS4at
rVoPFZmmNEszAJWNAGOu6wqSbahRsmPySXh60u1QYY095ZvRBA+E8F6+5vfeY/Zm7jB7HHQ7wBtk
36OedUq8vZ0+glFNGPsWcONbuKNa800mnfltbxt507llaus1W6Zuyx4Z0d5tssPCEECWyDPnvspS
dJS3bSn67L1E7tzy1rp9zZU5Z771KCcl2VzjY+3dDueVBC+eys/tiOSlOPi9Thh/l5wHUYkuEr5L
GmRnc7BxUWAXEfBvMygprezTPFMhaGcpE6WNppGx9oDPh22bh5NqThj4sOfu1/gO1I9E2hOUuwKc
YA26cgS2omRbs+GzHFl+gGG0wsIzAs/LZr+sZykT+Fjnrw8QJWuP2CXvRZHX0L4YfqA1ILYMJTZd
/TqU1kaIs78jAYrkLcLvX8YpEEhoKveW6Es61xKxykvLqx0jxukkOVB25GKYWhEwfPLHRMNxQ30i
xs7seDqY/ElizVYq1e2YROC8Ol7JO26AvYTZGY+zoQjXktRV60+p81fwDUdJf3wy3B547O3bpwTo
cbdxXP2OgzLtJXBIGPS6Z8bMvtT7deKM9eFHWS4v2+r3B+PQ+0HIjqK8jtRDyv0kfoWkwey0TmC+
SOmeNprlpw0wMDFhupZcWqkUUzkjgmyR2YCPiVdFfyfDVYIA/oVVMjiweMIqfMuDq8+K+khdppBt
mjmtwVvftigX9YjtNf8BS2iObpNtLtyUKU34gjcz6AnRG3Wbj4FpI5oxm1LjFMfffOxg+0aYXsBx
ou4VYYubzFu7xfLGC2ApxRFci59Pyey1PwW8xgzR/9qevO2xl0o9qbzkIo6GHdvbedyfLUJiTp7Y
1sIFIquGmpvpS4VQiWC5qWDc62AubK7rT2zq259riOM99326dW8cvt3XpfBtWYhgXuv6XZPVXzLP
2abXxreLVebQmqRR1WP6KaJ3QKWKr2YxD4rTVFzaswSfnY6ba6BKRxUg6EdXJCuZ7xYZud7v0H1S
Xx2d5VMuDY/xcyTOaBhoYnIb5V2rL6V9615UlkmTfPyozrwaswyxzErp7ai5A46k3HUDrhMoc4E1
ZFEI9VJQRV64wODkEemWoFAy4xvUuJh/mQgQrA+g1FDe87EJ/+zxxP40+rpgQ5/YlbfDwCj3hE3n
idzAOhM1rcuvQMYp9z9OuRJPhglv9beGXyEpK+w6ezTVdo9FT1nr9QkG3+ie6fmaEIzlCbO8nAbx
lkLTMVcfhK31Gm8RiobHRM6BZP9spfU+n0nII40B2pC+ss6CBgW8R5aKt2YVMf28Gf0y3gvehtjW
J8+yUTXaiVpMywBeLj3e5YuRENsr2y8azUoVbplw0klO/3tU0q4iPrfZzpogZtB/Bh3EqNABN4A9
gDOcKRVR6kPv7gI8SC960zOV4ZFPYXwmI3xbMOudpXPPwleFOtvOqaEFhRFxGvtr6uXPU2SYnxv3
bWhfNDo9/RydIS/la+/cXlS97Wl5iQ6vPnsns2XNh7ZQL6BxCaFQKfQzaNxxNvx9QzCglVslNUSN
zExSjo/N8pTkztGGTxfU4k/VJWA/IvESd+4CaHDqQ2czbNa3OT1WjiaVbyAOYNv6Rjm6CTvDFojB
Z9KbPrUelPxOihbcDwlrWnrbbxACyN6Sxmbaoh8rLot+4y/NTEDj/flr+sPdp5e4IJZ9ehR97muC
/7JOd0JJ+C8akO89YOuYCOZYriP1e0NOGiABmi7L/4WWofWcY+ZD+ayxbMIKMLBRhTiA37kI2xSw
9MJ39T15y2m8RgmSl0iJaBhm3DWJjR4KWNhASuO2ZOd0SVMreL0sD9dtMK+kl1DULnr4tzVrhU/z
YYPeCwD5Tb8VPaEH7b1zaPHbAbmlXXSbXtz9VXE/BLiaPRO3/O1flpE3Qekzzh+uPeTDGiyBnbOj
4eE4fFW8bE24AhIwvacqV34sY8SGNYxJVzDcx9ul0awot+29VJVqn05eeO1S9Cy2ABKIdl7dLdZc
YawqLsEgrj3Bn5gYpZgDvDTmrXOvQ4mWg3pZRGM7k5N12VTrVeGhK7+z525wB4yP/Uirq9QRK1x7
FJHZWCGxpCczJWV1R1f4j7TAfGhkXFxvD6pffg/dHLpKNFT9RTTjvfwnsVNUnGKJyN4SQYvtM70g
Cnu3AoF7cuiIrEbXqTQVy6GKecLhnV76zg69EkwpatWc9ZxWOtL9QE1KSxctAgKl4wh9E3WZ1BN1
hx3yGncJ32tNWK1ioO3Nhde/28d++Nj5UVzDpX9AwVpksfEK70ljTNJWd9baPkdMf9u78uqeq4Xi
DIeUlx1OiM8CHWuV+hcxHQBLKX5pzjLJRHIDaFnFpg4DHvWwPbuMEDN/gkp7fexd7T1kmOQEhnGz
IHiF6MfGiUrnB9gniLA8Dg0pX4LYA31tRfFsn6ZqGq3dyGo3Oq4a1h2VlVTTFGsfxowZHQObvpV5
/qikoNQIjPxXA3p6vZ2chDbzF284dIzNeEwQrxLpdyvYiO4RMazaVhAeS7aehskAMZdSqKs+kJYn
Ho+OX2VtS+mp4L4Bs0suCvmxAWkvRq+fqTfQw6RuVkRoCG4YgrgsRqpT/gyhvkTVlAT/8rkOJgYV
sWI9bVLrXTej5a/WGvZbOd56DRbkg/Hk4Szfp1Um2qmP01amexQVGOg3vfPwZ7FpBzLtGsQpsVTd
rZFswnQMRx5xdRtK9kNfdF/mBVdWmQK9gvdQTUpCSgkHWC0GEC1TdN4hXojN5XecKtn4CJFeAIfT
oEYyWnLb0/3jGbFuofkOqILj2tQXmoTcYB9pRDrTUDzwWUKdXgT8TvJqZdnXeFlBvY3zlXX6hn+K
2XgQjGUmpKQfHmIT7K67PjpsgOUJtXuVqy4cpzXs6G4VyX/+tN3s9jHmSA4xEijUHzW6/WUSAvZr
VLcRiWpQgf8EPrQXTUTvNeXLUevYrpmydDrf1sn9JiPNs9na35RbhCQiHVck1k5Kqucvmegm4udU
IL/NgseiV4rQPZrej3QbR05HfTuNhYNpGBZWWU33NxqWjqY2HBtmiI9gzA9D+x6jpjzRWM98iqyo
n6PhMO19rdTekkQlWxzBjB5hT/QxFjWse7gr77T+CSUcreG/OYKOMuV2HJ7NjtghhP2KoWclgD8Q
rlRf72RPGgxo+IbERxu9/rL9SwTgA/2+dDyk4KosP1jglHm23QiQBu8sj2PTYovbVFz46603tlgO
8Cxy4xJ/AGN6UWNzU08ISCvI4cHBo+AuKOltRskymjIoIug8HoUlAg9ohpLPqhjTDFwfNmxx3h4C
nw4O2fwc9ww5+nGd2roimmLuYDOXCmQsJezN8k+DULa5Rqt8XuZX6/W+JQnr9YDW4wabaYJDkI9Z
qXGyUsn20PYbUwCswN0RVpnLf7pvSIzfwI9eIoy8LWe1AH40MKfsgYdRTkR2KLS9x78Jz5+jhLgj
i3iteiv1hqDVcn/dO37A7sDG+RuT7x7OFjE2b1NxpeUmmeJi+hao+u/RtfRrpvapRXM6F80AOClx
z66iuMIKNWFX+bx3VdjxT5tWgMFjDWNny/wSLrqGJkKRkj2VDDbaPRoU8gsJ+CSv8ECzvL+Y/bKK
7FjSNOKcbcP0U13r1Dtqkbsp2tm7qVQj012iOK86QUaXamwX60dwuxqFyzqU8rf2y+vdOsWgmoci
r364Pl7YpaDht/KeEajKPNN4npGRWA5juyx9F7jkQQnEWo2tG5fzirA9L8rJ+BQdlQ2Ctwmd0aIO
01HX5AHENBVHR1UdyeBnSBjcN74w89XiCX+ygeeSzcG6phvbQR3opHqN7Wcuh2IRrKhodolSwPmW
ie4fW/tzAjEpQR4KKN3tB7w4y0RuZUaGYtP+O/Vcj7BbQE7GR9LU8eAOBwDHJuiDosDOxCDBztJ+
ocLJhPt7C/DeioPGxZPGPBfckCiWBb3sBfYEWOMbnZgJ4ihsbhaOkUM+zKQnYE6y4zQBdhaplXZt
AMQdEr6KAicu/ufi/nA1LvPu/bZitvazlvlCQ5gGflhGbw+YPLZs5ofwSPJGSuWhsUYMT9+1BFAK
ulOaLmT/nH5k35MgA1L7k3TmVJLEmsGPUADdXqYJM5K8ye9LtRFD/h/vI2rkYPhp0DokrCIeTWsH
DSEbeLEWquGYk48Ig4vll6c+j/GxhebqwjAEtQh2fXT8G68tihNnWTsvnVUCUB85xfuq3f08fXYD
wr7CD1IwrMDl3q4DnVnR5NTrNolg6DGvWCmhW8FQ3DF8N7Jjb57KYYQdxxiQGWJOjbeYnZCPaLgQ
6xOOcGgoyKtV1ipQAbVc2hTGOb04vK0I2xcqOeDqf4YxIDQqzlJHgnxEElXaYeBNkENm1aVwXlMw
RSFnDQPZk+4fWmx6GzzHnYuX1hmOqMr5YqlQ40rNN2c46P/yMvhz/ssMCCwppIIfufpTv4a/6Au4
NJZlllalfV59RA2wsQ/2rl/TMh+TpCaIl1DOXR71hllI0t5E9HjA9h63PvoFapefZqLFzHZrKxI5
hEWj6/hUre/oTkB5xDkYpmrn5hC6cmAThknbeWf2Jv7I1hwROCP1LCZKgyFjC/yuTKX6j6tkDS3O
yvpLzgY8Qmsk6TxqThReE7gF9kVkWzezVDU2dQFi2BUrz9/k5bygaL/SqvnCl62dHfPBCGkZ7m1/
m2Ys70ER8DMrfgHnRlZCJEn2WESnqJHenZQ8ghp8wa5YGkVKrzMFAX84I+pZpUjyMUkLdNxnnsXJ
MlEhGDNk5HkClZzPgjRi3UVP1tU5RFxV5w6Jp8sXyIONprOFueMJy63uz9U3j7MF2dmJg3jbgHVY
W7la6ko0PSdyH5CA9tX2mq6DFW3E1KWDwi6RxHEToJJBkR3MiWCDakGxfdruS5mJmr6Wq4eO4E0N
s1ULAh1eN0LIU+OHIKNPR2lW/1B8CyO6wjyWpG1HIx22WeaeCWRApGERClsVC2SWcXyaRFdyaZET
W0Q/bpDx9dA4veq38mCImhuVPK1ZPX8eSP8naa/b29gPDxGD6ZxhyC2sty+dUJUWiW+/JhtzbJE8
/9rj68FHShKzAPcuOB4q2OgrM8m5pUcvX1D4nMPEN80Ly79mimfM2hQV0br8ujPXSFfkBP71jCdX
VIWrZhc0qe2KOj6c15gFtCO4fkJg3xgeEJYigxcSoVrmsLF3cFKaN0MQD5ituwVAUoo+r/67aFW9
ZuMvK5DYYCLF0696CyCgtNFtHgcRdBdND6dXdondJsiJhqenhXlJV3hWFAIQRh6F7zYfNrhI2GMd
mklkjH0QMrfork+XYBb4MCBAfOqHlp9y2w0Kr/xKJ3Xo8287/QQt8KR0Ks82JXGUi4RBdKyBtyJ4
c8O16dPP1dWR2DfEZAU2ouBuYpTFV6Sbdl5aBNUndnRtEiQd0UWZSyaRKNuHf2nnmYnY0nUoAU9r
xTyFJPKGtWBTntLwqmB96GbFK2BhXVMJ/GLE1ja1XO0Z8xXh39TaHgXLetmcUv8I0KojaErhXMq1
JfYUd7iV2XiaUmnyZx6vKpBIEOwPOf6xF58RdmmUnlGsLfca3ZVl/uE+JNtTIaDJuj/xQGXH9roF
lKr+nthnKNPz+e7+TBzFnr2E/DYb3XrOvd4syyPyjS/FFQGy16n+QaA2Q5U/1b4lGPVVVRDphDTL
g0LrlaqJ/yThQN3Glxp8496XDyw2jNHtwsbaXl0+lkZ6ycpkjiAf+OE6rC2wKQq7u5fjz/0fe3F3
BnUhW5z4GfoiyuSDqi61uvFylRf58SjPusOe/SZwuDdR5+dpn4Q7LFVRoqVM/JOE6dqa9qWGXnrQ
C+ujxAUq4WRh3KHRvs/g3gZN8f2+1oy7nMVIvZhtBsWKYGjq6zZDBLzI2FfLrmuqK34Pn/ag+YHK
eQH8Lt3FDaG9jlPr/lU5hZLHAAMdmrPEWnFkcIB6srz7+wo7tB+ZxdcgImyo4d1C/74z13noxNko
70Tn4ckUntQPxR1XuQULiRdtSD5e8a9VRz0ITysBDonYPWAk64oon/Efm6OudtrE6aUmh8VPjmgL
r8GFBM4YpQ/9PsbL/jxuL2x0vgWEbpdaq+C5yRjZJCx1yXOv5Ko5gBkRamN4WPSdxnAb+2QVUHn7
P6hEgM1yGE1Fn6HP3/t857L7IsJ6I0eRuuqE7qOFv4DMKc+WHEJcEe4Qun0q83DPxcRDP7PJMQVH
kpzFTL+QDFczvosjfX20rCU9AVQyzembFhuan1glaHZH+cwQkt82dXOhp0N8MmyQ31O6Hz7Ijnd2
rez2v7dgAWItkJ+ACD0br1sEKgcSoA6Hc+pVKF8ROoIgy/XxHGaAcfeAkVyDpYhEbT1WNpcahcSq
AE5cQHLwyBkofIQL8e7HEsoxG+b7a7tBhLZj+M1sMw1dHWWsBCsLqOwdw8VnUc/m6jR3qb1ArFpH
V0AAsTCkiPq/hUMfaWua0BlRm+UoixA1K/4nepmRmVn+BA9XiYIPTbuW/tLhcQNxHAAdJyW/4riJ
32Ajky+X++mQqv0oWLF4GEliATDYecS3rQll4gvFwJNM9vdPM1KrHR/tNKM7i6E7yH/8kQ1XAJzS
JO9hG2FyA7yGu3qFS3nht5TPNZZ+bTuuA6l+O9ndjZLgpKN3RKtQWb3FpNrF5xIx/TpEeyComh35
Qm5FQs/YvS9/LOlzKgXaQ5vzhWs/ccH4pfpba7CqINNkI3PM9wLFbHVio+TpQvYZs5h83kc/Tvtk
LYnE2VNHcnfb4qhvew4TSAuCD5vRzNVLqmUfEhzybSHIfnh42c81OgOY7pPTuthV5AqlIr0bJqzR
aF2DpNtfcg5ZsHVmMs2dWJrfnf4Ywk3tK7vOGH7too2sDZn3kwtWg3hErjeNGaGFS9v5uzKENzqu
jdfGsLsPrbduj+K1x4Fx8n+10f6Kkwis4LNYcccXG6p/zrwFrVom2KY3D8lsjtRhQJy4Ae/WMODW
VuhbNkDlGcJ0FF2sjbLIzl3GauSLJFxDux1fMBBCTSqnxkBQUvhvub/+WU0r32nSgZGMPCch9J1i
ivjUxnomJ1BsjhFYF0bYCr3shfcQwnyjJm/g8owTRqu9fRMtudM1mgApe64ITL5of7GbJFY+3z2Y
eIeWA3ktPPa3WTUS4LS+jIKkUOYg/45WOPTdfIAtTVIW/Ya+IIfT8S7gycZFsSWZdekGRNuC6f4+
K0g8E1wam/iNeF7dHO1DU7hBie0T5xV3iTaJWqAvCZffl/xCJBgKJ7ZBXby+1tbAiz3yoWkc/L/M
/zGYKfeGAmzY6A+VM76VX1JkX7MTI6ybMdF6ia/bKr6zV9b4Mm5VNhDBQwdf81vr+FdVl9NiI3VT
FZ3141mUgMzhZIZViMK6WO0AGVnh9EP9PmKCugSJoDB3CNEWiee6y5dB3aNrcJlgCBOU9JFV+6Av
WD/TuDi/ht09rs2BZOL+wlZ52z5urZ8idhuBC80wrNUjfOyzOOwcrWCja4UaMURHt1Sduk4zdA3I
Jio4SNtqfQ3YDNHHE1EjP0g7ECvTEhKNgaC6hoEZWPQy3bpvzUjM0ol7eBfq1WHkUySmKLQkKmo1
2mkFrx+qmyY8MYvTvToWLhxF54SglKAdll1HplOSCoptOad8fAUj78PT5kYmAKJEhrR8+amDtVTs
xFnbxPhaKSTfJu8xPeDshApsFs0BAK4xpqppLfdxl4E/CspYtBzvZGv9rzLHtMIJUiKscsJK6OJt
KMF1gO99BMpaLsf1nwqshAMBBgnijDkIoeUfj4ZPwJbW1UXTwBTg34KLeeiilFPJHaDmk+w6l8Tx
cdYKURSs8ntSHAj0S3MG5fRW+2QBPQRB/arkVbcgOZPKnm+xUJxPLHyLJbRB4epALpKiHcqvEdjt
n6/6LTkScYqpBOoa0xslXSR+7HZ/8Nyq0dLbIvJ8rOGwJRQLcpXDbM3FJkTfJNL5Q48R9DLZNQDO
fHcww1nlv5PvASSy4GZ76LW3FaQBPVRFQ9QidEMO/HoDdGUCwf3lrK69/49Grq06h0KX/yNQyJut
8zJNTYztpinTEyN/MJeUhA76J8/O5RmEWmUSp9H6E3ni4oWg1CczKj9uxEMK+cxmDMhn9tkFii7Y
i/S53qYIoTuSv8m67q9mWMSVW1FCXpQOViMa+iTBSFqYNnot99321MmNu6XvwoG5zh/GhbK1rwbl
AIWN1UdjYk1GWE1n3YUce2QgJw3NJAF+ifUI+sIS6GEpoa/8v5BGek9VsWTj1xVbSE8JsSGNVvVO
AI74Q4uw10nj1/oL+oF1MoUPLxc4vxd0FbYq9N6Ymfj9lzC8/NGNE0SRWXfVfpkY8BmJ7KCU7MUs
BvGUeMJz48VY0cvhnlPqvbA3Dsk+dqlwhQxGJoXyA7CldtiVBtVeDUNfGFY0SH5GTGhfQGj/GKCT
9CeEAcmxWMIlWtEAOkKOGQ9H8VUrt2HyH8Pmjcb9nTEo1O01nuAYq8HQVyligaYnEtsqUJWTlZtE
9eEhrBsRrShl0us30L9UmptY/fbwkL2uJY4YG8wuC4Ui2oZFqxi12XzlCaGIWQW2XcA4HIQD1xnh
DCmZ4z3AP8qQ5yjHA8yaBXKTI4OUoQSVpG/kTFZ+1tgVPr0PebFNIKmwFLD88Ms2J2YM71MdbpN+
FZCXor5dYfO4olE9Fm3uBCio8VebII5FImv0dSHdmXoj9dbAIiilnPp3o9EHXARGfmgFyQXwy/oq
YUfh4XYJRDAyXbWUk2Q8n7ClzgWfW0MZ5pVAQaotebHKonC5HNzYBBYENy4s+5A8i0h2RQgq6rKg
mbsR9j6rRXUh/GF91xxgC4Pjv/nUffw8agZT2kJZb3bQAkk/DiTA5lSZCtj+Ee/EcXETzS55rmjM
lIoJP6TTFc8MKfbTNT0BDpIoLD32k584VKBi6niG4C6wv4csyDLbuECCCyNv1tbEG+Vm3IBottaA
8DnNfKGiXeXtaakirfqAQK0hhpVYYI4Vkpp8hLUX98zt74VIDhlIGyEi4cCQiAuEHdTRGUdTO6MR
KTLSSbut3k6sxS3U+DsIWz89cHDoJNzmGOS0F86fCOJO1fgh2q+bQGsfQ3ENTjk1rPV3k4TJEjWU
2Vx1uQnt4H7sQ7GPd7UTVAEBrM/IAdRgd8JouGa8p4XyyWJUpkSIPf7reNqqUKgO45U2nRA1jJLx
2NsMMNnQ1snWaFNIzXwjPJL605Z52aEXqvV95xtxA6TWDmneswEiSPVsYLoN/+6apzBFgHpZSMPJ
abzroFcsWsh2KWrFhLAa2C6K7xeUccOMXLJzKiNxOvCKetzTsW4iagj8kovQIElAXPn8oJ0jOdg4
LPnhNGpY15Ee/Zi0Plo5npeXAJzEwnHRnTII3ex8ZCX59kz4nipwCr4LPdJi5IUyWhxYG7za2v8u
LAW7FLH9AmEtO+QEv8nQmID34JwH158LJJRRmE+Jyr/HwoMIr1Np8V/DZ2Y62iZ/GW3Sei8qNhKi
oLhYvI0PRjxqqEKZyQH0oqC2G98lxCc31nHDu4PUMFSGvrCuqeXlG54bO6MQ98ToTQmGIroW97wu
ADPVKEq28DuZib1i2CE9+SCJutSNgbYXWXowLKYDJghpC9Ikv/f4+W97AHLueujvrGKX5pV/I+E+
5HOAAHwEJd2WaQyzb3dL6Yim0teMH+FCaR0Se6vabnGG5hw8IcNsmRgO3ylX1hfpei/KsXyyuHPp
EOh5LMT5L3VWJrcjS8zAHx32ep5EaKqL4BnRLXvhxMR6BtynXDdJXzdb3bz9xUrYhHVdw4zQ/nkd
bi0P+fLXggMr7WWb3hg2cnlnIrPvZF/Clsit639L3OzOv43lJ7R4bK9VHo9AlFSqAuEPVW7YVG70
k41+IuSzW4+TUjpE1SKzFfEkRmaCPPmz1sEdBnuBWOrUlTJ/jwaT1qx7E4zBgNGFIsRIn1dan+jk
IkczQ8jIez1wV5xyPZFh/LB5OU+uDOATXnC3CQ8aisznjRTWck++G7kGX99YcKhsAA6NVFFazefh
3gxOjFeFxJ6LHEgNcy+l0tQwl+xsp0FticZa8iGzQDqriDki7cFGMGEszfk1UV1E5Shulje5tafZ
+YKm5NLc8jVd8IIS7V8CkMESMZxd5liIrqmDLoWmAg3CmAll6xTX1WSc+m0ATWZcT138BCxTbhp+
cy70xfnjT8j2BJQZCqpCDfyubuuaPV3eaWLz7u4WvVVnml1YQAqhNF5i1S/+W1xADA+V5oijnpzm
dF+He+hEeVwgnsUss+x04BxppQD8sTB3vtu6DTy8pxME8Xq9OdSR7Xb5iZpWWGIJRjOOstk6/Fdx
nstu3aRw09B938SZL1nYP1a6ly87BJjvFM+PxZVKv8BodGdrwdS1aWR2akAHdF1q/lX14gc1xzOo
fbkUC3nZSRMm188Ikqfu5H0gb1nyDcyhIEu3VVqXZqCsV9yRlRg1IgoBnOyFNDyACUyO/krk6WHh
Ntv20nFk498dwAMYe4xhtK5O0iM4b60EA969WKu5mfMkIvaiUqXRt6k6RJay85sDFl43jJmiaXjU
SJR4542xLSpcPYwBrKuMcu0riNaasDv9x+yEUaJETOaUjC+2njJJUsPSJ74w2x/m7XJnyDXVZbbU
XNiCuJX55KU/expdpcfjKZmttgB3URwF4ncydD6GscK7ZKKgTBkgZFgbWYnmClw/PsKHvkAk3ITK
kqVpzvKHjO92TTv4X4UIXMF0rqLYOs2/8UoVSwNVk89gXEKCzM1PmGRaDQ5L6i1ubJItRzV5qc3H
U3w71DMt9xUS8F2sB+JdM2ugRnOOUKyPBndfhFPK3QM0r/7haFmVqfHL/qITyEvj5nPc5JUddmK9
hvfgJ+fvdKmai3Tn9OKu0d+DgxEayVejYqo9GcVCv/ucbuK/ocuHLjpzyUVpCeGqRALROqo3nCic
ZPHTvqxDRD0lcclv5z+OUUQ3GI04CMqCL3d4ULpF/lQeYwKrbWAd0d+tVgnbXry0uXxm4oLZYUVq
QUtG7/igoEXix81fnCqcklQGfI+OdhCKNV02XtKGj5pSMNZLYVW8G9LnC/PBQ77kzWAIgih/rjtb
zIdWTjJqKm634madygjJuTCDlr+AfTtLBLMVCbcMym/514vZY732H5mu8R4PR4NmqpJOBZ7ymmSh
CFmvCNuCSpfsg/Fz37TsNWnRI1d9gXWDwHrfKh5untNX8XWTtpZvZB3XSLmL8pEYUrpy5L3bjdxI
vRh5LdO3PDyABUh3Abb2G5d6rG1+QDoGnRK3aVBpFIj+hEIxskEHXi+QuPlV2BBZypWSD47joyRP
1joKHV7Zt0xVdNBor65liYQEDOgcnGV6hVO1rJ1Xp0OrPLBB5WcXFW7/X+plwKsilQZxpKn17qk4
fiZ2o7Ne45lmxdPZfyB2z7kgSBSEcG8xmyjsVfazwmp7H9q+h2B+ryF12KPSXqds8moU/ydNBLFb
VAEcMGNvSkiyxddIaoJtqKqxI6f8amx+i5NKpvY7UTdlWUNT8/my1hgKwNUQ9gpL+HYQdtVxSAIM
kIukAFCdI0rGRl1GwlS2bR5RsCwbjmuy8rl854gO5448BfKoWg3l9eRXUeLfUhkwJBi/lzk/zXuH
mCbfGymu/51BRWfUNfeCQ6l8+RnMtr44i9HbHEg1TUU63GXvmROpHAeF8wQcV5pvl+cpAJjhdWwR
WcqwKk7TztkIZklHF4zzcuvKY0bpyEk7d1fGqM6Qy5n/mdcGAPZvM4Jfh7K6ElOvSAuv7dXDMtYp
W2RQnpPTqR4VWnB4qn3L7GkEs9atAZwX9jnB0Hm+aGipRcBT6+bMJuGvZd9WsovY7pLTOfU1ir1M
ptL4N+aU756ViXnQO4OKVR27l+tLqi4AU2pp0WRUIAiB+LOEvseKdqbVWbBT1kxNhOjI6lY+12YX
6t9gDuyb8SnQ21Oz6sejQt6IYXJTxx+r8G0fE3lbZ5xQAdOytJzp25Vo1wdACOwR8UvKeyTpGP7k
S9ehnl0kMfCmSzDEXn0G12Ja/dkId23VNilrOXzEpfI13fd/opFlOAZQhZPHPml8dWLrgjmi2dNY
qDYrYr36qbNzCofiYpTdvcbba1JgS4XI+BxeGcTtHA89aqKjgp75C+q4GHrzS0iyOO5nhHkYOjC/
MnLBX/Yc9a73A2SmW0iAu8hGY1FtfxfCCdSwZfaDzcrf8MaJDJPrTj9uO2jYUhis8FyMXGoFP8yg
cx6qYvjU1t04w46IJ5h6KgmNbkSgtnZldKu0IKBkzAytG4+l9BCiUZLKetXcgKC5b2qcHzrMFU7m
oPJrF1DZRMFR7/xg+z/KVPIzG+xIlBwffTfB42AhZBSM2TxNmO8uravmMzej1xODyiXyN+6ZfLfv
cbEMZpd/0neC4Rh9K6RAfPG+UhMucciKnWQTOqJcrSIipB0wZ9GkF0uPD9wWLGnCBarDWulI0JOc
FOw2SX7TsTV0Po+GPYmxjthy78gtUr7+hMZqPgbrgRGHODGmR7gr98JOspSxU8Nf9yT+kWC3O/lp
EcKXw7DUtat3ZE2BA2r4672PYZfeB7Ml0AWWSyIq0b0KkC3lNm3/muCVCWRz1EY7907P5mjIPeEH
FZGsZJR5qww2qfeBUDYq+PF7wzhiOEy8n/H2Eo0EQJ8mDxlONWOmV4SEk0dBSF1v9sz82vF/EETO
l/ZJ0XDUmy8Xj7cBu8OWU2BnhAye3bzQxGw9dDyKusfIee+C/ZLhdp30sBvveKisdvX25nDmSZWY
LXXz7d8mMg63ktq4XU7tOM+WPxIeQwNTURyWvUcco1g/LHhgOyivFr9TtI7aRHeUsTE3vd8IHsEk
p2A42aeXGzpRBD8++HdJt/gHuCchXtwA7zVO3Bp9RiPqk09zxu6u7QfSGARuJkOE3jWdeoPftxHj
BbZinh4Oztf1eXtrQcdvY74S601xIaI14WN9Ap142m5mNIJQzoTRz8GIRTsOdqi1K6mQ9OvlZL8U
VP6sj4C/kQnaQ5DOvt6Kbbe3Jennh33KAB0z18TXMGWjG27k9w3foCChf0S2brnvl3UpcXPGZ28Q
K3NJJgqUo5hruaQQL0Aw1jO2Lti4uRvMGDmvuHhBaYa0gu5Gy+ThloRJLAOveAUtbyjuZU/TvwOx
XGSAsZ6YvQ4D84li3CL9ommSCmYuJPiefBpZufAj0vH2lXebq07/cx83cOw0kJprC9rq5uvMmLkP
bWRBKa2gfgoap7JhJaOLweTqeWp/qOO6y2eLcfMJIZ5YnL15JlPWGbH3yweXazh6ZetssZIqZ0Wh
++1giIC+m2oEKNdPPooKu3Cd3Bx4WGoRAmKfSXVZdFdDP9gdts6q5bXw8cPTK6p1GR70AaYY7XWM
yzeGqdA3B8WPKQPGC5j+SEBMXo2SyVUAOIL4HBWoFv7hssreqmpjsUoBPWuLK3/9MDswA43/Qbj3
InVs+GkVLUfeU+y4o4tuPsVSI4GIw9iGesEibTxNGvHvHrXdrZFLKidpVznU6Z6/RBMEMOurz7Jd
2KSWp18Wvc5Qo2JywszZZwVbbBmqN1ZhjbQk1cKnWIXizsYiw5KYs80mNfsDU6Vy6qqZ5pqnFqI7
3ZniOiFzvU4MayNKVaRO6DWypUC5DhCg+eFRv00hTYAZbl71RBGQgQA/nH7KansgmGfRLVeIgj7A
gEDauZZZBTZwIMBYWbI7gVZ4sTFD9+/B0XwLx22EeHKoXbH5l274aOkXa82lCm/+T71VQkzoOjE5
tp5klTpNyU/TtFB0v/eNTGjxqpC4wzIk9aKJNoKceVF+a+32Pepzl97OqTfDzsfwk2itXAHfabA8
gI3yoiSx+0G2pQNGzWMQUu7uonz6xd7YRkcXyYu7G5wm0df4mueUxhEGYN0QJ6pqkhV9KXNbFcIL
73HPIueN9SbHTzQXu8G7lsu9hp9OSI1iZApU6SUcGNq+RBGbmrXTieSMexHSIs2LflENhBjvJl3g
aDPVAvs+opVcgmKWUUl4kU0OAz7gBRqYpmRVCbcSbjhRpwvc8+ItVioIHUCeDkTP6po6vpyA1xfN
sxCBYQA0LwnRGp3gwnhhdJaiFFu3VBr23fs5/wpp7sek+k+jv4SsmqDCeLbIwUCZqoW+U506FyGS
KXyBE8XmsVSHagx23PCf3HkEgKJieTfuo5p4dNoO4UmKt/gM3MC8mn9bzGsg35N07cU5n3pOMGrq
5WKI8uaU7Xy5YsIHgBZf3J8E5TAOpEGgwvfAeoTEggfv+eYVp5Bw9SJvdszRMzWOfztpZkfUXfQv
1SdOwVnT220ZKMcwg+eg/LceLCQtxYfQ/4LKbIXKeBVxyTe/Uf3V6o5Rb1mXRMpmz8LxRKDBkPy6
KO5q+sx8ZyM73uCGCPvOOha5Fm44UgAmYwge9L2dmUj9Qh4jLIEwW1qpVLdOLXXNO8uNJRkyp5Ip
xW6roql/+csAbhNTGNtMRxGk9U/zEfrnGzqisdz9UylGRDQvviDVHrkqvOnFhFON6Md/kZtpMHZX
tphDcQsZoHCvd1He69rEXB+iPNR6uknpbSVyoE9nAr3hPIsLnn+9MqBAlc7XPaZZEQHgVj4cxJAG
XfCy9OhEBfUHmIY65BPu1WueBNmUWPt8x5ZDRN4s50UKVWCdTifmFBoUe5jWg7/V6v2Xf8jEH3ds
ks0IQNM5ag5cEwByiupuch6/FkK4mK9BB7q7S3JMEKlmw87H0fiFBb8M2DS1YL6lXZSSL8hBxOWG
dJ29keFpuI0gH6Fxv+dCptOCDMSMKrBcVtGEwXt9aW4MAhsY+CvUYd7Ep/Tb5vRYUtt0JBtE/Cwo
r8PgEQAFOx/Lq48LoRm6uRvoBXd3duDh6Nb3XuvzCM6H29x+KfT9iyptYA1N7QcopYXtmXsnosB2
3HNcUo1cR1D4y3ike7VIx9GAXFKfzBB87yJqAzw3Dsz3qVSzGRt999Z2MlFNH1sHE0eKt9ELF+4A
ywIvIvTaBL82IXgkfHSbZXIakmiqqGTmcnRHm8XN4if5zoHnx58AWnRwLLSP6aRJCC0j9xF9TRA9
zMu/Ii+R6ErO+XVvQe8Mcofw7U/XVigwkn9n20UBcy5rQeKcYS1lAfPaMqawMvZph3jI3RlZteWS
nSLOS76G8kYXvr4n2N3p45hajYwaYzwdOZN5EG6RGIZtNobTxjlm6NUxTVrFo07ufZs638IqMeB1
aoek+1/IFZVicxwW7rl1iBaJ48awZba0JKmUEQsRtnQfxAlaaXE0JSqSjajW6F0tisJPUmBMg/O+
DwRnoCkL6gcRUM2yAPbqzHRCxABiAn46QNmhFFf33JcdcPo9b4nMkpOh8GoUU0VbLw96eySr96kQ
HOXCaUQ+bYKu+wpFm8EOGTPjBS8yFTqRWKRnflsahLbrjhu5nipXmqHy6pSV7NtwhCcOEvFX3OwJ
g+JQf1hTrauT4h46NqUcTVPJ1brWvT/jiN5zBuqwdFXaur+W9/QrdP9I8oUAmEvBk3Bmqb+N9SgZ
n3yu7XnLvxrGXwFbvuMseYHbCaunXi7j+tU1epwgCfd2mwg/0ewHkvNd5aB+TEy7QpjNbBjHCtVE
wVU8oDX2qnUEx7uLvfZChQ6aGu1Wjjx6/4LvW0OYXr3nghTOTWdMZp1yJa4LYLMnD0WyEBrkHw32
8Ea7jtjBzv8OwriuHqE1uBcvxBZDdCydD+VCpEyi/DtermQro9+SIl3nnkUpnueuNK7zuQ59RnzD
zrRw8iPJq0VZofMa4yxJfNO+nONlD9oRFvNbGmfZFd64wa4Nk0dEoW+NIQ2lA+GFk+JmTtIM45Vb
tMM5B0GFjQ+9ePdkECx4FPzY4TwljpQ68ZZD6VKQuzcsxF/Rxw+9hDRUz2SDnyUp3HlNQ1izqAyl
I0/OROeKsxyJeTnYOff/5f/zMxGIMgVznBdR0IRMGg1kC4D93r6nPpr28JrIJHU4BcSOrzrbFECb
Pwua/aT5SbtKwpZ5QUuFzwtFoZtF7KJ8mrjY3IxVM71E1jfR9RrSf7tIEByuU3EQkXVI6WGyQ4mI
KHl8q2CF0hXzUvYQJ7G6tp3zLiOeRY2FtWDebqZfwdWH6OMYNosqrJnLjaGenMgOAFSZThOHqXmS
xvjEYlSIk7p3wkFMU8QNap67gzOFIoXIMi+mgAUxgscVtmKPashaodYGBte9l415b6v/K0hRue6r
ynpkHCo7U/d+y3mQAvqnW/L6Omka+ZW6Pip/DPuTBm3+e80VB4VVTFI7RUaWMO1wn2IT80di69J9
OflVG83PiplPT075MYAZRi0H9ILq+l8S1GkxXud36dKzmAUDDFQGK99OHT+EJzPp+3Sj+ngDFm1E
7ON7cDo8zeFGPuznU4ZzieF7xR+kB2nf1q9GE9v7BaRfUg1n/WbKQGFr2L0TBS973v1lqqjP1a3m
0AeHtYN4DXPgwY/ElPvdU0RFS3FdO/t6NNcOQjpLDVlJQ+C0mtE+0x3SDszUkNag99lUs55BODKs
Ehk8o4inkhyq1/t89ng6lTU8Bi1u5GbjHb8OeEG4jZunlJ51KCkZJg6RIFSnbKhiYoXkWlFrp5pN
1ES7ab3Wo8oZlqTKRuBJPC9Lg9GWKf7PrjODPF5qZNW/C36g1o5/3M50YKx6EfVFqlVydcx6lv6y
5CPwbJjeuAjZ31pmhucwPtcAwtr2OhdZ1DkYWI/JD5p+CN8uAhL3ZkaKr2GGQ4dFvyiC5R9bcYbz
CZY4i7pcnQaB8+8OzuwrFxL6SSPeanQbT+AqwAD+0p4V0CNFJoVLyhj+X0g7y4yEaeKLCh6kU7p+
zTN4DfyDLv9g3lFolzKWy32IB+WZqz4a4zaZ/fnl29HFeLhMdatAOi2kmoabmnI/q11kfWhtUsVE
PkZ6ywqftnJ5CRYwxfA0mCsp0HrdFr8GcIqrDj3JzWh/8UQVWEoGoLrpxmvsphdQyjfrgVlyKJH0
jcTgVDRlnLuS9Wlaz2jl7qFSHxd+dx0jVuVbGI8DDYczSuy6B9Y3UYbruVs9OlKJlNI6OY0xzo5H
AUnLNnbwvd1F2ZK8zgzUgV++b/asswHTyNvAru9ToX8nQvDtsp8RJOAK57GIi7pv1kpaJOebvx9E
UB4vEsoXBJFzV6vdTzAvsjzhXLBLgIGEYthIto61ufRVIuzAH8PSsQbi2Yw/MchtasYhSZYeBNHn
EOVNptDs/+j5Wzu09O8Ykok9jfns2V3daaDhUXcV+6DHM3k12nTMYb/MJm4e6mSfKedRCd1ST09X
XwaTxBytu2AyfmMzdVuPeRW+t6q08JxJ0Ur1A9BTnrtbamkqyDJR2CEKq4ZhJDnQz2lEG8zoSPbg
9skyjObVU1ld//izRZ13SHRtEewUi5wmbZuf/sDFGrkmmx5IPURXcgpskKS0LxBiX9fezdPQevgE
WyccfGle3fPE030rJ4QvHGE+ZnUsGd0HRqPBwBuDLnDwolNNJUPnhhNyWQc8g3xlxjDHTfP8BoGi
q28O7L3LnmKb+Y35WAsbzMkrjiPT1Ay4p+1fng+Oxgr/+UeUfsP4e0Eq6NvS6psyrARAwmUaGyJf
Xee+SZlnRLFWGV8ViH9EyFmeTG2jbuRIWMG0z7zazMClC529jyK+nRmRKBnv0tPPizT3w87wRXKE
Iwg+BR38a4dUZDIfxwZKRF+xyslNYjh7saX8P22fzx2yBn11ilwvjsDRHDeOSLLjik7TZ2rTtnPF
LHcQWUo4LJ/hMHyFamYvQ6u/1wNrqi9fdEprXZlkJyhLplobUVF2TaNe1ZD4APzh8Jcr8U6jkS/5
Yz3Bms2HuuKF0TOXtiKMuPwCTAE3oTgdVzgDmMAL1sQLzKmmo8eKwKAmVfDdV0aPUnmDXneXG7sY
kNwfYUZT/Eh70eDWLXFhN1qWt/jGdy2P3dtQVOgMOrIsPKFp090PqNlXzFvkdsRhzH5KDUeLkg4k
RKzlVLGdlVtoIFLY4w01XzyMToYxfg/ED3+MoSg67Q54GL1GL/orGYKUL6gVnjlAobcAFhblOZXN
d3IgD2Z2yFW4YGpd+KEG7OIyFIp1u6NqLJolPJSh/YPDVF7vi8Skke+7XrHstv5p8gmF9Jyz/XN7
qOwFjQdhuKONadkYpUOytx+LADmrPvqhs2pWr0VsvVGgHBjYBcFyydDgs/vA6oyOiwGobyNpExys
AfLZOZ97/KsV3zoCI3rkNkzaxIYDMxBXLdtAXy2ABcbf3GleKXe/KiGx4aCziANBAU9mtYBTU8Hr
uOciB4C17VF+wvjfbbk+pNb0XfzLSY0IBRixb8jEyGET918VPPHReyj17VM6xFcXetsDmqS+SCbf
2CYliGsCjDijBW89Vgl8InKNDn8H80iILayoeKHE81jOgV57ZrFo72ZKbE0bT5bq7y0wntr83azw
st9bJOAtihgclcObycg6lj5PzxfRyr81LgP5lmud03yBkDTFpNQUxPUcQUZkF3APWIzwFubMI1E2
PjKvbGchLGwm1xNcw4pYyNZngdrDMYto9993FDc+aQtk3q3lh+RZyK5NqDxeB4JryR7pJxqXD/fo
gtnWdqllhWJeEMImCG18bGZWoo5whD2RRuJCzuOLfb6wLjH37sbdoS1bph1Kx5LhP0kNQVc9VGPw
y+Vx9jSNYhVGtK6zDWdb8DK/S4Y2+QmkFlgZGr1KLppWZRDmhtvfR1uZCl1UVEaphVAATYLbF9jS
tyFomhM21Nghms/L+y9r/YmSO74QaFSdg0bVItsYZe7eF5oi2gvUhqRJYN7U0fkG9M0cSVzaS7iw
ZF8iYfQBLiZR243IwkOohQjwkMRD0848ls4uf2U7OeexJV9t4G/WXHCC7Nh8LOVNqWWXEtz15YTM
vFpTRpN9ZAnct4PZmvO/KwjN2FB//BZzjgIw6JQuQ90/O6Xp3Cw7cJdZxGRoxs4dKTz8Iz98aDxz
gJkyXFt6O3TnuoT7QE4iU9QvU9PlMbmw8jW2ULLtYU2YfjBgzqsIHC6+3MbZDTgyhTENucAIIX7I
euYq4hybF1P/ea4azv+/lacWsxtDGzywjZWLVhAXMLR6dqI/b9DNeazZ8fnEZ+TTlB8s40OB78xp
mQZEWh4GpIOtN5W57XZAc2gIN/L0Ab14MnVOfdhAqNiHkvyosxbKqeYuSmqbq5WbGqg9ETXqRNi2
PSAuhakyooZwRd9jSvGqp28XF4O9GUWzQ+Bpm+TWXrMsflqvJweSmyrk/Ya6BAnFHGsN6fcb+f0h
lNlo43XTll2cilsFaFESRChI6Uj925mihvlEHFgGDvrkRiq0xjpoMOwzxog15JKCObTdEudw5ERV
mqI0X/y482QuTetReY1Ml3T/Pny5G50otkjq6lSQC47cy/mLOmutGH7+PBJHJGIgLK29XBUJun90
RB8weFhh3oEM99Hc0qLIshW+dX652G+E8OJTUK7IXEUyY16hYwniX+6jC1gjpPTc1uOjtsIOg7bt
jqFUTTjCFyhhuUXdd5rNC/CC8GIN2f7OMg1+l7WQecV0mBkThLjAmgcDTXqezK8P7O+ThhrkWvYq
jIa033jHv84CRMstMd/VUYugru5Jv1H4TLQUrXV8elAXUy00njo0gxejlbF5SZD1FazOLs4PR2v9
KkG5ts1q0fRuxxY2eO7cWfAUJ3GNUK1lJj+BVVlJbr3IHwUkWsJfsXfn/4f1NGEXN1MbVZLkOqCg
5N3kIMfJkWmA2GD/rYHApgPjVfQnzHGhRWH3D8koeZcRxO+LjkzdbGsFUYNxQ5H35qq5cBibVGMR
Cz7YDxClumuDMbA08ELVc1thAj9y2I6iGubkcz1GNSOnasCWz9chH/xJI5cvBu8wJBNsEqQI2xWD
6d3to5wcGQAsmvbuWE7jr/ZTE6VXnbg1yjV7mtKD/1916hF4cFsDMJpnTgOfG9hqi4novN65WtK3
zpgQPEF2abE5DLL4iN9W3QfzE7zhRlqvTWvlRmbcg/5aaD1L+uDC7vMoeoo0Ml+A34FWCcV52iDH
aVNcSt9Y73C10/rW5qSg7AVYov0DPyhpUBTSpGDy5VYepTUa+arj6xJt0nQi5l1DAvvYfmrVtDJi
a2+Dh2drAnvk4C3CYHusOZWwejs7A6FkdxVWydcyal0YLKoG6caH2esxGKJUDmi8zVy0+PdJjuF7
LYEK3HxA8vQrT3LYBXq+dG6p3JG6p1UQr1nZFq/IPAgn1lP92oPtq24+4cnpk8Wr9gRwtFxaRflg
0FgKUhOKfAL5e4jsHCly1eYGXiMHGp7a8iioT82cw+ZQTtAHVXZWctw7JKd9DuAV7eDInAz+B3Fv
BudBWq/ywDow7sWxwE86MXlIqaxn5Zb17L4ayvVcolub54f9COj+Ftz1wfSjELUWs+u/U9g5atJ9
RLso3lSqhuZHeMkPWFjIehGo4BBmNSekYP0+eq2W7eGET3oh5Ea5CHZiTm5ZCqUUG9cdGenPHn5g
EJWvbFiSnI3bjuYbOlDXrwNQqk7jNgZ4Bhefd6QJFB0KsH+m4mMwNb1BvmCx3GMDW3SeoGyOQxTF
BxqHlELtUNcryBamw3Gi/AlplZaxeWJaisN7k/qN4VxDV3QLg/PdUgcBJBLrY8VHHd435AZ8A7L/
WXiKcxBZUCEpu7/V3hqZyFFjF7V0Sajyd6Hg0tt8ZtZlUAwunn9AfQ85ZpQQfZXUWz+HNF8ItQKk
K8VK4yxx/fvcdkqtwVqSEiBGvkAg8WLaFWjnKIcR4PFA6EIrCVUPxJjT1mIcleU48p0KxFFoyuLN
7Z3er3a7emGkSDhty4887IEpCF+TL1NrKASrXUhf7kl5mhDiLmfTEUwm2Ao6wlU2tJOH5/BsreAF
oo75M1e3SZscKtdX3yWCsVwc1iGRQ8MJXmQBQQNI51IRChuz4hQdnGmimw9BzmsgDocnBBflxAzc
a84UzG9MN2Qf30DlRc9JopWpEEFx6id2aYzj2wEfMmjGVX/MXkywpJ7VXFvf7zqBGeyuvpbT1+ey
UxBNSjI6e6JfZYzBCg8niOse1fUTZAoLnUb3zgQCQAXpHceXK6RHAx0UK1di1BQB9gpdw5k+hpHX
nO77S/DPNKpO8lqBqkn2YUDGUtCVLqlMwZYhGxva1HUsq6IeQBUW776ucYg2tJGn+y8o3B9F6RDI
+BzxBo2EiXOdT9Q8KAqgiRUCHg0fZpuCI5ViThD8wkvaAnibWofcOfvxXu/WJmBvsgDD0VEOl0Hm
OlqG5mw2iD7w6MYJ8CLth3hWCmBgsU4pq1WpjWDsZVTUBZVM3amW6f2S4hRZqz8Tdq63WZw8hcLG
p/NcoYkAQusfm3Xen450il8nCt4DvHeaJxPnU4d8TAqmS5mTv5DKSXuUY3ctyMKvg2L84bImOsj8
rDkdAijCZk70AsCEgvDGsz2+X6sea+vTSsLWaylB3A5qfFoyocg/VdXz/qtSlHlbX9D6XgZ2TyOR
ek/5UDeA1gU84jiJtOAN2t2p0rwbKEE/Lgv9d1J1Csit7fJAlgyMdUS1QldeJn2MdnyUTBhJrN/C
NjZl1AgnUUy0d/kxdTUWNIbUUETq3/eeWb+iDR0m914UmJxa0MIkafjVZjb+sJkl9MSDoLA4hE5B
+yp2sqYr6E268pNok6ydEikfI/QZsnwiyDHYIGUfKEHqk9vP25voz2rje/Gpo4f/bUbRYrICr+G/
temPVpxpQC6ABKKDvUZY3vtMf1cCJV4GjDkEVOox4pTfSrqVJgaTUaQmy+NkDRGT6mn9fcbkaMSV
rqI7ccdS/t86zP786EXCa9Y3a0SmYnMT3RzlPr33/WqmjRHiUOmKLRWFvETWDXWAZt7LmJsAaYit
Z9bSdQxFlezejm9FfWPgFEoRps5iZcMWhunCrluGNSSbd3wac7sidbik4KTBLBPs3HAiCtLvcLm/
GoJRR562lLsDs169Hcimwawkh5gocGRSlTcglSyPPufg3lDR/DkcG3f4DYcx90a5syChe0xt30V5
bH1Rdcqz8lHZ+q0PGpDdLMMurUJxz1KGWR8ton0ZwNay7cI5Onvo7Xmynokz7Y3NF2EGWcJCiUTM
3bbZFkDFFECWxDGqLMmxcES1i2dPywSvDNqba1KSN6bDWOwpO9j+aJ4RpyYBPEji1jhFdsW0W5MR
ZMFCkQND5GJX/IsNpfzu7X8HPvaGMHI5G5myuuCKJTa0cJyYWNK0uBA4fV6q8yHBBPUFQwbBWrM7
tRsl7/wkhRhaPn9oXWE2bqSMVyaQdKi7WXfw9UlALySQjvv1cYzpLUgxTmq8xBdyNJjKYdpOw9El
6CPhWWDarDmMmhFkIhUUy3mXMVJV4BsuaJqTN9Rw04ts6vlgqC3EZu80Q/oqbjUNqHgYjUhQCYvm
SbSp29C1A+FdxKLFEZQdnrpU7Mv82ymwLTMS5WVWaZGkNCYNiQbBguYmKYQu9qz8lJOLMINc9TwR
kYBICvwdiO9ukHfNZT6qeUvwZ2f4ZFBgMQKfkWbhC+uFIsVkgwacuAS4RMmS7R+WubqaeobsazNV
I56rFqEIKi64abi+jR2q33jHXQv7WCwnDlPAEbrOBMHcYrI4LIGfbUoM6oVyoAbVu66lliboxDNe
6x4BS1oKtD+6cb8fVxFddFx9rNlYMxIAzaezQHnYa0lI1fh1lnYQszMAywW8jcQfqLkdsJo67yFF
1EAKnJw8Zx7+LD3wbPTz730X2uChiuZ9DlWKgw5b2MnI9jLY0ucmIPXbIVg/YeF3YQLmvdPMORXR
9dj3fp1TPILuPpZjQkVU8psTLsf0ChzpelUsOv0NMW2JpTwmNUWp4tLcVWi3USlzno7zlbzPMvtr
dmU4sVOppB2WHosKuv9ZjiJH4emZfw3OU5Ud/HZY0VMPJdL5R8EFo7T69yJ+/R9HpjU9z1MVC+2c
60FE7TrRl2IUIxr07hghzXKOqYYloyV9ESx+qKryXDzlS05JqrLYEijwtfz5GDAY4/7rE12qzMT1
KQEUluCLfeykHsE7+BMRSYbF1LTEMaqOSFvMYyIEFWPBUl8m6D3uHBeI51NVJMztSjb7/RH3SFOs
2GjjNy/jef/0yHXhiyxwW42q3VZPw9cF74XwbEY5nly2l0mgvrk6IoXctTsv60Lfnf9kb/439/RH
UGf+CvlrlvrrlmuOiKXMPNnlvNNDlnP0QFm25IVWcOuDBgW4k180U5sytEBy1MMbSYRAx8ZoWCEN
R6fCJYK9923sEYIKIOxLQeN4CvHibpj2M7hlVpX64KT7KFSJfQUm9p3XnKiuwoWe1MAT8izMmFn6
uUkIoyLodgf7eaAIKfSUHmbG5z2wX7fbOBpah44uVojkvAcqvOoGqYNuO896brChrKw0ejcEH2Uw
KeItfeiUVlbxGaiNoyjCRDXW3PLdl2MAkzXXJdIhpAW6ao4voWiakVxOCdjWODCoHAuGzkovAdhI
sKb/R6mafHBxtfuQS6yKELdvIlP0BInqWVCoMoTtX27Zu5cNSCrJAItrMqzZIBNB6IogyvRqHsbn
NcuOYQHO8MQwa1gwgk0O9uvk87nOI57vsLuMBcp4QvnJ39DhXL3sCnHBU6MxLnxNB20PZHFECkaM
4oWoFsm0h540QfWgF0gmJEQy1PPBvDgljHAG+K7P70NFNNqXCnx2a2yDirhOE9El0D2iXkDcGUC+
b3YWcuXtPzSLR62uZDNSv9rIjw3jkbNJmwytvGfQHz3UgrsltXUX8urlASGOysWSlF8TX+vBp+rF
1D48/zP+CxstA0DsUk4FXKQPmthH4JE7aWKZXKERk1JfDmjpa3zqVGPL5vOlv+W5ZoivUsN94e4l
c2yJ/1RJRpyim1Ap1Wnj0XjKUTG/niZzThyF0/+CfhG2V4L4axNiH6FQaa3LicXQ8ofQXhOZDV9X
Md93jm9ADTOluSVSJMQlWq26nSHZw6PPvS2UaiHYDyDdLNPOkViOeg24kDS08inDYXn8U2ayMgVE
6MRx82AW0V/39uzsqOQoZvBPR0ZVusbndmjre5bxeMZaDpVJQap/BQE9XbrSj1HdjQ3fWMasbLOe
4vIdQ2Vn4NplesonnIGP5GO0+/kPaRuoC5xLmqNPG5MybxiNjFUHU0oihG/ii2JJbX/pq14WKZM7
JbCRTdfpcD3Vn7nv+NOUY5Ij4Qhk72098LjAjF0nj2D7TmM8wRwksmcduVwj5daOf6uWnHR04GgK
sGfB2v8/wkVHa2bUrapvHb9y/qOnxaxzZB0enUnvaSI7ul3lStohO/Aa0qPiNb8diNLeaItO1Bvy
fWcTNlmym4WBmcSIXXEr7ouat58/OL6TGJZwR9m2ZGvL1y9HsCOwRllvVoU4O+8QC2VBoqVM6IGI
D3Jeakh5H67z05PoAqkhY0NYfov5phiwUAHBSgWlamanjfHutR+uBbORtBwKyICQsN0qkgowrxmF
TKYiqETi3kyTMqEUry1EwXzoBPWf21X3ESbYlOMaAfq0vNIn3moEaY8Bj7UKOD0cLYq+RyL2F6RX
WCPQmYSWd/BlHgHMEX5w6z64j1CckN7FI+/lzfnBqC5Ze2043ffOnBUbQgNjn8Dk0VM1VlUpOmr4
TyqACOCaeunr8UW12dvk/+QHvenDAy8SOshirzWrTmQP5gRKqh++4qejjYiVkbFTK/qoDekIc/tw
zzH6VFOaawcEpBsNLYmwnO9GbyAP5f8dPhXj6ziFAa+2svKYNjsi2hw6+8ocz2ou0px3FgKJerCe
txDvtEUPHK41cZgGBUZtmmD2U64gwbEA9EfbvDpUP2vCMPkF7JkjmMHiddfwyQFo+bIipYB0opq4
/kuPgK6K8s0aT6FY9xBuISRNlXIKyfVF05dPqAN0zvXfpSG3XEWEzgKCZ5ReYrdmeQzfyxeRI293
bK0H7MNwjV/AENFO6sHNfmcPNRp0O0Uu9COnDgT5vUrh56t5guvrdQFv5cQKF5w2N/xMAfcOMP34
zh/riE+v49Q0umPp0pkEkz18qUgH6Vj+BYTZAFOroXAdRoO7sGjks8ShhJc0j/AvxMvApIi5l9bb
EfC9IWp9X393xUxX5/kb61Vyi0x2qmyfN79VtUuQ3jXTXBkYfubpAGxC5vyszteKCbLHovdI+UU3
jVDhxQa6R6eSHpK4ClIpj7GwIk+z7T9fVYyh1cBH5gaLy7B45/iB5hrflfPsofGBqiVW22fIITfv
atzm96hAlJKLLD3ZUtvQi2FXukfj8R4I+q9i/OM4MHqYngt02IIzqVEN2Ra/CdPXWRPDss05Vx86
e3D3d6xg3h1ExoGlbQH+ul0uEA1TppvwCNcIavbFe3trl7+0DqbdrxHSX4+iz0/1iGQ8LuIiTrRQ
HCg+QvfKctmj+1i2n5oBTx0s5IT6+ai5ydgvGyL4K6OpOZytyYnh1sx812riEWOkO4kLe3J+lVZT
itc0XF0zeZ6DpDgLZgCamlV3SX13KfHZnCzq/XGE/0QL2MX7Ih6J4EiqZMLdiTXTRzqymOCKOyS4
REa2V2PsZ/GI/cUQx+hNH70ZnWF/yMazGB+fzsgGtN+ZyJG83UYZv1hC//70bb3LcTgavsyohQij
0ktCKwxQH4Hz24PBqxtASyB23D5adxeyGnuV6myHimpCOectXuAdRvsGvBzGpJ3Ag6X3VcdIkfGP
Au1RvKH1v9Xt2ISIWvOXU+3sHtepDU7xsOhpy+MaUp3T0v34N55+D8veS3PKJjadixnjHWEN3AY0
Vxr8KlPtnhXDunGQe1hhJ5IiT9KUjx9+11OA42jSdzjNbo+pZAX1pn4RpK61eqIAzAqGcc6eirKg
4CNUCYofKhDGe87Aiqvnvs0RrZGCgyxiV3kQc+fZ753JLPpGbVijwV7aqTrscLDOq7Dymxr9Y88e
l2rnMA7Rb1yWr1q+ewMsC+Qqy8bafD6U3TULlGuZtpR/TwA57wo6jPZD0o14Y6H1GxpNZPFXtScj
exZU05JUcgKrvDk+Rf1htiPImgacWxueAIRUAHY3HmEiORnZBFB0rkhOJF7k+ME7/aqdM449vkaq
2/pBAhy0mI8/Gr4iH+X1M4HgevXFl5MpEesomt4sG8avr98Veph9ltygNeFk/z2QjD0ed2gDh3Pg
uruRv5O7O7c11LkfcQ81ogo5eUkcLANRlN4pqhQ2dHCDwBDP+JMJazCR+dvJ1MWvl4djoZOQ6ZBo
uOBXvWbAEjAM2Ni7LhfvBOHKRyfb03HtxA8dnDaQW89yR3OLZ6cG40cw65lmSVjqTGtcvlpS22oC
IN2xasrN40BUOO8OoXeWmQRysd4iI0qR4kGeQSNN6az2kQlqbAtcosqEuMJMk4Nu6bwJCgfKrJqB
3tsmbhsDbEVIflJdRAr/7xV0BvpR0sp5C7q1yHfDCxYmJSsbOXZ9Dv+7TaEauS3yGVqqix6TufYY
PsaHusC+eEq0JW0GqUki7Af5USfU1oSe4SRnYpNxh4+mJsjz2ZNfShX+ouSj5GqoBY4p3vHau6V3
vhT+DwGFvpimzSE28aIE9Yv1haI2Z/i4w/5KOar1SNdBi8xNK8gdcl2stFY/J52liG063HSxd27j
zOpSl5nAdQFj6D4+09lTOtbt2Ho0nIHG+j4T6zp9uPtZtd3eKatnSSWAhdfPGLFCEN/VVZo7QSJq
+relzvaqJ9zfK03/Mu8ZW54jLPsgQxO7yV+DS3LeiMWw/HReni9hQOkCHe8WtZC3saR0isfQSQHe
JgPdu28d6v23FT8zAP8a8dHOz3djh7jbRRHlsnrKfQ9okQz+jlkaqqDiYx77oictWTxmkmJhRjrI
Z+casthpsLFmgHA+kViQqe32t7Us8o1x6dIpkoACqAI1mMrlTw7rgtDzD/Wmbr+/Hr9Onf+/is3P
RQHbwyeqehC1f3VxKUWiQennhB8XLNJfRn1wAqygOW0NOowOaWrclN3qE7t1UR4Xxo1lXEq2TRKb
1MQGk6NIXHzNHeOdj9RFC9ewGzVICx/wgHBCOmHSzQmK4GsGnrE0bWJ2H9WxuLw5XguWMulCeSzY
tQ7bfFm0/yXs1Z2/tTZdFEXoM53W1SYtKUPTnkCbCG45kvAyZ59TKoWQqLue8CqsSphU3JniHju9
U8rrGAEGmSzQRpMTs2N/xb1mRAPPPUFhaXGWP87zrn6gaIUK3Jc1Cqs6I3zi8FdEcJaMlb5yhHTl
qrJLu72rZByBgcpE0Oydf2xWbSIrk2OZkpkeN1M8IYM6azVe51DMY9ZcVnThuBPlDPxl3YRAJ4Y4
bEwmxV0N8fia1eAKKb48C9TZWJAV9iRtX0qV1ISkXVQVY1LCGFUEA2J+16WWjYUWOc+vIG0DlPyA
JGZkoedGA90qjiX486IZoLtoXZSxiOGiKCPoE/1wjJQlepeZhqnzZ1yvxOuTnhxz+rbsa6wfh+xU
MX5SywsQ9KMGxH1Vtwm8C3RnmDJCTwI6VCvMmfVt58RhtIzdvwzAlHR3pp/PxRI3Cex+bZF4UYo2
e10SQ/1CwsfsL+EOoPy7cfzI1s78URpCQeM7Pd+gCqycuu21m9KLHvugbYAf6WSgxsNPkwX6b44U
yWO1+E6wpJrxCUgpXGqNYegpgOmNLTI3jNrbsKZJEmElCaC0XtdnRNXBJ7eGyCB2l/yCWCylESTg
4Vl/ZDsrVsptdZFY3/RW09IRa0Y2EFrbjSgzUVVVw3F58p16bP5yU+eQgkjptb4j+p+8AFPe/WJU
y1bkWqjSLDyXxDf/yVsA7+GC4gZEEZMj7njbVRkahyeguCcH9Yg9ABjVc6T0oECtU8CbQFIoj2EA
qbkPQaUpoNIi7bZvLubgUKLrR9L5xHccFjM92pYtaCKOHPkt5U+sANFJ6fhCd+hJBvai6DbTTGbh
1HkifqMxKafkwIMPW6hWnFOLSALYJ/4mVvT1XPYpdYdms/j1wpM7cf6rGHxLX3NvwT7TZjwo/n0k
tLd/PrDHQmoieQmBCx9UWwQchZ2dDqbT52NrA3YFGOlEO0VBKBtyU4aeLcTL3m3xtpQ3H5pk8znm
+tJJ+e9hDMUofdjtmZiFMpxLfJfzx0vV5GLloOpkeqYT2NtZgIeNseULON4ajpURutLu4PdrA7jm
JG9Gnzx1TQg93m5zdOPxbbk1ZnzGtXKTiemyqD9PceMQu4jTMamDMfi4ROBKv5MiJZy1DOLnjz44
E0sbUJhoUvbkWa+kcExerj438Oh6kdJpT0qXn+k5Om3g0WOWccd60jWwebIOfT0uKVSNqO74Vocz
h8TzsY7yRDvuz7blqz4P+kaZnoMxU+S9hblC6gm8w/M013gWD9RUqD64oLG1h8uMpxqT1MSmpTBL
N3rPdWL4B6er8D6tqgHuqGHHRIpw1ls8On1E5e+1zMtmwc6c9UdhndXoinu/eAQGbB3d2DWZ6Op5
DCQV8ctRFba0SbRZyWyUHvZljjXpZU10Sx1FNKYhLcct04SQFH8nbnmiklV8J9d1jjGkaKsvkbAl
6ZnSD1TrO8Y+ACJ18b9dY3I4iKVXV2JVO7TCRMWqgbU7pxSiz63sHoxjUmIpDSMSJvmUexG+Nq69
lglQc0v0Sgn+KXyIL9cj6XEToPKXsGQZQEXICAH9zLuKFc6U4ms5LVo+xNDi6ZE/bSzqqC4gtQta
YDPm3HAjyThBZn5HSi8wOXo63UBw8OoKdW5U6rQ8ts9OPAJzOQaecRjyIkdrqBQq7yl450h7uYQj
FDtGFGIbhRYcFK8Wcgm1wJ28Dk7wqWORX/FXfiYmy4uJjBZc+ez3JsghHTmWjz0iEhOwVIX/yGw8
Jgs08CUMFf02aBu92dmXgt8KmHrWT0ZCy7JH8/7AeNXawuTtcWNnzyeO/FSAp/yXDFaA6x+v+eGN
G2yt0ebgNtqKQTtknCeA+/wk73dhH4qhveIq60Q/VVCqIhV5GjRpE5fjzIanG6NOfZ3ynEQhi2vG
JZTxxEIXiRnVBObPVHeiHqlbUatFGri0CcpDMup6+qJbhDOsy8rswNNWPGE9fdJm644nRUZkL5Ih
YykC+DsWSpLszz/vhT/doRkT9szMLfGJ06jqr04V3TvlwZY8IDdX+qK/LumlsTTFyZOeM2p9WOjn
xbhQSYz7NO4rpqcNCSrYSpUCOtZwnj+sdw81em/B/bTKKrqbw81E6bJ9qapOrmJbbdDjIuGtvoS/
nPkUXpe7vsgR8cweYzxZh/YsoXo4ln38kvxh5J+6QSXPaDW724tgRAsdY9da/Le/YCfnxJPq0sU3
bt4XmGKl7kYzLXc9nslF+4/yD5Lb//ivuRE/mwBtd1ro4653SozMZZJjXmyAtuP7V2YkC0shTWCo
GMs9Cc83g8PSo5IdcnSsX+56gDDqTp76bEIOsKNo6Hm4kf6OM0SZMRTVvLQo0fggTn3w5BAdYEdY
zG/Bp2UKhNaLS4DIIMfvUL10tuuB+sJVxe1/patkalcdBpdSw+CRh/LXJsiedawJCD5AxCFsImLb
dXTDjtYn6aYyXQsnTZSlX1/vQ6XqKSDnkEMOw0GBEg5eoOSe3qxTUnCh4+fPfMT7iNxCdWMq7HmG
blEF+wgjk2R/bDAyP0QpC9RIyBJZh4jMHqZEQAUxmmrmkoHSb/bDp2gxEfJda/1KyaOvUhRs6iN5
9ea4ben1lfPYrMrV8N5kIX5VmL7PRJMeIQajfbn3n08jEhDAl5mvMy1DH/O37Bu/Y4r3CWVzqB4E
NyH2lit+YUsPuTS8cAJ1sp4JmW6O44Z12uQbObaq6hVXVQ4PcgtYHBSRAubQ9s1bBhyyZdAWMd3B
4E94j8XMDns3cNhRBnP0dgAVp7dn9rhgMzHBkgEZrAovYAbN7qBDubsheO2WkOotZSLlVN2seWR4
1f0WlRCCi7kdpZLzvVRW4BN1GrPS2j1WyXUhTn0N+XwjIfe2U2KvdZq0L8PUhtBCfmCCi4rG1A0F
duS9qMRMPop/0CCQL1lMLLuhj8Q9dlPth9wnygT95o7M/6xPaXauLNeCtg6cG81YOV3/SnfGmeBw
wRl5MplwZtJVqD0EMjqSks5VpB5E2KigEU1YZZ12Ne3YumTOrm6HyYTLz4jC/D1wIJVHwISXtV5W
pD1W5VmiSDrkY5ul/ZJoitM0pew7NlDR+awm9DYdUnn7QjBMOQYHMIdEo+Q9sN/A+FfBrlAXD2yH
y1mtD8v3vKBFWB8ZjsJJ/fGyvH6mcRHxdK0VUA6gvPXPxwShV+oQdHr+LpsIA1Z+vfmKKxRsKso/
avA4tqz2Fu4WP29xYmixW5wJGLFNAz8fZrz1h3r8WizwPQBfThmncHyGJMZkAVex4096X0fCaAGk
5n1/3Ik0qSXvWGNEQ6aG+fFJXC/y0hX/LZynVQd+ul3vV2RtAGwI6ytnZfHlyrK78eRCk94Mo2Bd
YT6IrftaKWcVKq/eMfE+kWC/g3nLHE7FFJqoNHnaCGcpieoU9RxigSSygp7TOMIHfVnRkv2SjrsO
d03SyiXGsDkJ6pjSxUu5xE3e5xF+8VrtOghPl9LvmfPbfXZ2O4c1dZhtyxFsStgkliL2MALapUzo
XbbaibN3hCRcDBO8GXFrb8C9QDd9zTX23bEoUT2VvwiIlmqyAr+Zab4IPUftK8jcwr7wV05Sp3QN
4eQoYKVNvDLvLOLXrfzzGLpIEq9j7eEjd//7Nr4u1c8qeFAd479TdjqSXIeKTWUh7fRYfzJ03Ysv
D4zFxSsXkgWE8k1v3UPs92lot9oenvrzuSNjtp6JFkgDU7k0hmo/WM5tIkMsoZW783zQJGIm9owr
p2G/uzJ8fwkFs9Ps0Z0OisVYi3oWpsqJoKX9AhUAtixnYiTLs6nkta4EN5OMt4goTXU1Q1c2ESwG
cqFNw7+R9AHo4eXuuhdO49HGtERbNioTCHPKtX9Crj1ANXopYAbwfryzv+x3YadjOtu4rbdG/iJI
gl+tyFeVvb0szAyGL6rYkpvf7BEHlZneXhs+T0dnym7J8lVqtvBYjR9fYV/3kqQYXft2qTwfEx5z
wMaSeU7lcGR03ns5Lye7pEP5ohYaNYBQ1az4UW6epkdbJm7QUPoCLHds01SWx2o/6RIEi2NWR0FK
4NJsjK7cExdyFSBtUt778BeR0pAyOwgLWatSucp+jbN0D+Rjjqvn12mD5X3L30W2WA/8UGa8Rp7G
innPuOIhOz9VqKly1zGHPNCNJgYZ74muvZqaY9YLz7ICzzIo5/RA7mwYQuXb8TEtUe2F9RcwkA+I
dpZUM+mdemVoy+v4WYr1MNCYuAsieqUm+nd+yzxS3Z3FPNTkOV4lCjz1o9j+3EkrefDQ6hsKjUwo
Mn49c0X6fdWRZvHpi2kGWsWibStkclDu6P72On2noKyKdsI/wu1vaQpz7x7BZcsdA9OoD+gdzf0I
uTDIM2PBYVdwHkrF+S6tY6alrdoonWO9qxPk3ez7D4TDl4HofxJpKelLxOeToMYrqnkpEi7SO6av
1H18HKPkf32xzwsNrK6ECQgRZzqKPP8BD8x6tefOOI4BxCY4T11XVWY2QhpRUsAl6kitI1VGTGst
B4KerkCh1sGn9hd60FldT0O1GaSBIvqw2+DtweeeoBeE349LLUOs8OcZ3va/4zbvqUaeTJvIPAfP
e5OGGUZoiJg8iHx/6S2JsKTBvnbMBLqDc3YYDqK56JTqw37gI1VWseJvxQLQC523xNS1UthfTFIO
9zap/Gle9bA92cr9sSve4hI6m7tm4jjuqpl+WTwFW7fCFIeHMrJkvDEZGDVBlF4yz03Q5XSrqWCV
cDGRkdEA1Fy0I4JKdX28fk/TrMYIsYR0bMT16onUNL8Y9qRE2JaiQa9yJj4kvaah8xu327IyGBQy
grJx4mG+5e69pqWU0jslv+uGPYVke8OyVqugVb/5f8DKc9XKLniOG+nGIP1TsdyuQrxfUGXLTW3Y
SZP1DwbJcys/XeG7WuEvyzs2BJkSBOiFJOSOlzUwhZLXiPk8tzpMeMPK+wYy9kTYiEUNcbClMsEU
Ogdw0Sk73UM4g0uh3bgMiBLZ4ImtUjoTR6iXR1ltpbTbjgOksLeuA/sbEBXiyt4XdUzCnp+SzIC+
PK/vTd4DOv1ayoCdIjre3almgVfu/jm0uIk7xteGf8DrffwjcbVchJNpzcrdI79c/J4X2+YsMqlY
EUsX5Jh9NiDcxHGPAMNy5w9qH80j9kNIRLLORlr60+IC7v0AQ65rtVk4sgwE1q2wgouUCf6XUqCa
y6NUo0r6ryzIifCfszRcQRTl2cIGJ5C/aUIPNqlfq81DhS7mGWD0kEKT1IKg0KZyP5r1ZUFGjQpe
ofo8JjJLojSyKMzDmb/YJ8iRLVqgT8cMSS5SsOKSot/yIyzLG+gKEzakgTQYUw1FqhBBB1gZ04DN
7tw3/V4U0yYEEs6yYVdVeKIp8FMbn73RAPEcdtCQeC1aUdPeJOgDl2NntXTpW7VrTWCaDxCaOfkR
UMm0SMn2qz2rX1STjMNsIPI0EE3pZ7ZmgQudQusmESsxkNaT0hrTmy9eI2iO3yc02AsA+fO0scRa
63ZlV5ccLgmHVDPMCbd9mh7gneKPW5K0jBqeUSKL468IyV8MOb5rmWa3afw+Xpis/VwoJOkVI6gw
s6QpmcvRy3VwOGAEkkaA55iwbZQ3EhjXWP7YMEowyUjAK3xhv+5TeCSnsj/Wm61SxAO7dfa3pKpx
PMXsGDLUvVE1iaixvs7mjRPiEYLhzY2lW27V0J6p3hGryzI1XYwf1ngV3mXCSynRkjCSCtsvaLnD
315kzNHPwpXYl4mp/mVSUnAFyPAVRwkfqEmX3M9PKb2IPmmIpoRPOEeOrk06307DSUIxllfri6XF
06tpGXoB728lHzm1p2iF4QpA/UknYB+h/Y0U94RhDXDiRwDbnC+t+XAmLE+1pxDM1IY1+QQ2TEyC
B+f6lnkCSE9as1SZbqL4wbB1izPcIQIx6eKVy8KjdvcZH8egFfiAxCf9aADFDeoPIPVynGtdr2uU
C4aMGK2/SyegsjqL8YOZZbRUctLL0X1+VXUn1pGxHVSP3esD64iRedX19hTg3ltX6ApqGn+9nQgs
xnU1OcLOgkYa+yD2hawUVy8TgitXYicW4DoAq8eh8GI4JjoMAsjF1CkJbsSHW6amUWym9n6ctJd6
sWAEZoZsYDbLW0yMk6+SNC24SdNsMPaFFXSxS/fujWArzyzEfygVvdJT104k1Bt/NflE1XWli2MN
uKvCEyd3QM1n2RPiv52j8oK1kyz2gz1NNspR7XoBv17InVIqyCIcXr764bZY5hDfqdd9LHoR0Y97
DAcaGOFYKIlk/yhiJTDvTnOLEDk78VAtMIt/a8syVULBmGPlk35NP9/VHd+9a/sPG0cmCIQtHc2n
KzcZxMDM1KL3aB+ufHha+sh6Qv8RlHrYp5IDTbimOfLMqTIpj2C+hHIE8n9X8qHgc1/5Qwbv7tmB
QdO9DXtNMAKburP6txJ676hBPDiKLzuyJO6gEEErhuFqrcIAn7WSVB+wrKQZjeZ/W8GM6U7yW7MX
XgtjcYR9cS7tdc31/tSUuTNJK0uu451J+MJ+3KmCPjqK1c6BwAsIhG3BH7gfJmu3NYCBmprNukmT
gxS//dw+tdJGOGorQbRDzx3D5S8WqON7HvPtJw+x1yIaaDqfjEMFPnpCPd4osQJ6Ea9HlMxjATUp
rjPnqo/e7usa10ZGEGbvHxqmqxl98Tz2QiXGlejD53t8nHKy8OYcNYUNbZID9ZBxWfnsmJF0rk6M
78KmPQJHRC7dsPDnM35CdRe+lc8FrdWQwcd4N3ePBqUYREEg5FG/FFgtvAiqjC2NA5graaiXp+LW
JcSieL109WTYAzLLJhcwA3Z50qw0q5nvMqEuRwbOMh9ewANwxIVxPmQ/BMntMw6A0XApMEGzA0hw
cjiDI/r78OpOQjvWv0mrsYWy4AazzT+jjKjOggwQ1vrIoKaxyqRexlsmeiZtK0by8KvYFt5eWfZU
HY3O4UlHz3BBibhQmFkbjr5L7R/tawHmL+GP8crJ3pL0DAUu9lSX8tQlvwqQvq12Q9L8NwgLk/Y4
1TtGc5lKwAId1wQpszmQF4RtxilgmyTnsXKURfPy9WO6jaknVp6FKqmqy655IisuDoGnKr7nG4jJ
akCBSpno9gnZKCOhK725JWti+mfiqeEWjLWj+OMSpt/Bmvul5849H1EUdqpLLBeU+f8Y4isg0b3s
vAgw78cUyz3/zTq/JJ8duEAXNQbKW2B9a1GMvfYzNsV1kfGZubMrlqQUxixspelWAWrjr4SK8rly
R5N7252J5Vf80f3BvheXfDJ6rJ+IpkIrIWf/glVNsRG1vB9+BgxbON7eRVXdi0gsHJtgzMi+ssqz
MbxeA5F27pfESqQWLo2UdNxYhkNOJm0CdFH5yLWkQm23vqsgdtIw+StFS/rE0Lav2L99v0zTFz5k
1cLD3aur7FNsITgORQDhbV30+BBPrU7ZGGuMLDpE524gErJhCl7dC+5PCFkg4jfMB8dQzQXcel72
SCHmG8FnlvU2YRNzmdiYrysSFDcKrEqzHfD80hK40jzNWjjfy8PbD1g2spSdJr3+YGMGZGm0B/YT
lsrAyMuSAErGqMY1wsbl5tPsuBwaG9KGRM7A+HLDt+BwFGsHyZGf+iBWMQMYFWUYavuCrdU9xL4F
YUxYHE0htTLT3ByFEVmpM4T7pML7c05AwRgoQ6FYqV+24LAOGNm1yEFdu+J+QiSb4jJub4U1bxm/
1cN4ruWNg83t7JH9ccCaE7egiTQxjeUsnQfTKDNmtbcJAIrsHmeza3E2ZZNRI9heMu37x0L6ytQx
ClFqHEe8pNAUY5PTn/bX2QRZbDuOJYNPGp6nhGlr8MuA9UNhYWsD6FRtgI3thyqafNM5GNdNTsyk
RFP6oXwlUCh/uhMc+YhSY35uDH2vaFsLZn7V89EDjl7FMM4381dxDLO4rFHjYOjN/9gvrMm/voEs
rlfS/mCN3riX4w6P0+YsNKQbRgQK7GVW89YPhrGy3/O+fEtQYz+UKMnXB4tFN+Nxg1SXuoZJa+Wt
NeN0In+yeJrgytPXPW/QPLaBDgB5fmwE6rNjieqPqWpBQty6qPCMj2ldMxXGKZKMFPwaPpns0HRD
xYFI/tsFcMYWdQmmL3LJXCaOH4VG3p7pbwSiyhOiYUhrG1gstmxzpW048yL0YaswTFxkeqZdH452
Y/mHXr1yAUQMmnUz/KznrjhrY9sSidkHbJg/XFJmytv7GHSJLr8TGXB1fDFoKf1H19z0E9lKukfi
x5xuQ1P7CFuW5Xxt3LnhTodqbkw10eLL7mQ/cnMfTQjTNJ5JHFzlv7DkrLWY77bSk1qLUjx/+MD+
T+0nCTnKgYnkw+trBeu/myn5lQKlFnwHXlSixordpjV8D3KW0i/1fSzZDWKz6ZWBRnO3rQHikJhd
U4pkzULNF++Be9zIDxCXW3l2lV8LkD825dByx1QESJNTCyBAuxwtBiWYxaSX5DYhv4LOauaZ4frM
14PIl4zERYufNNY9JynCIBSFrcGO6r0hmxl+OlyhW+CucG7l5ixhIaTWYd2LdZiro5kL/rw4i6Jd
6kWKO+XklzKFlxFPyoZm0MJFj+w2Wtrm0W4IoprDyuF7jwtOH46xJAWVjdyNGDuDLzgXWTY6wyHx
RJf4ozGWz6xPhIJ1IV1ekv2/IgoqIMYF5oRKgykYK3tuYnXUt9H0YQI8c169sWS0V6G6gxnEtfzS
21+UOXQ+hFzia/nMN/FRPy//JpAzjkI0O1PBbKT6j97TCK33ZXUd1mqWR2RJnIfsjyJ0krxLTY9X
gVwCNxH6MZkM6qhy3TyK53Lpf+wrY9uDZfN1R6wDud+0vrHWKvCbZV//4dJNxKCnSBomEzFFT5YI
l7/W469LKShnIhHpPaXLOTmnklJkTo8HyWDQmkdfnq4uGD4QeOobQSZYsUL1wog2kyowZKe6I6m8
4ERWBeT909OVT8UOjjs7ZyLIisbu/euHMRiGQzij98bTV2JYDXd2Eji6froE51yq/WCXzQ5BvYGC
Q63k5OkiHaq35WsicmUg/2/t0UtyDFvPgOvx9llKEsR9r323QQbu2G7SPcxYAeDHLbRpuc6bBGVR
DYBWwpWSdaXMhqpuenypPCf+wNmHo4QwNJOfjj6V81paS8o5bsK7AgH42E7d3Sf/jSmJmaQeBEdS
Oh0XA6Rxr3LmcrF2jgNRiygN0bNmGozu4LW9mWpTeSkYyrKRzqsVZm/QNzRtFKwgfWz9Z2ZYO7rB
oKIlMrQjoDQNhaE3GlNpAZuqsc/USaVjQ+rsvJXFIipnAXV33rb2ZmonmYxO6MVnMq6ip6sBJayC
wMvyosarquxduGVpi5l9vo7e0BRJsQZFamp/6JBIsp7gA9hOAbSwtY6ImCUGh7HHtKOB5HoapmrQ
nH8xgEbfCRdX/YJEN1mFYjXn7FxMWbsh4ujp2JrM0fEXyY1awFtT1tUfYg2o0oICGuDZhdmL4D56
DvadV14wSLhkRUmLuAqlJ//DYgQ3gxCLALZkhUs78pqfDSrMu4efiXUmRXwU95cL8C/Kxl9g2yKf
CoBOJpGjOcgzxF9Iy17FcOP9sWPZDUvcOr0jrMVwXYH7ZJ9QuxLbgVAP86if0lXc4Sqrf1WFIKn3
rOQN/qKg+T099HYF/BPyzGMOL177OC6VjT+LwiDhIlTZu+cVjCSF5ipX9c1IppGshHtRnrlzz8t7
djaYXy42Y4PVtDqhhGMfqDtfuuGQbBEYd5v5UavDq+0SdTVs5lwH/e0sDrJwPvH7a8ZsaJT4JwAH
+N3a8JQVRysRbUZQITaF1obq36/Oy13AfpIyhQhb2YIDT1UnSh+IbvfsF3u0C79DoEYtxtyXVW9y
iOjCA5A9OY18SVp1NUr8x4kTe/taACF/MAN9D8EJPvvwUxzq5SOFVUM7r8wE7QaGcavpaxznwju+
WETUweSISl9ppBi0DAQT0vL5qsJSDAbc3gEqCFsxpisvU497H/SqIzz2J90Zsh2UJLMpPGjfV+YI
8cPVFpZK/ReNJ2k7L2jh7kKlEm/DJXKEezH8+yab8PRYG6Uooi6sU7hpYTe250oe8N02MdszBa0k
p53Z76MGZ7tm2oAoHqRVWtoIxugExdlKJ+eM8FJRzlJqGsJfXWnqKkI95NyvNblDRMtNRbP7ZMrW
q0naDLlYUF+EN/1yTNBJ6E/9Uck1t7Wh9J+LpGRq0e0nn3L6AFjzpFjJlD/9nfWrt+NviHM7IfiH
q8daGiLCT+dtKt40irPpG1nJo7/MbZV8ls3upmxO5y28hgEwFFhFphnNLyoUvBcHNnwY0j15Vbta
49tvxJ0SfWjSFUvTQADe/juLPtRDpHVHG+P1rz4WUGLdWvNB6Ylp+cDbP2e+XWcKL/cGmU8T7qCJ
I/GVgmAsnxZ8JIfLCAX1lMCgccvwViUGgX+xblfsxifqA3ARcJpvjpkiXAJHriiytYU8XDpyniM7
UaMLoPVSLqj7dl/2/eVNEIDyhSfGY7PPTzeEinWAnHEcoz2P58esAyWV060TDFwWIuAayBbrRqEG
zcVQRqWdcDC+32FC6svomlVSv9eHDemrnwARqD5Y4Eo514BjiCHUm7xevGE5SFeaYg+iSYylbjdP
82puqec9WbCXmDd13GD7zrbxYG8g12k3lGKY9Mqn2NJjYlnsfDCEFb6YmiP4zCzPq/9M4HEcsmyg
l9zrrfqNAsd9ZpBlhxnGJEEE/V91gAvKHMhYhhz9X87vNdgzqXbNNco56yTcr66ejQ6m7KebwSfZ
h0WU2kwOwcKA9twn85TcBCZx+02cEDrJusg9qwCFUA/s60m/Q2HpOFsCTN+DJ6Gtq9vYl9FdqJkf
MSSH9WfUv0j+gQPPX3Q//wRsb3R60jvBQ+z8TbhUl1pQnr3GD45m1kSib/VTEb3MezByEi9Iw5ZY
ceZDtJyq0UICorbhJtc4KhYzuL7NxDfnLowV4mgNIzGm4QFyxolgROy4qYUDGT+9WmVaF5X7+Vgp
DMVZGR7ibEcH4xocv5QZs2giyLuIIUyw477MNneprFJD4mB+BNHJz69rYPmTuBitFDpzVKzCVgrp
iT+V91ryQx6obUpuOFuVGLH9h7CBAQJQtCr41yVlW7u6NwFWW65sYDAAzOaV4vEBUM75BF00xQo+
mYQTHZKSqSvUY9BxR9k0lvw3IfSsS81jR5nKEl03OhB6QHXZCxqjgCJn3FfPuMtZ1fW4gXeCYE8q
+r7RI6j7mTUZjP0/F2VE3fhmQQxeRppjq/maql7ILBCRINT3a+Sz+eZtVEG+Lw/q0wGqJChd5rgc
ye6qw2+rwdFO+TAJkhTecsYZnoD9IbPkv0M+/DGtkCoDFEe7hVC3MiRisbsE7GcAwtRBmIWad3Mc
9s6fjCa7+80Ax10V9bqnT7vfdkVhDjRqDDx1VFjUBonotPYQGvzl4UdTQpxSiHDp/kI9MLaEtxWK
/+xMiI/Xxjns+ntMrKtg4w5nJrSXuEXFfD9sV5neVSTLwYr9YcppY0cu4vyqiGnsF4svqmpT6IKB
Qoa3VMwe2gzgeQ51p1RRcCC/ihTPwjlzssn1e/stxFtDPSxf3d69pBeqL0wJh4X70yFQ874yNUXr
lH7bIqAL7RGg5KgwRZ9kt8pNGlvlXJWYWDqDOr69dzQR72GJVgNWAyXl38q+c55gvuXtu9FzLFQg
wVk8EOSueUGdh0zBaISb6iOO5qp1TL91TWbYrPqG9Nj0TYPWYYUJwz89xT7/UsVrmkfQKgJfmPJ5
e9viJ6MtdjQHw1JHV/5EotuQhqIGruoYGh0tmDhHiGDpY667FF49gLahUoBaXVppAiyR6LqW2fUX
2sUkCTRbtz0Fop53iWesTr7vT5LpuG856znxEpcDSOLJep19Kcw4T9ufY7WjFwfLbq1+f674NGNo
Cdq1UllGDM5GQfi66l2Lrj/R/Qpls2vJ1OLHXVc4cxlfHvkbMhmUeFOhY8OtzECJ68rm8jfJQQ/o
DeDz2ObPiaHrCxnhvB5eM1NUIdzHj5hIHOJJWQ5eqRi48T+WaT2/Nns1mSSkuejLd1Nzu4EMSh4w
DWJXlmgfeVIcQH9wjMMVnYzGcYr3gM+G4wK/KuwU0ETH1ScWKReYvNut0TB2cgD5Ey3A12Zw0hOj
KCWX8FtBS/zC936/fJHiDWswxlz6WNH694h2YiWp+NuBnteR8Wxxmrq6162BoC5XbaeHnS7MXIlU
Jta8q/O9B44aKTbHHmyUPVky03kWSgC9urY5b/Pky6FxGE1adrWgv0+uDp/EFSz5/2SDQ1dHaioj
y6kAZjLPDy5eLnbfeWJ2Alxm17H7GdnXy+YoaUHF8MSQwPNWy2ugfwC+UOJIVRYMuPRVCxZb+mQT
43654nQk5ZGQd+KPmValHLZ1puvmdaZGPikhFlJJ5dilfLElvsQQC2zfajrlB0A3014LidenAsO2
Ey/OItUEe1TgPa/QKDhwuYpXIeDLSb5+Gte/lZs9SR+lE8bLAhmbBpAPDxKm49l/H9v8rlDWeAFm
MCWhDMM3IBnivCZBtX3J8uK2ae3nYfWU5sGOBZmN8t4VLNTLuqntWKRLJgJ2ZQe83U5NCvObR6bS
UTaGZtKTGG8nZZ1c/XwwKFILeL9P4WwsFKgX1Y4nq/eIUxeJ6YE4Sh5a6veKmpj+oe6avyXEVBZe
KSrJTUWtkqNcbVDh8naCTa1Qv4BWIMWZvQjvYqZt5FWmkkKruc4H/wTGNzu6HyYNLQFDwgCCbGH7
jMijuCWJIhgXXvJiTCWDcqahZ0yDG6RCtR/PMFs+qfTELt2NujgENQmVPekNL0kkhAyM3+83mipV
YYqohzCmk6tzc1G1/sZi2QJ+OeVWV7Qf95hpJbp/Sz2mSyx9kuqxOGb7wcdu2jRcnCVP/l8nqOkY
f5khZihDTPC70cfq7ybyPRzpvB17dzBP3NtzOHAx8erM5CmYjj9caGERN4Ge7tx1X3fFXbQicSop
bdMruEjc9gBHxs5A5AeFFrTOpXVYrcKGcKo4aPRVRYup14kQk7/7rONdFpXHVwpIuvlYDTLAHt7R
hpvKyGFxOILfgCNsGRjs7viOse33aW/IYEwbbxRrIM1EaCo2z0MVdnfaOthZZGpOtpeaksnuswL0
VDmTPcv67fDGdk2l8HOO8/pQeLxq+ueHJTub4lJEwERg35t3XsNlnrughtEauydhby5wvr4Ysbv6
PSDyh7pCeYafZTKX02xthoFpFKGRRyGy7TNgZWgTyvrjhTP44dn8rXCGrkwLCfhN8HGF5YL+8Z2y
yqiFWitbGgL6xUAGoQWP8hM9qYL8Sb76cMMWW0sa1FebjQNw258wkYa/M+15KjWZJTm9oJ0Ebydl
8ogBVVBLonyX3BB+3Mck01bEUxZgLmhVT7kxb75SIkME4/SkjgWyDqEqGtzKMyq19ODcKYmtyv/7
OXAgZz3V40LgxjS2aCMLRwuRCioCKHnBuhO7U1E08CQXvK8g88VRy5bdobpV1jGOugYTl7k9IKwQ
v7rqGgAzaC+AbEti9YXApfmJlecYU1VI11ddTKRQWc2nVWvN0lVow80e39BfO/RhvhmFZowOMQ6O
xfIE8YSrxz09X86UuQec1OOOIBM5kH1Pqmv5UJsyRaLCxKI73HQnNMBiPhgrREmfoYFQxjxYPNH4
wgVlWAWQwNfJMc4sDuXNIuk1h+fu7+nETPBLupyXbaZ6htLBItLi+DPakMVZw77CD8HALhrfDd5O
a5ktm5Sp8QwZR4THmrm5ar01JOBa6WaK+UNDKy3PwYUlbSIKQJMr9KIYoFzrV41BZNxkpDhmhv/g
xWZpYbXTaHuUcNXgsfCuseb7eOaigRgc5MNnFJacjzQhmI7F2hHsdlAwG15EATYFuN+lOu8oW7SL
Nr7WtOslrSIzB6kuZbq9zKTtCoia/8Tk+MHtYNgJUjNwpwjaNYH/G9/4bsO/bKY02CJDWP7odcvJ
eD69WTnxzwVpK2csH8HNScMfAVbACnQPU8G0D9Lpe6iVc3H09h3OsoMTBt0GG1V/7jz7Es/bjwHB
WZBB7Pbxb/neIm+G+XewXWMaZDn5BH5SinRdr3H57Gz0ssGah9GAPQcm3z6TNcjssVzkR7qRbD08
mQ0UqDDTQgewvFkvCrpDSCuFmsMOaMnPIGnJEKBRCENlrn90C1fwjnbJPGjOlXL4I/OfNDQ5FgcF
6Rr49G5HOKxtNVU/mRI0fUv1k9e+tW9fXHyNFaeqnLFQEDeCRU3HdwPQnjGuGQiRKBop+97sdWci
rjpqpsAuowKw9dsPNUsOGprfxBKSKA65Iad1fYEFWb+zOvGRb2jnk6FRfRSagLVIfh/VN3sA3UV3
7xd8CSrftQKZqBH7vKjl97XZCuzPVkopm7pCGr8yHXDL6YyhiGIOuySvzzu7QuBVqQ2iQf9uuLD+
yx1KP11HkUD+l/fOuJDnx45CpTDmJek6mALB4dryJWsRIRsJG+WVqTyQTHBnfj0JPN0MOasEuOk3
VLXVSEifxbaVf0/9KPLFg1/Ndjj7kASjicuJ7jucBzvwdZqCb9EjhIcXrTi2L5v4PdSxeEMoGQo4
iM8oWr9WymZ4/C0UTHApjUu91HrzlAZMd5xEUzlRhUXoAn0BKr9DSzPLBV/pHCHQkB99frrkV2vr
zFeGvNkJdBC8psXqnLgistGcWIKkIFd5fcANGSRDimd+05sDFVEBjVJs/z22bBblVctZ2g/8+fTV
I2acGfmhkWPefRGSJUkvGKWPNB5ynHKxRqjj/QPJ0kbFhdJIjHgkj5473C4W6CVyOyweao5jWtrB
oyShFJ3R+12YXPJRDj7YyoaZ7sXNRP5fPLiVh6lzlIwQ3Tts8/NjYHBmu6z1xmysy1DcmIS/AoJ4
wXWKjDbGbaufYMFFlcTztJYf4uTHc2lSq9eCD/KToJ9R13OSb9k8jveBAhIYuKVndNMHRGNnN2Cm
xbbFGHBmJKBOGCecWBahV4Z1BzTUH3zYfT7H/B7kTGa1Sc8mMF65//wwvdZq/4n46qBMa8MhP72Y
kLBdBegOfPhnaMelfXrM5uF7at9T2PB9rmbgWna+inCpj93rjUAnw/5Dd5CWwNE4WrMt74I2KvOA
XP/XjyDTfICJb58VdpKGer1rXYJL8cbEVyDaHbszwyhzua+KIBMSWy0FnPbfV3e2aS04ek8t6ae1
VVOmusAV0JNxoWNvGsyk9xvJ4BTPuT6sKdV4zf8Hf1JxKqhtncfZ0qxVQNeOX71CjlcBGWUtuUdK
XygqmnDj+hFfqBojJyXtdsHd5RUkhPlHSGe3h3XuMqaso9EeCRkswC1Nw4fLuo2xHwmjUKLDS+Zw
+F965L7tRBz/+RuCYNQkqVbF3MOVhbigaCCXrcPCEvOezL33a4iXEvT2w5nRlAw8O0BAJZvXW4bX
Y1SYg/vrj1OHZqdoHA+agw6xL8tgQf1Dp6zxeqBDnVT6D/itSKYfeWMdCMSxaccAdQ7/UL87UbjW
wkgzSqizzgJbPyylgq+UGuYMopxUT5kll7waSOfrc0ZTrQKk93JONyjHQ74K8mrZ1/HAv1CGL7sq
0sYuxITEbQ/Kqk3gXauJfzgwmWqhoShjSwNNdmZkg2/f8SoPvpb+JV+pHVOM57JesFB5Mu0O2p5u
nEUUjHfMQyJ+6z2ShC2qMmBNityrfdprdlp51bffJIeqgupKjvglxYSiMak12gAtUYbqIByYdeIy
YgqXHCWvfhWA9Rxv+hHGtK/A1/KnquGEBktH0PNkhg64xURecAGQ2f+YJVDeOIHAqQ8v3QXvwP9n
GL2U3M0357aL9CfUV49p1KiIU2tkI6kP
`protect end_protected
