-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AFeWVwcmaerB2qNDb7zZ6jd33hDhCPXjaqQ6I7rExcFwLnwPg8dQJy+zs6LWm6fSGV0fg6fer2KA
bzHJ7kbXPv3IexcNTmwvSgv3WU+g/clnur8Bw6vIE6SiecHzMtN3Lzm7+SEwYHyLLnjnklHIjZkx
gZl4v4ifGjyl0fBvo8vdp77Q0R5J+qTdhvpjXmK703+9drFY9rLq5llnOBun+p/0GjHmmVjcWvAb
q/EvMC0Ozf2LC6rddL6pmQfBT7BIeWR8iNCJyqTIPs76w6t+NeyEev8blidsPOPLbwISfczALRMI
i9+bzO/4gzTRKX7PCD8ERyTcjk+pCkMtcYfDGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
6bUbjT3iAnPv6wW9eDvGH0a3Q/3VFMNcAxiU1TPJ5pu+39mf3taahnhEsTuZrCCFz4QK9H0s+HSt
Mmrb3LyBIVFgjQv4fihvkzdPsPIFvNr9/an/8QP71m6BIViVUqte26aPRV/jubc1mCGJtmit86aO
1V15cFqjB3TZQo0mI+wgtJ9QA0KG9HeOxInbngPgtnB1sf2s8QPe0jmrbjF5Qp8HlB4zGmOp9pC2
V8X828atUXvqHlfsAIgmzMxI1oRAhnt3TdLVtdNsGDqL/UGbUGm9VgnuV+R8TjPB96OXgK2fjz+Z
hi/F4loVNYwhjtpj11vlRef4xAnDiLHspRrLqhN+/azkXDzzky7ylhc0vWAXcbfMMfef5+6ILIs5
GhcQOcXqn6zj0Oncbaeq6BJiy3tV8Ua1n65GH6rSCAii2EDjGc9s+V/YSKF7U6waH2M53Y90hV8I
Jvi1J5XlJ3xWMzwW1Sl3vSzrqiE21Vx1fY7wQlqQGB2J7UFycyP+NuhfakFHcOE5Q6Z/brIuhJUR
Jx9+Hq0bWkX35oJNUH6r5NZ0Tv0JZkaXNAcbVqMDr+AXFGR4c9hMk67ca3ntt/Ystrhn0aS4ReBg
AbigQ+kTHFZinvKk7TWcJyeWR5WC+8W5+VIIechGyE+NZ8OdFNSK2e9ILr99veEcasFZh4QSSBPd
wU+lBaM7DWd1dLBr9cbyfLEquTUEMTsXw/linYk2MI2OmK1QdhSFR4dR58WN2TnBJLUnSwwiUYEO
6Q1CEEdwDm5MKNYEeKItNigh+gab30OPbunwLOzsDFEIVXgzkSsMGG0u/eUQDFKoF97KbabLcr9m
/AfdesMKW6dxOVC4O7l6tdvJxOMh0r99OmUzn87IWjIySJ24haPZPPy8A+RXCXCTOWEN0HB0sbiZ
MQKeQb6GlKn7ABV4B6lpeVXA7THWqr6dqJYdLD4GRiefEaXCdf9FIqy34v8em9U7Eo1yvjliwBbb
UjkfWVKGVtl6/leukm4yyAdWdl9Yxx8x/g/0AcFxUvCjGOq+tO6s/7/5OdPe26rdd6lvKprEVbgO
m6R6IbPnoquysj+ZvGSCljbF/R5JGCTz8lWHsYFtIsoYbf2BEHIF1cX7+LAYM6Eugh+3u9FFow+p
3LQqmyECxR1RvmtyoIFx6tWnLSNNmJEZl7Nw0l2vERlg8IX+ELvwRou1Pkkm1xuDA0PFRD0N/DsD
YBrtpfcSr3ngCDk5a5KaUf/aE3z1RgjmoT/IoHfJRDWJrs9p2QMPRkkgexp7yRHB+ucI+gvkSMvV
dRusgdBtff0yCCwKG6XCI4hqOkWR8GfZFEyrv6J6gsXWcMrPdxykfaP2V9ID8l3S3o1ODh8AEfwZ
catZgOcREBU7ZFt233FJtfuSHFJg3DuCiyjoIVN25l1Ov9rg5KmY0Qoz+D5TiRTikvqvbwFTesan
s7Sis/pMzTbbkyEplqacom7SMa1RItxGQaiZ+kMcvoGyr4/KgEYk1zYkYPkaA3bFMI+Wwqoi8j+F
iEZ/Yp4LGkLnCZwhlZcSF7TMZFwx/Nqllj06GDgsmpaWcmBZCPOczubEk/3qFmozgqswKOoOCMUX
oOysKjFxjXdPu8L0E6cHPNLR2ZOcm1YXzpXKd7b48J1gUk8+arHmD6myir2fzQA1Qc/IInGLZEm7
DAuT3+L6q7SPt8ijW+AI5NuRod2P93rHuerorQwQaElxqqDOM+Yqr0qu9AXkBOEw8/RlonV5mORc
4jYGT4JZbyI5izbAVWGNPvwIHWqEkfeUojeBSYGnbX9QbUv1CKwlJ7DYx21KQyyYrhg7E8LStRyk
gEWB607sIXi13SRjEW/OWad3ykuzIa9oE2P9MGxKZGR4EQ5pJVdmpW0LBeN6YG160h4/+d1tognV
IJ+Hfd4Euny2xUS8JtYUzhnWDxV0HLHKdQw1uWxY1gbwmrhS6nqR7evKjrDV0DeisZaA4BSxP8Lq
XJg1BTayToqFNrnE5YjyF/BjPBEOECZzC9CrJ368J2/axOGUuseO/fhX+GwTBr+lLHpGz8zvkjhZ
Zzf3P1m4fdIpdLGYLXbGWH2wzicajtQB9a8jeaMx2hwvxKwTaLrn5q5fuwTZEUjm9UHF9TXGu3K6
8DK/8dsmGbgOGLHAFkYeCxGTs+IeBuvMcHeQrtYzaWTsYId4S7eNzzvV88TscHVSkXoMs+wmlb31
s+itqwKYIN2SdV7+/88IMYTDxfmAziLO/Drsm5jTgyoFQntnVMiH1CDc6FKYiHLLVrWYeMUDjhYF
ci5qKOEikV1m/UoYy509kl09G2QfMBhJ9Uo9d7qZaaQqSuFNjXC8YyiFkYCdUSAcA0wtLv2dJh2Q
RX41JCoC0PMtHqzs4ALv49D/uY0yIEraUY1jlCMYfnqW9jWOI1yb68cCGk2PD2CL7V2XuQqGwJEJ
4svDbwNvdeWt8s92+eIQDwh2yCOLggC3Knv1QsoofiZX6Dkr/f1D3dJD63R63xD2ANxlRA0kbKjF
k73K9nKZS/S6m+Oj4OoYab4FdaDGEX7bwomrr8w+yrwvqSbrRA0f/7TKF7kZT5YCaofz0RUCadPW
8QfV20KCfxUUm1rN93Na+zSEpipAJ81TOSA6qRmUC8AKVeHF1h3lP1FzS2O/kf6Qzjr+C3N0LW9G
ad1cCnW+QBLTgubJYUb21M3FiUbs6C2gkFvwjjH4R6pXygQ9XpORrpCgq03QxfBJHka5hR7BrebY
fk4aOUEQRfej1s3SSnqujCKPuLZsrIoxyFw0U8oswXvZjEfzG9zWauwboFND9Ps/+pw2wVvTfHkU
expnzPiPWvFfZoW8jCDiFBJGxdcexzPHrxifLHQMp88+daVcauhvuMF09PV3hVDnpiGJsZL/cYsq
OEKB40rHTdxan4aQi3UKP6PCT+3SE3o6TNJ9cUonsyqL7Ak60gRRbeptWVfD9UQa6CnAey6QIjf2
FFMRArSQN/4tyoDAqTktoRNHtegMu7kfp7dwh4ewSXbpDO4HdJF1E+bLuWAjNG/RwrT0fDNpBhTH
wt6Xqn3DX9CZXZRbH3MLWDvDddqfQWg1IeIeNTimn8hrVfwRZtkgNyObSGuEAOQy+BbdwXvz54ef
S59LjnZGaxJR0lKLbx1uljsiSI/9gzgI5BKfUa/vqDdj8Eu488V3Rs5nqjC4gzGl/U5UAEL0BwFx
plimc6RDCyuIG/+LkQPexvxY8kyFbEQx3XCLcXBVrdpZxMCFg4IKSVGNRJsWLeE6fydIC/lHPJX5
T2zR7XL7nCXmkKakeXIWmt0w0G2Gth0BF2HnLeapYmti1zogE+YStfb+HEIwmpl28G6UF52PWyUO
KMBr1a/BfMo9Q6uOEgbSIbBuTOf4sDnxFX9GfNMaYDQO7EVJEtlDygQIzhUaN/XeT+xN7+jzjNMW
nV7q5BmA9MiCofhhTasm/FKhJVWcmDxII5tD9nPGYeOI1L5sP9orJAi6+XOYZthxVB4v1ZarWi29
QJ03HbAhZ269y0EFxOeRluu21iK1RF8UPLnx0aB4DnP67hmGct8U3Kk3UETRh4xuGUUWxGYilCTa
KbKxVUik5ai2s0hA37l5r94ZVN9QIC+PPf5kNCZb9dImIX81EKDiJoQrOFDPrU3eiCJ1cev92vYA
Wqb+fQ5+IVFZM1s9J5iU2BHzMkcPB87rGsjLec45VE/zrthXI/8PucDsFRfH6tCKNGv5ESWhbS6N
7+JlNR7Flfm4kE4okvbK1aMsuxxiuh/I3OzgUJN/Eg1+H8dz3tnrd8dCG+9Q8iSyVqE27jdwArTp
LPnJErhyPCJ4CNrc+617bdYBNxOp5f/IIXW9gzA9zBOV5SF0dkg8ULW3pnXqaSCGwJTM94Y1eui1
FBMQ6ey51LQn8VXho40MQO2HOjmySyUwehXjfYr117p1VWKkpdfM2hNlrXpi2N5EpOiWUeK15GkM
dp9q0E/7qf3hpJgTVJwNBUdON7khAKYadElOxrLdIpYgdZh8HIScJqio2DK8FQNM7xh12dVt6JXv
obgp6rF0V++QFSNpQddujhzfI/sBBXN6JjZgS4oSs2FZWJ+p/WGIMfA0MtFTPNGxul+IHdWKymaU
GqD/t/rPR2ovd09R39uArys99pjBnWo2j1FF18GnxX9YKtHjXy68956ovPAYjlcoDTLDJsMdK09u
GOBZQvNVZ8vOmOGP0MMGPI75+5S01QCK3GUA63tJwD/ZguT0XRNnP11KVl+a/5BZsXiwxt7zT90V
Ywlb/SJ6qxTHPcPdUjcaplyhv0VeC2HPRh0Kg8YYji6a5I6X1FCsTQJMlwmLK5dpDyI5ScKX2Doe
esykAyV+9KbfHRBu6h8ipugYTMIHanJJI9aKvewUsYsSHeT4y/rAkRgtZ+2v58jK6h7yqRguT7y/
UfMbpUj+v2zql8RZXfI4s+bVMECxDzY2Rp01v1EXmMQgANQ70PGX/dCeK51CJa5Q6M9kEQB+YiDe
gntqnyX3cleqmZORJM3G3vs7rqIsQVakHHzFeCl0f/uHlIzKZOf0/n6Zh/4HD1uwjs4/KFdXCuSg
VFDgGTyRAgi210jNUTAS6vr8eZTeibM3kg3k/+uL/Ni9XzG0V5h3MK1jNxN4ngI/N0r54U1HX14w
Gq5EnQQgtijFcZGWyevT3u21MWOgrr1zhQIs8ERUVi6wtkn21D+Ga2tsJdbPhc+FDujRjUlSoabf
iv66+kj4PTZe9xhIAaDOQyIPfKsW2kk6TrCY7cXwbWXTcwmRFE1EC/tWVehKVzNH3kFTrl4tl1gJ
Dc/gxVN/clu5X81GVw94L0T5BB8TZJq/uE25DHmmhUFO4nQrGkNcU4h7qHit4Zm2cfWNUyADjEQV
Zpi8gY/pG8FeTsfMZVM4bBoHGzAneAT8/PHEiHaudzcfZyfyivHLIamy85UkPNy9x4xA1XDt9EUG
emiE1lziY4+2X77ogV5/5yWjUaSAjcAQozf2Jv+fudsLrphcBvNt9A7XeKJVyXinQzxWGNp7D03v
ao7KP8VQQCRofyPb41HJniIQg4fNg8cZyA+4vycRxfzps3c8vDgu5d1HQ4+U1ouEepLXSNqGoDeT
gWQ6gd7kn/3G+E9ZIsHUmBsStfwyaxiWYO4RW/wqm/3Cj4H9k4vFMTpa5f7Dkq49c80hgDxzh36s
We8eL7FxmguD7tGs4k+hhNRiv4eh7cC+D5GNGFiAnlTTA54Eb9DjYYUScuxjov/yqa647GAPrm1Q
FIT7N6S+0zCPns21z4EyC1zRH6SrtPFBWRNVkaCHrn2Nqwfyjo/8E+BeFE23rC53Y9NHZooE7eI2
vk1wTbno5ic6i/1cQerpjLQzvOROyQ2/LjXO+z+BcYrkZiFvmU4yWKpf1Axt+IyeSKKQbcpiDcrQ
O5Ugl0qm7IPss2fbLBsS69LsaynJNg9UCWQrZnBtNYw0XqrAYuf7KvgEQC9U2B+9EZ8SfF/yM73v
2Z0dAcMTUAMjSejptRhJWugjkEzAUkgrO4wIYfWRRH85glAfwOrfBuojM40/oq7EutIalBVKRFIU
ba3ak/8U/DGvS3FtMTJZfTwnbDpG9y0W8fpGQPBr62EDGb4a43tw9sAw9KDq48qpIspZsJgYsovB
KTU7yIHqWj53RcBEwFYUlmUPMX6ewYxOsNBg8RCYUdl5u75P0J6zH+uTYVHbwS1wc6TTc6hCgHeR
DO1syzgly9gsiZ0B726sZIYPPJVuKaUeooVgDvRxWv/blacEWNh56C+1QzATe/THsTafuvrqeyBx
xk45jqhHjzzTKT7XamSJIYDBP1pQ5RoQ/GRiTMcT1dXKEjvDHMQacSmJEMSczEXfOmsrVvAOHTht
6s6sbYaY6onzMI/yG4PI3N2XANmde6NosS9igxthSAIAXv3blWYso8zMYKZA/hw2Z5KfhdtVnsQc
Dfz1v3t9SbrlHH4dF6EHTWDoUDfVckEdbQ7pEwXipmf03vUAi2pnKftSvmb122OkxWp8n2iu9/11
EpZKK0A3YqFzRRqe6FK3qa63NOngDrx+ulKc/67h+6UXKDbHa0FkUx9WIs+kZsIifUHjhtWgo+NR
c2u8qMTTo/Np+9I2TmiCGM95L0Tf2a1izv/lfzw0FgG/fiY6hEBXA+41H4q6nJT72FnlusiWTeLF
myEMCA68mheq4HRSyC80w3kgtp4+fnQPTfMgaSdR4PyYwclkeEwZGJYkwZwukqndnxo3Y5DbVzz4
DBGobUZimoa1CF+uGfRG6i+xHAKfb9C+1+XIzlLBPYuRNemYGjsNkUrdrATNdPEyvjxwZit7tcWS
QRxyot7RLYnv3Ll5fOG3pPT1LRn4TAwnyYx6AZovK2uBxDTtReFJtwlEajDawFmQRHH0c76y0MnG
2mH19ccDmtSh36uxSizw89a0XkC1f7rXhp6sCspHYvkEYwZ4OF7LVxK6fegtZ9ADM/HaFp7DDNrp
5MZRkAPRCB4dPNVWbtHLB0Kuv+Hof3F+VFTNsZBWuIvidk6MyUDBphktTHJhWcteeoxqf9mZj79z
FNduQayWGY9cbWV9Yq1PD57kJWF2gnXsCIdu2Xp6gtmP7dX1paYCPrHFRfiGlnsHXril4xID/mii
AFGY2V9zPaBHLgkGcWGBDFbssQnZqEd+LhouBSq8MAZeY6jwoUZ92LeXI0cd9ke4y8R2duFxIiSn
C+Zn34YBtnXcvF9mrCdzsNdBWvPiBf8tk+GcnOQ0DEKBdF+xaCKCHTqIJRnnZulTs/QBBhO+AJoz
XH8HAWks+DJHfy5t4V4a5hVVaJsejuq0hPpblSKo//5a7pgwIr1aRnY06+NDcUJ94q97mOVbMRu7
dQqJHsHtUSmNrJ+CAgqcBruX5hORoRCEpboq2OauWqmMKlYxQVM0a4lH3h5NY9mgjOtprOWEZkbW
yD7FYHbQVmij5Yan8Nk+gX2goX0lqkO2//cUGVUvtnK2JGYUBi+jogguNANTY1g+oLGgkS6BpPaS
k8oT25Lua+rxtF4Av4Hm6ouuMe3sb4OUlukt0ZoervacGBecNhCbLh2DxWUPlemTMsKyDItb09/+
X3a62do6nbBIDU/PRCqQU3ZPRE1oHdy71KRG0CInKEo50amBQmHceqvgSdfYF4taVkCnS1lsZTQe
kMsrEbTNiZRL1zbujFtzn1eWzju+Cb/oIXeGdpNg7ZN31w8UyvLGa+XZtEMFbnJrF0mUCvPCogZe
s0yPdWmYiI5Muwt4mI5OON2eeCxGNX7D5pKuurCu+Q4qqcktu/9KK0DWeQfauUfWxVOwKXYaW80v
mDF+8vQLLbEyC/PP+Bm5Hzxk0e/eJJktJcf7MkVL9fPnVK60pfWyom+yzOyiYdtZhna5ZVEpj6YN
3+JSlF1HlZy0ioTJhalqZVHC9/k7EfGmsENOy73/aX+B/GAeqKYa9kIM3ZyM/npVvaWyNg0lGwNl
K/aoQ//ehDDxx0abso56G7r0h8WEFkxIjhadSfA3WE2MUv2KWoUNqnQGQMmTbyNBtz13z2QPuv0V
DBse3DoHgGm3SxpNMPCmgDHHERhCNEi79JSffityCDZvDLD9QM+vU3Rkd3KG4YroN7yE1Gx9YWzj
LJ3g+N9zwonrQ7WT56mzzTbHz9TI4w2uDyuwbDVhOWJhrCZfvBjkf6CfmUNDMaSsRYKrmRFpaZ20
KOxLPTUc2PgQLk5yeUvUzTuCPHLuX7Yb10S7yxQaOGvKi3pjTL53JHcc9K23k+cDgLlsDn/bWtV/
pQpicj46Bw7fu5bMlcNr8BrRCdcFECNEuFihQAHn/wpKyig+NM26Q8wWJPu33f2nvHkIhPVoJCuK
dAtCo1g7vR6buZXO2aDey7/wh4H5iGq5Jk0r7ACdBX9XM1xmifALGn7Fzv7rUF6RKfbvFm+poDa+
R3Z7fGD0NpGmRDrW4arqytWnL9x5Dq/t5zugw94s0uQuQbJG7Hy2BRKclL/+8h/pdcg1tzTfO6ju
PmXR62GsBuKFmyIWrNfajxBObqi7yQ0gNM7/LOetGEkU67GMZGvJw3l+Z8dXXqF8Lgg5zOIBmJUu
vDQffXbajL6xX56oFFoCTGaN3YF9bMT5h+ccL/ZzJjQHzTQFy2Xh6L8UmyQ0m/8vuh8HLRCFQx0S
ct/+PFXbshjJsvOBn0rKJ9cE1Aa88JgHVjE/VmqhcEJBq5SfZtABp49PaPKEEHOe5edPJ00hdhWj
5HDbPMpzknb/oKcDTHWOr+TYEsut6HpfqNmYZ0tMBBQf9Bzs1ZbhYdGspnCGEW1U3F3B1SGM4WZj
CQLWXQPuAP1ruAARnVhY/ziAwBZu7fmUey+TyuXKbkS+Xk64cYoboVIJ+Qyi11ju1/oX0nx4M7/t
mdB2k159jAiO9PAwiS9xKA2195dfSiXa1Rpihvmrq6kE9aQaeq2qvNBuAt75X4zm1Z/ofLEpdCzN
jXqis22ga0SODv/2BtzjZ0K3ZwGQybgZaRBDed+y5klnZN8KgxLhnMtXvG65o5TdXe07wL9K8ex8
GEJYQFp3Nd13hVo7Vo5ZtDWDHL1k8GuWpZeq6atbGCNFBgveFswh1E9KgToCT0aybTZNyA2sEwCv
D/p+9Vn/NoIW6MiXpZCjDNL/N3B9J1UEnL2rvaUPWztWKFYIQjF7YFWbq9hv+rE5/u7T4/bAnO8C
8y27q6CKGIuatl7M2Y0iQ9TksGnyz9+G4UKg86D+IpyJRzTR4LN9sxufmtNriM6za/CfL1YXTeBq
1D77A4OxWnFaNK/FlHe5ssw0r6vtYGiuK+xYiA+IQ3FMscWSEaQDOr7k1Itw6L77/xnGoZeBr7Cc
UbFhG5RAvZYrMMVEAFxfwiiYnWmLZGO82igGTIqQia/08HFjsCrCoGMKfA0HCI4Aer3XTVw5Uhz5
+ynCY5EiWV4XwFILDJvrUGaCA30P41CDV+ij+xjrjs10TL0/VoWLbt59onyPk8Y3iv+gLuaUPvK0
5rgJYrikEdJVTx/HsV/3WcBkYBL6fyAoJQhUcvklLi71JocyHFi4SK04SlzX2Q93HHVPaCfF7TM5
rn0/ar1atdKLowQA0PFw5uaPqivHZag2pobiXf6CITmPr0Twnv+fKG87Uno2vJV9UYhWbtangnkX
54EeVFsAAgJ5uqqacBxm50g9TZI3/Cl9P9oyoxWDvZIQOAR47Zv6NRp7gh5B98LSJNz3jL15OnRv
FifbEcaqAf9XgK76FkJ/jL5jMrQgAcj+A1kt49WXS0JF7X3nDpCWeudCDXsuS7zgAMyA3Ym3kLtl
a31fwvboKAU/l37zGyG0kl7uBdYabvVY+b7SBgLiHv/Wh+XGY6guKs74n7C+KIaZi90UMpO6ELoL
CBXkbi/GiX0XwQBJwIt4tRY8L0GDOJ0vC2WQBzHyueZXMKwnf3+q9Dqa41A2KImg5je3W/qHa+TX
uI1NKT+P8MpHz12UYxwfnifYZyrZ+8b2LGHqDQS62nFbx9l20FCBkA7PNppoONixcnAHjRQIJtOU
++cBpNs3ui9DEVgeBx5dKQ5Wv/Ixghr/zLJ3to1r/5QxoHYmkw/HqhwNIqH3AQ54dAzocfqfe3v2
mS7npJqyZm24oSHlAazUhNPLFE0dZ81DN2vAY1mC8elb2VmPeqo8McsfR3u1/MVr2psYZkDLNmmO
cgLFYsHLeg1ZQYruu4AbL9J2iiUKnmY3nwy8MAuiBsh/VVtj3lE9iPzrDDeuCYIF5/XJ3NmN9JvR
NjWtdjiffrTtPmJGn7GonUie2VdrAJK7pSyjph1gtyt0L4Q6b/AG74fAryUGyZ+CtLw3pUD6qlGM
lYWcAhL3ujFXZDjQq0fUC8TxQlJLHjVxj+jyCZRjBZ0o8MsWGPUXjuL3C2hPfZqsUHTjw18ongpr
AhzlbBfh0ZfIdzKch07eCOjN5fQ3GRdc+0bRJJvB33tYiZ+P8IOreYw+p3l+vuIUDUFphRISjgm9
1FMZm1dXAD0FOypughT+Btn0B7iRMaHVGkmfJ1KwStk90/wrC74Iha4J9y3F127yq2eMCoAqNc2E
fp3q3i2uCv1L1GMvP/ufYPPXgSDKGB3X3pLUXzpuoyC1y7IZgLMdP9Hpuk6bc9vp3ZDPSL61F5HR
5mSNgZBR2Mg+5j8sGNa7ptVyzS1sVac9SybkgcKEhbBAcq4ST6GkwH92N+SSGCjL0IK5ryoz/JIX
XkXvwo/9hX1qDyrtaVUtfIhsFgTJlxQyIXjhlY1a265H8EmToi77u5PK8ktfwbo6m6QevwGCqKrJ
hyatkfSUTRbMriljhDyRS1U=
`protect end_protected
