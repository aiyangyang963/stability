-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tSec9jzCiM4o0OZP7HwaTSlpfVi5wUe8axUaTiPaSN+cm3H/QarHVnkwzf15qAMvbdAzn5g89N9s
YXtmEWFitSXofiVQB4R/6Kd8Iq5CWvnBYtS/BFF65vDWnMq9gpxtrz3EU4I3FanmfkH48+Gf/fyV
PQikVrF7oMRR/r5Qf6ZMBNdOPrCoq9YwVnPi3YATV/EdruL7gv9cY+Mtiu/iK+6VarHTunqoxP0Y
D8I711GP4qNcCZd/Kgnggw60sE9Tg8v273lBRJ/WruFnTSSARuX6u83MN3XBhCPRQ9sLt7foXMT/
YxxV/AVHwjR43V3h/DPLnETXkTmgcTal3j60fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3680)
`protect data_block
6CdiFJSgkgmlC3uSVziRxnr/f4XyceiLt0AYoDeZ03JxmVbMZyp+dAmYIygxEScTT2ZXYefyiEtR
v/DxKD7Z+INbhN28l0+99NjwLe9T8uYNWUjhbdDXqLq5JhZuxtKFMf53qojZpQCjbdlFLwuYmG1j
rn/S9bWGNcAeETRsPuE6yzoSBVvASGRCyjYFFi/v3HdpXn1bsBEMTxkcKcTdaFLq9j4RSJ5mx2J/
bFzlO5OF+xOO+Uw36KG6Ymp8s3WGnP6B5ci3STovuNyZQ/7CQ3PqmbjDVkY7JGVc2qBKvqHTgplE
0bk4l/CiNKL5AdsnFwjwZNNUwO4pG9Z+Qi5kiwxY4i0jx19BHRRMJKEzug+I1UDBU2NtdzBsdRmZ
FUeTMu1Swh9LsBDPcQUTvTqtTvN1Ja52138SYe6RMWyiNK0zX+YBMr7L05paR4r4iPC78eSwlc6i
smWKLdPZIDLZtDMKk0P5rVJFM2c9BGOHyQriOSC0ry7ipUAhldBOCOOr3fEaJc0Rthxmrfca+K8V
Ys9MFQ93bFP1x06VMChLo/MPATm5HLAo+DsWyIY1pxdWqPTGgphEXh41rZB/blT7urP3npbIpEHR
sD4OVSXGN92Vwz58SWmlnT1Ja9cCuoK2hBy39ZgdSDv37rADmeFgDfH45RRd/F8nzCGVl9KlDN65
U27KZkDDeBu9irLcn9WYJAuUmb9hfZUYImCLohzv4bxOpCOvUzV+scbY8HNAgn0ZHTU8pCyo+4AK
1aTF/qf0fLUxU46mVKgzVfAxuMY0lYG8VWdGgsoe8kXKdeVBS6XS8RfV1ZkZcO9IqfUY3/6Hdufl
l9Ed8jg3FFhVr64aJ4CckCW6fXXBhRa27es1aaMs9mWmovfIt4ak/zqW9iWaAP4maSw6QMFgVFs4
oudmdb2vGi1hKOIObEOrWF6mnhk3L1Hb/QdYBUiGS1V04eV9lcPCZzoe4bnl7Hwm/rpkFR6zDc5N
4awwdKCO2YfvBI+N+rPatbnDhDDJNQrkIdKeeGYLyNDezlNYkCunv3nQZc59DD2UfjZKXrJLHPHC
HwFFuTB+avjsOrUsrqalXjDZg1y83q+6ls6gC/c2SgPmxItnOUG2f7+tM71mtKU9d+3CqfdJ/buP
SBUtGVX3HCSDz54TavbeCEKM2a4InNNaeo/ZZCuonQWStcOvW6puF0WbQVoqOA+e8Bqr7HKBA4/4
PWCrOZ6XLtYDT9yGK/SyIOh8g3I0L4OFL5hMeCCipOOpclEdeVarBtAz4HU0MrjvRkENCKXLLUEs
E3e9HAnLxPwSHSGC13Wj2B8ktE/5h6DNJAilXdAf2XLj7tZY0Eq7BjLH84XztVq935eJCqA4sKAo
k3DXmzBwpVP++7R5JMCcZFRV6dpfn3aLdi9quv4jeWl3SAYr2Wab8y7po9IYmSrAIz/LyDi3nqpR
sklT/AN8+rqom+tQA/fml10SYWfh0RvV4ZptWJlhNnIqkjR0jbEghkM6g/OTraDdBLfF9AZxjyKz
iCWj9rKGsTCiGOZjBSidR3S6mTfKOYpy7848/ViPOLjw7at5Ei6ClfgME6k1U4QUWQFqmw4Wz+gJ
+N0NSaSbSTKRdUvyPle8h8iOYOPi/iFR5SIFskbn+z5TAFPAsxypmUDK5oiROnPr/Sy55NHjOajJ
f81tuSF0HErHiA/PtBd9K1ehuQ3ObSzVuQLepI5nYVnFuGK4/b86T51jxjeVGV2PKCKgw1/CGMNn
tRqq5nbppgvGx/5JIgsZ+CAurkiuW2+t2egw8xx+HzP3iP+OcNL/siJijWcNgAb5CmnB+UyhHHix
2hRmj43xsKpX17i7R3obTuFf+SDWZqd3vTy4Dm2sO2okEPpHJcU3D1VIn3OmnnXjyEGN5HEbSLDX
BMWIzcX0D0QdeknYu+l7yKD76ejfu3LpH/xpzWWbpO95yexKe1kD1ZMDCwRkXsU5jBuP40QFRKdw
fdxBga23ZfnpTGFiCsZ836ataZlMqYWShlmrk9XKKZc4WqesYQDnrvLCTzUYLbwy63jKw6rlKJsg
1uwSbgyD/6GytwkII+VGCsZjrR/jmd4WXDx4Lj9ADrnu13HH7itz4XAKDLtmHEaUpq6IHtq1mwf2
zmxk6l/lSU9A/dh8b+SG6ZEfBGFyrM9K7ovKaMRTBk4nApC8zycVkjVt+iXMMIxKxv+vsMUWQ8cn
kVsCef2o0O1wd491+3XCMK440PRtfUrY02S6wB7Lmao9ahxfqnYsRnT1H0Ks5BKHhHTLNrkLIeU9
0nPd//0bw7M4RNF9j8+SQgqQIF/DdPWXrV3ytg/jJIlrrLPD+hk0KZcAu1utVf0giIrqU8MKaR5E
PCKQMu/VSfqNjhXUNy4MkY0cEbQwcoX2bG1wXk3W2ePuWwA6exmKzCbktbslhBnntqfvJgDKxqMa
k8ptlaTPcRSWPwnQxOfeavJvFxLb4EgVbHfi6jYtLN5IWof4FPN/GsAiaOySrhBrxdWztoZWJFIl
AGH6yyla46JwOReK6eQu+cS0Avr0uofMif1JZSFTLnonj3E9Guv9+TROnZunogL2vAZcwm4cU+j9
y2xYnMwJu8xfDJcnm+XpduhNYMoDuBVyH66mh7BrQXfISwuxnald4/cLEBdWvcak7DGPLlWVDmKO
G0X7iNEuU1271c/VX+mUgFlPQn72YW2484k6nRilHVDi1FDuTxlzq/DnG5CaCeYUmn36oOOGVm0W
x/f47XC923jgSRcwyX4npKCuKeRFWwAw8SGn+Y6gyRYtmq5saTUdDz+rAA4phXwb5B23i0NOyXSB
1hkWwYL74MJbWn4PCv+FY4O8AmmC0VinKSirlMC7mCPS4lIBH+fFKEdy/002VBmLmTSthNaOvreY
Oi1nF02hhDWCE4LSNIUK5soiKMXrBHY7HBEsszDZw801/DWVgbZBDJKjPvysdHrCi1+tq496Eyws
TBWfYjvf/sMKxZlkyQHwkEamUwLKq9KEK51VKnZhZLzlD+NkEfsCjSISSh2MvBDmjgRSjmDfijBw
fRShmhDoc6gagKd5cFiJORYGWMh1Omso0CC6xo+scpdgClYCRl51KQeBxSl29fdHcJGyYyfC+s6j
18RKQ06ubaMEmyqlKNAzWPDly1ZhBOErCiOaE9HbYPwVHd0/xop53Be3/GQGhErSZShz7hhBg1J+
8ZJYrQ/gdcsa+j5r5QOjHAyF0bfNQ4X+PEQKIMrgtKt0bHdu1o7SQyN/3Fuh1NPx4XdGttGY77Kk
6bTVmwXgNmDdVMKAg4SSFkmFxrBkBfy2xDLfCmg051i+8JPkahH8NA2FQV15rP099vJ72TL1cWpG
BDCs/oz23tw9FTYfGbO+3EOQazt6g2lSFDQoVudgF+ZuJnv/VAtdLvBmXC3bR0Pk1zJpRIrP2/ez
M680s+c/tqJEvNqUWzxQgTe83k18pnw6Uewy24YxZwVUxGJK05blto64qUewi1psfyhNocQiJzfR
eFi8EphdASfiXeQG5NChFatGPiJY08ExBBlshGCQDJavUaO3QNt4W1AWRSuup/h7hPrG/yE8ywxn
8Hi1tcXyytHg64qas2TqcUj8fQ+HrgIi7XdhTpvssQd7BzVxLzEreKy6E1fG82Qag5Sxwz8WTH8b
pwNFQcPfaGTfyDESPCTZUreo2gYiXHvqPqekXOyMX2kep0g1PLJSFH4ZAsjfXZOCf/83NVYr3B9X
jNmOQ6NEQaCuHADtmwlvJblAVpIwU279TQ9pvE/RNtoaEXS6NfDUJV/22eSrZS2e9TyvdNEkk0OV
haeEfwl4bq5Qnn32+qaWBHdTklLiKFEjPeM96a3fPhDoAe7lmjGUWj4mk3a5KkBvTUQlxhmTZXrZ
fFvzr4tF86M8NqJgTEi2UkT12tFynxAM7O1OPC0+MXAI7/80bnb3RUbWgEDK9Qdd8XCtQrwzXkCv
9FVjTL5fOoWolyObihUaeM9clmvwMZUoaY2me6NXCS12JxYRfW7xB8N1DBlbmtObf/qzfa2dRA76
gDM8cERBUDNuC3jsNcycbl3NKcELgHUdkK8saAYzu3m8ujvkIkP0JeQvcZM+9GRNyYzeO8QTzFL2
o9/YqJmqIh5bd1T/tSEDYaHT0Qvkmluz50m8aFMod6Rag5QJ8i63xkgK4CF1q+IVdxWUXoWlSqM2
jvdQbDIE1bq17GZWPR2zLqg0HdBAXY56epiBpmxG6lJPzr2zK6ApNGozfaNk9uAwI7R2iru7RGoO
r3NlEgv2xtq7QmJ4QtGyBwj77HQzCPk3CeSBLvlSQlzR/z0MmYv0wiEQb7IklbR8FBihsHiycqFA
6tuaPre48zBkAGKILIFlqICCKChzUV0gNMQTU8MVr9czPF2dWgaaPLO70/laWCpNH3qhplDFCVGv
UCnJtQIJBJ9aNLST52ipeF4PlkyYIZXJKNAaFYERlRScgmYwkUAwCLzHOhdJ36zY/+j+SfLdxhI4
Q8xeFZ1k91eMk2Camxuhi5ChhxuKdHRJElN8oc3qUCNG3Yjkmn+mWMNH+T1HQ+JXgrbddB0AIPW9
wFsNeOTptAoMvaPFYxLVHUunQH7QFtvQ8JcZ/YaT6sKkd1zQAUaptEShvQZPvR0/Fm2tOwmqso4m
ZCNHyNh0qkCusuPtmqK2KP67Fm3k0MUazATkRKVrt50MTOXDJklSuqlMCrIKuCGHeNFRO4nyLuqN
9QR3g75UzQbe2pL5S5ooI2vUYqybIrehoAjRFYXr1aTyeXOZ61X0zPAHUMCnJxHeP1K3C0g8F40I
+ZaDdoTzHvq2QwEnAibhp98//1hZ+qCJpi6WdZ4wecclNqN0SpHZjo8eh29MuWbnA3fJuRH+Z08M
KgQlKFdsS9DWzg3TdrmMcI4PWdXKHqXIO/LGwhNfrvs=
`protect end_protected
