-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
isK1KTKVX3SLT4hAxIJew+qdvXhZMhfOR15mUz46rUPa9nHGc4daJHeRIwPiuJAsCnRic04Ys7KN
p5/zMCyC19S6KrdbCwzugc/hFcW8tLbzX5S+P0af6RMN8xtAAn78c5QNpS1Uti8nwPGB99Fpn6N6
YC/ddD/9WPoWSBrfYRdAu8sd4BsRnetZp/K+mw//RRA304ewYMhVWqquEli1wai/toLidFTm9Tt6
Gd8yePeYeXXHJ+Pgj59LKzKbcGsSoToX9vKgbMXsGviMgKjVFpCz1f8Em6zvIwWsxXZ5p1d7IyTt
qYWAp0Ajsa/kC2XNcqmt8dejQuF6llaSBihO0g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
CXCVGuOOO04ChoG3+ePByhVvlN2kY5cev+wo2GsVDPjBmaMjNBB9EheYg08K2R9Q8jlpKdKEsz00
lAD7XS5Ld8OYW/ANOgiqDukCO7WSlL2FNRKhDHO7LVpDCLTyvWUsBKCur8UIeOB4XQsZZJRhbvTm
x6K9RU30IckypRlL3SELJJqQJKxcIcVaATBsm7iOySFwHImPnJqO8s1Af4SjhuKXsZShaS3YFraD
qxgmK5qjPvZOc20aHJBh8iOTDnAWD8jrI2MALaXLz70rUKKDQhLWSJeAL7Hg0L5OFhyJY0+1xpy+
5kpeFF99qSI4/0iOrydgEGXgO7agirHHs8PDWEJNi10yP1TyWb6e9zQHum67rhHeVmONyWznrFaT
65zUYcqKbnzygHbE1re4Q+IbiADN5rFGPY3hETLOqWnz+WXNgrkhv8QvXL5nPqt0r+HDHvZptmk8
hSub0ApKYiqThGj0R1Igx8E5nLV9QsQMvyxc/+sveYZ08kCQqwJwpjH/IE4q9fCDnhxGlTOklQ/i
474bmyaehQM28UDj1aeByTv2ql0am/U+UVmgdvPl24OrMmGPz0ZRZlr1xDNyFBuWwzd0XFVbO0rP
HkRLtkk2WI4uG3gBw5YYKj5Y4yzpr0+/vcs1yErS37ApABLrRQC5bQN/HieOuBHw8sJbxEwnfyF2
Y+HdAduehZylfq3pv3f34MO4fZo1RjZ9U9vJpuv9FExwLXXh4RdxQ8Np3AO0GF+L3XaPKwvxGSiQ
8c65DwQioIHEkR/iYGb5ASNjVXsr6xh8zU3EogvJm8/OhA1lef/AjwH+KVB/Rxbc+GCYNEwGRZ6j
9Jg4L1jFMybCw6SBvIEpIjQOhwI02q/4bism1VWCqGYZBj7KRF1g4qiTi0g0yAoJeT5x/Br2gKu2
PDxajGFR01KwU51JFuHMXZmh4COAUw7YUtRq7SDH3MPDyYkGw0VdmyFbLFU2uWQfpwz8xFn4hJvu
ptC1sUXFD/XOoQ3JDvB4QVHMuQXjx8p/iTM+1FGZchmnS7hlj/2Bllhrf6/UAMHMmaYspEJEBBMn
1GRu+psyrOWISwcguf1/1p4OfDMEifp3KYr7XNttPeBJFNdyd3a1fu3lwyEQppgKRdL4qpZ6n1c8
Yj1ZxOBeynJYZeda9UPNIuwv/imkUqTiWiy1rYJeS88+NQV4RFCuHi0mWB3u1Xcep98Ci5cord/B
uhOh34walwyzw2IUv8ZfhKvHE/gL3rKEdoY16sEIkbDMnwiBE05gaynXN6/ipHJvpZKSZ+xuoUEL
QNvijK8orwo3iKX8pfzNXSxc3XNmT3F2fyNeakR+o+bCWeVTDQHaAnAk7ewsUbhVErSfTHSzkKlP
X3O3hdMBLuZHb1aLnKdhsEPH+B5g/getB8Fx9Lpu1D3n+yGooWuSpTTaiJJcpTjab5hfcuRFtmIj
jVJzyVdwqXd+Q/YRNXxniGtqcSrd4o/cLzHD9rcDLqbzy35FdQ4AeRYTMbNPjvOtrNzyeODSJy1U
1mVD37KTv3E0R4bcI+k5SWxkft8To5D5EbWldHuVmhpFnNWlzG9Rmc3ZOwEIm0i0ckt0MgIJfj6E
4uSqZ3H8wgJeiVJVP8KxsK7qXrdgETwR5/NOIorL5Nhsga52aQvXrrorJr7qh2kk3pUEwnD/RG5t
fLuLRmoSRqH2F/We1WXGsr6d6PjUEu8KY7ogc0wH6j1MbgfLtt3AEQZj+tvkcXx5ZfPuFswVHDY4
OpoSxR1jzoxrDRkAo8qTniVEitmsE7XZzYH57k5VJzD4NdKYVjckjhhxa0Pk/n6USBaaIXdN7wW2
GfubV6ZV8scflHipBF/oaI9G8vPMyTCsQRFWVLS7BUsKh+PbSNhCAbaxbPfR8Zqn7t+XX/xLXkiF
/lPGma3FWLG+ww5snZHZluNT5clVsErd1EkCJkJa5p3UQUMBdrnf7otQ+XroB4L1yTeb2AD7X0oT
GIOzGEuoQ8hw+ggPtsOHi3j+YZr/SAdzFWdRCWT/bpX56wXwUO3mD4pPsbaiZ0NUZtb7OvcScSkH
nAmFHKb3SkcxsmScEGEpIczvftyr/D6KAWl2LRZcIZrUMqX5BXKpmqjk2m61AMG++/7Ab4+TVkSu
k9KkiRXL6p8a8bxnR1KmoVKtmmneM2nt1R9kDfO5Y4+LtGTofWfufCAho1AMt8ewjpKlxhzCI8yH
UC9+UOwo8JUBzGvrSDVzQT1BTzV0Z9/HI6zqpzHGBxt4jYxShiGRnLNIm7Zps8E8eOOJzS3WhUFx
mi0gYLNX+A8XSa6Uc6bUKHy4wbLMtJr2GhHNMNSRa7b8acaidQWb7RhXuZEFE2+2OkhKpQj+NVjT
4ncb6AblOBQSZ9zUMbrYCeLRof7FE2xMGPTRsqarWV0MOGy9kakhd62wFRC+ORXPwVp28tGbRdX7
Qidu1BjapCMI3CT6btiKzx4uObiNF9BeEb7UZq58J+34PTEEmrtOCmHRx73RIdH2ZZuEYG+4ZGcX
Aso/H8bCflR8Y0y3Sp/mULylThh02APOVod4HIGF36bue2chr+/slvQcTX+eZg70Wk8semqp/khq
y4CfmJbwj2jXvpIW6g0cmk+Fg3AYYSmPHv8ZKRIiGFAXvzi1wfhBmLY3tfxWBdT1JWwikqdz0hK9
sD/cemN1LZzE6jME24SpWouUqYSzwc3l8RohG4vg5fb+r4nNnbC4mjKzmhMe8boF8gJ21z2+h1Oe
n5Go7XNq6FFvYNcARpsxZsdDSz4u0wWfIbfbYvTvy5dxRd7P9WqyIzOxBtuzsMp/kQ5QiO18eerY
KQU3h0NMqmWiEQ7Q5c/dzxSVq5iljhvgknk4yomg/MRv17++/eWUUp/oqNDEL/7EN6naNJziofIk
hAYj6AqFuZjTVx1n1FXxTvxUI5ZreTRCX7DY+7blkYhE2jTX+buCq1j+JNQoLlKGYx7aZNT32tma
UgCjcMH8EFC+krN20NzFPAxF4RQ12wOxXsfP9UNU7GfLhhOJHUkXRTvMzVCfZ61oZn6rFVv+Xyuk
WZJYgJ1PjZyxigA5mcODFYiWDoaKqdnCtKPp0LtG5SnkMuQgUMY8+XOcE9DjQx3bK+Gz90FTFRXx
ucM6BDU8+P/CiTvNVGL+wXXcYQJJ4k8nrJjSJFzSdxC3C63/vvFPnzIS3VCxsA5dM89dqnPfKB4g
8O15v0p9vyTsvTtQ/pjsD5RGS3DWkagQyjyoyOSzg0lJnQ+xjOmruso7Ug25E166sZnUrYVuRkYR
mGnkIrWx3YR0W7RVcOi6SFtq2g69oaXhzWWbqj4Q9HzNFSQfPDqjPiq7mUOvEigs0TRGe/GZpJc/
Z0vm9427jvP1gVVpvl7E6mh4rYqUT2doVkKV8zcGna78u/TJwsm9nYG4awAIyFbeF7EPYOpI/x2d
+kgkWh1IOJoUQ7pez/GYLs19yoWmgVEdL58XPd5QWZkKY3zQR9Vlj6c9HsfGENPQz4N50ReHp10E
pHwPq4SPA1H2Raoog+tazNlxtGufCnXyrgUFFtFbn2Ld8kZVZDmLx3jl5SAdi76qNdS6jlf3ecJz
9J9HXsq7vaLK/5no67QU9Q1y33Nf00iOoyqIUYCEjTpDJ7xOt9dQZZmZ+YESimJRdeO00pt3yhmX
6qVranNoZyiTGI8cFjq8y9ITzEbD2qIj6KkLMC/Z80nxmVNnvvvtnOpBZtvApaqBH7b8wpkrOX5R
+qbQPjWW6G1p3fWFiG0A+g7I/x4LchglFD6kHGYnabmjfsJ9Hr0ypcE3EvCdV386VHWBOoONTt9h
DHYIl2OfCZiMsGNgSDPrj9zzNxZ7nvTRPBgnp3qe4vep3nv1M89QUNtfQvgAuzRTtsO+vFsXAaso
qA10aA2ruDGmeyHqW3iGNSSl3GV/AWcfixPvqFbZa2moz4BlliKoXwpE1E6ldezNLLK6US+JdVlh
N0Lhu09MJQvk56eI2krDqTS7EuyLx4XMSFebh9ZYdhCRyBjhU/nt5aBxOgOPNB1yjs2SGmK2TNaP
eWp9lNv7NkakSS1w1T7P6B19G/krX0CXUUZZTpZdKb4q1Tw0s1cpNVxvTtIZijfFTHWk75ZqQmZa
g/IteRPAYH0IUWnHyijoGn2AQJ4yqw5aOkAfOeWK7igPg5DsSh2iKflLTBKjdq3hCxTKd6Kzb5BD
qRgVzii4D4nsuiT37yc10RId/vRYUsv3MkOSdBs48GEFD8TNPgq6/PVCbHMd4/KU37sYrolmgTHa
/3mabX+WwzU1JPj9P6CCuh9N0CrP7kdXaj7n4sx+SEFu6Z2YECGrdEouav67Wld01HEUQ73Hge2I
mufUF1Vuz1ME1B9y8pkA6KcocTramibdIiT/2ageeONQa+Y1heg3kj5WFHXECANQJ57b05OaJfgN
VKVSsitcxE8UJ5djwABj2ELPIkoK8wHuhiEV9lGcYzBto29hQU0umGe7H4tf8nlcAsKJv7pSGhRI
S1aqbyPbb6GGQew9Kc5qHb0BIY3/XTYK1JY2iQ1kSPOouBOLxmWM4pkkAP5AwMzhns/McCmuAtBv
miLE6LM2nmUpJ6khtm/SozT+VptNcCVRJqy3G9pJ3HK0+lUmaSGIQxAnkNg/4+/+zi2lVWDmrZXo
UJtEEym/vppHfQCT59aHo74v56SWbek/Dw0r4wHZA4gm9Ov91KRXAPvLTsro2azniIWhWvcWs/zR
HPP/IKz9vyUTBKu1+e8VOfO+nMJAtR2EI+bclZhZE+HeHUSXXhqkkN8YqBFFoo3WwHXR+W80DjtK
udAUoz23y3Mnd+4PFoDkhwRcZmuchnyVeFseooLAKC5PL9rag2oANv7a5st7NcAFu3kP8ymHATnP
p3pKaj+CZjy/M1PSaqdZso+cll8diyPDqy2KYcGx15HPFOAFmnL6GhPFrdUnCoSmkkL3z/UJZzBz
CtdD6bIsb1TkEK/+fZXe5poIf1TgNmH3mO6UhWrPxUy4GbbR7If/gqjIrS8YWJlKDrfjXgbmRgVv
5guD4IoHA75jW2b3cGrDqKebuPh4e/BfRoYnBouH1UaOA+Qhdsj0YY2STVsu2RuqR1ADbAV5EXIi
xvuK4/pCNq4Yj3uIGZZA+MNyLgTmxREJqBzlWZCcAroyThhwlDyW4N3SES2+hSADbcBVemZmGKig
aSfZFCwfQfy7Gm/r3mJ2n3dnNrWy7bFted7Xe6U3d3aqYPXSZX3aBkjRV5Ua9nfCEh4bCGDYEng/
XnsdUerLIHNrfYMzmu90WOtgH9hJY36Cee2do6S5dMhhPj9MxjzTMLmJaTak1c82oQe1GDJWd3cz
kETO68T8dnjedpO5tdr3nrW3xn5StCfw39DdFUIyvparRgq4He1urEmPtePt9bSS+dzZazN7wynu
Q68KB7fsMzv6d8Bdpasu6TiUcstA4hxSnh29DQ7+XpFoe2oMnqE0zsfR15aidVyb4f01zLWar73t
ZzARAvRpmttEmrgVaEYKn5dgz/iLDOsbIsJ3hBZpugtEQ8TcHvF0BVYUr5ERwx3gaW8LeSyymUWZ
vvFsu2mjYZautmTvZV2zlbQAt6ed+zjuAv3qjEYLkYks5SxI6lJZR5opBodgrDCTiv9pxcjcYe1L
ZewbG3kecyc+sTlziId3qQSYreKRjvrZOjywBxMo3mGfSxJ6nUbfE0Z2EluwZcr2BxCYrdUsa9Fc
YZiTOPfdfLVmbBW/rLeHtRMYWaKmjjWBwZb+Y/q9w/Qf62XH36VT9PYkNtHu3EIb+/aum6fc34OG
VCndpDIi9cKS2gTliD3K4kZ2s0SrVTVqS+66OWRbLyDwKbbRoOKSaBsYDfiBgnOKGFOieV+tT3HV
z55aXz8QOdzQRLsDFvI2k9MKoIc+m2L/axlnrB4Me2yf2rwP7oSNQApxOyfJ2VEX0B/hta2j/19k
YfM3kAsYkREQwH/mjM+ybn0ShAtvqgokmnYJmNtgMPUS0YU4nVF4x84UDudv+1dw+/IFEJLXZTLG
r89Xv4S/T1oL/b8LJWwUo8s153zTYXCXuC87hSK2evPwsFHvOPzwBZOBBvhIeMF9kmseOoIw/1t8
cEUD7g5MxY/RzegQPLX67UeBJJeuNNTGu/CUgPDgX1srHkueLvvUOIlbm5HgJIavMXxy+CBPwp7O
2AGgUKON3kwYbeyUtdbK+g+iYvs5snJEOeZmqcLPLallmFat8UO8XAyxp0j/GNE8WvCvAHsOohF0
pu6HyL47fRUJSZqMaIl/9Ixd4485J/X/QkRjEonmiyaBJFZwQhSBFg1Q+qVYwHt5MdndzWSfUUj+
NK69ed7172RIqIxWTDZo/ylO737/HK6y8pNDgUq8RqV9FFJItdOxIf3j+aXx6yBakgT4Cr65d/3i
AKlhOBhLU9Oxij2xX+1q+qAlB7ww0hpBmRMp+Zgj2fFMG70okoVCLvJ20Ff7YYhtZRoO0fB7i/+i
myNZ+c/0ryunNOMq38mGQ349RGScBYpR+XqpaZOAGM0bpoXNC2Fcwsx13cgQL7z/ChkW2p7l8Zj+
RP/j71IRJUiQrTmUONI+3xnWIsDk2Yz+6uXbkDCmLZeyl9gVlqXBtDTWh1MjSk3F0VoPqhZTiRa5
HtixL3ZXr9B/elsvjYEPWAWM5WF953dq/wgjfsmc+dvgvd61gxMIAxoVzdDGxt92xUntbQa3ffxn
TLMng/GUyPXnpeNwAktbbL5K1Z2kivK3RPtqLrNyKEC30wqQIH4NWIuAvrzhQRY8icPdv+ef/FyR
65biIUb3HAGQrY81NIK4qcBsaA9vxMpLdGsIb6T4XhNWu3v0dvvTA53uIsU94vmYkgSjAp6/nGcY
cIjODAEmu2eHBefo+xDbomqJ03trla3qcbPCvTwss/xs/BDPr/fv32/luugW59f5+NUcgAQvkr7r
Zar9rExPT3PNK6U36rkvj4m26MN0r3VRBuMQgugQOQKeZxYPPs3sGVqb+ecbmLbZPe9/Dqh8unY7
lQ1qgfrvXIi6gGvNxlfCC5Qjsz6PaiKqUtHNgvCfjlCP0BpFGNUfKUcl6WOd9pYTZDuePDma4fwh
vKFsFzimxmp48ZTxF/SORQaHpGD0Z7+qfU1OE8UHXYnbMW2HFPuh1jtn/t+Oc0HGRnhRuJj1+Pev
YxsnV5/TLLkYFkKpwV58m6k7L0pnOLMHl88BU8oOmok8i7+tpx+5/fBgrxDl1sQlPRyoSchQo5r1
+YW/yWxmA6AZOEkNu3dgGcjWOE+5KlOSE5hCF8FBUZL6a4/gt6pWHApeZzpJTDZXx0uVxUZyKEH1
TZgQna9SNt+mNrMsGs6XUyrA7MIKA4il9gr5+WZABCwMYTG4q2MTYxqedSyZoyr5s6rTZccK48a7
nhUXnQ+29HLCer5vxbxxqdiMvq6DdimwreIx/8qEWBVvIekeElnWa06PZ7olLIlhakhINqhBs5+G
vPt5zaJ0aRsRPH5k+t6h06E3NO2ysQEDQ4w6Mg6BBc8OlDqgtWlQYWSDcB9yR9L4QbLxh4E5bmGO
OBBPOiYowpY547DK7Ttk6N+Qc42fICSwk+GHd+RRnTtyl0Z3bbOBZqpIrZqY/RwO/f23P94U6R08
UI2b8CKbTpqk97oYo1v3IQnlafiZqr1fFxEGPDej43Aexnh56cEz9u7Sy3pAx4mMxKQCKWLSWJAR
izscu0rKDI4g6GFW6a/BA6ufZ1voPNO4xK3zerEgxINaTRgjD6cjhu1WzHtSxq3DrE1cL3Uhj8tV
UGOxz9G1Y7Pk0Jelzk/6l06oyA8IVxdXReQOdF2tKoUztDIf+IP6iumbhUaHzh+pLieQGO0eeLWa
UMYc5hqN3ZAa6gX84HxoTkgWLPRI47a3izBn4RYQDlDKbiHH2OsjgqUxk29xWrONT++oj6VhRfnl
04IbT1w3LtuSD0u6x58Li8EIRlV4xvmFKk0pLjixQRJcT4oOMWz9rHAkbSm/Wn5+pdKRXl2ouXJy
INFRxBVprG1HMBsVSNgegblvzjOxTA0e2F8+jrMMZsrnWtYqgyePqygDWv26ITFgxc7R0dyE08fI
2NX9VVUUwlPFsdq6I1BvScZR5+4wRm/UHJoXp+ISBcL/k/GnaF9VCq4E8KxHvBU48o+/udyLU49A
VxnM0HkLQjfEpoUgZnPqgaKRXeByOGby6g25NdzIF4T2F1ZSV2Ojc04fGgcf++k9640H0hgLt3bZ
hp3gZsQnlyxvqy6O9Jdl2Yutv4xNC+AJZDdhtrjwMHqxdCIU1vVLnPrqFA5n6hLmj8vWzFFZdE/Z
utvuiXewBFhG6yeWhepKyPcSLRD22OW4Rcm5YRKZg+QFUfs2UjfMRlUkl0oKBZkiVxAKSjsI4eqD
VuVrGO8ft/pKaSjoJW7U36QTONldfB+eiMdren2esl7N5U6FE2TAOjY66J0tgZNj+lrVa2yCj8Um
YMrqQ0KS5aBRrVKsbymNv+8WQ7PUEhwYP2hisfzhb2Ar8IfxznZat0kcOcFZRU2WlVQxftZrIAjP
MBKUZjnFu7IcQ67DaXjBSk5xZpi1bf5uQVBUPpBn3L7jeh1cLdsQE2hNnKamBYU1WeV3w/QxB0zh
uaVKdm1TXkbLRENY+Ap5AGPxJoAHBceb2ntdRU7+AmUTTkdZMxYTak7XgXk9SBNxvzXr8QD9HRXC
wM77bZMMRzdzm8HtfQHHnUYFuQu2N7jOeNQ1JhlDcA6KqnfUV/IoECqs3wWhp7rXrxYF7OUFfSnN
a58rFsLS8V+WePdglu+hZBaC0vHTyHoiJ6WR4jDqWafyY0tjcnecPQz0qBBwyUyD6QpqE8oMQCXI
aNDzUMm8SotO+3nOirq2KIAlzeJMH64n6lHZOZzgHca2oLBjPNXdBdMj2VHhGM6aA+MQeCbh9e69
AzgwGaRFyEchOuMSA8yFvZUWIf0M5WgRPaq5VkxChOQqZN00akkz/pfiHd5X4Vjp4Qwk4kHD9Mv/
GRKdZ5MdvCgocB9JIQDih7As7pZ4nnsWsDC2ZEg2KnKNs6wv/F0gc/f/3ExPMcE1rvkaohjwryqN
qzIOQpVTZr5wUZRV8jUplxdxigchyAc1jGAd+nsLQPw7ZKxrIKDEkuJLTUTQKeGZPVVvehRtPjGF
StIl3sDNN1iNp9WipMmROyA0391YGUr5NxhkBKQ1KeM8+L8M2gVYopmFfp3xtwiI1N+1M+Gy56S9
V1RCmx2DfRqn62s6U51dKhvvEEI8My3Voo6FjkB7IqpdVPBCveUBmu3M5mE3VmkDkH1yTRdedYpJ
E+FGuXoyoLaByGT56z1uRZxl5ofFAhDPx0qlVPBxl3Zxg7e1k+fwJyisYFoF1B1MUUoAT5+iDFU9
kaEx3DU6deByS7+4+t31ZIx148D9PKDn9j3aYZ75Db2CQXWy46ikmhC/AdmkZVsKgQl14Zr9QdAe
kmn8YG7V2AIGDZYiCk4xW59MnAU95eIP1cmIuHK2U4WsrAW2N+kbuTm/2F94kMYFp/t3fW4A+Dxj
DbS9IeHgB0I0LiKEkubkyN+kD/tL8resiziQ8q3mBZEJRIHM/hF0VRUfox5bLDiR1GZdCsjeYcVe
BZ5ZubO9xCVBTbO4ZNeJOBH3QVLMFrZeslgxe2Gq7qM8OM4DUM9XMi9YSe85fj8HDjjZNfg4AK86
6eoE8OTBP2/1z56KG3/wxofXwsOtf7C49APnBXofv88UKnSKZx/SsXI1GYbvj/I6x+ZVh1GbpHWJ
naUKvbKTwl8r8J/AgEeWR2qTTrLAESL8RaCgeZLma91ald+bzbpjtvbecTKlkOb8xakbZ3XPW6Mp
1ds71ilMVqBgNj2+fo8qjMMg+x+5dnzPxAyGEqROkAMi6c4siFf0T/g3V6X1WxGWj3d6txNNus+5
g8vTbzW74N9tietEZ8ONhlHWN9bKpNXUpl/uzl/NN7PfqIQeuJVc4BHsQDoRcGgrJVCzrDVdM6Bf
xzorEPlS6MLEKyVDcUNXwfuASafVpHBU7i4C1Ae7ljNTWEP69lz/jgNRM9S+ZThT97LOFBYHpp6z
ZgSn+XhfR0KDuLZoadneULN7I4KPwMA/4HwbuNWIOBwybzzk//6w/dm64aLHC0mzZHYjUcBBGta0
u9IAZUG8+P9ipLUyrgQzVeoaFIpdoMVQdFDRVJpxqA8Gjcl1bqOnjuUddYif/Sc9YE6T4IQxKw8I
5ZutuMRnpyDl9jaUV9lPHpddkMjWPv/RUN9z1J+v3I8a24nYwbWHbCXqNWJ3BTgEzuRxHl9FltFz
i9FaIThdGSGdkFEgi0+r+hKBi/1QEkjhbx7DnX5+ahNkqlhmqlp7QUnXBJAtxXt7dkPfP5ZjzMfh
eZmzM2tzJ9An1cGXeJzS520aVMA4O59QJWKydU/9I0Ten7IcbYJ+xNN5e+VUNArFBobDb47N7HH4
cMEOImJJdfYzXag6uAoZVCIR9vEMzuIg2hZxP6uU8AISU9gre+Md6NmkUaZ44oU2eOBAmVLnYFUi
iTQ7mEK9E2xpdlQSNhjGRrUNcd6l3Lh+/MydzKN//tYHraNNF0OLQgLDAW6HMs2L4Qzf9SiDh2rK
fWYSjn5XfE43ouQYKPGM/IyNMDq+JyAnG9fMl4+yJz1mZx8YOwml6DtvIol/VOr9BKKq+XcXVRAU
kjUWQaH5BsQqLMHGr67bYd8pzlDrl+0PkNUaRyxiqX56uZ/g3UPqjMfxKN4Z3iW95wTaB5OMfnEs
tHJYB/dLMeqt9VCg0qaazXk25k6rA7oCUZ/bhLVwTsIrjPFEuU7wtBi56B4G/GciosKBwSw4SMDh
Lqk2q8JAwNPObcv11b4ZFGJo/1M5ul5MeZmDPrlG7FAI2k++voNwJRvZCMxjwulLmzo0Xmqpwuet
V1OdF+LZukP1Su9UAVLtSxATkDPLafQsNGRA6dkoeCjw48dyZ4myKZ7KFaUQmqeZV3L3kpYCGhIQ
iqIguCDCcLv4dMZSap0qOeewfFNI9skEJS5PYSn3ZaTmF2SJdaL21bej42bUJwnnbyDmRrnGvUw0
HYYYnBLcqDaZVg+ViTol/VQrNj7BCfec5WwAGeNhgrW3cXN2nxIIF2CpoPHNw1vHGm3qpu5ai+Jp
h94q8OLV0Y6+paT2uK33bVIuhDAX4lPyiUJBWAZqziCF3UNR0hRqZz8YOC+d4O//HiaHhhGZLu9i
q04p0Isv2kElcafx7UXVNb4AH1YIHNZ68iwBwA9S27atNyr19hCH0/oDHam122mTorbv/+1+CX1Z
N5cJCmTPutaAagshXNZtEOXgv5YiUrz4DuNl7a0oUGwYkPOcml26rwtaRYulkisSBnr8VBc/OnFD
ew+lAAJeCOHd5w9NimcWFhsMgo4o6tQLKt4lwD/JW3rytl3p9sJcxOwiVr6J0Vt3FfR/gyjrOsjc
0Diw1y3i7hYUKHvVpEX2XZR9CIOeWxBEDes46NsSMt/Z8k4lGk5cb3urr1b56BHzMW/dltLNPWHt
MsvAHFUUOjIacEfMXlWt5havLAauiLdgFGh4MC8Y3St4ga3QIJwG4gsjDXpqH5ZnZoiFyWDOxR5l
tSPyycv9NZD/ZgH8rer/EKoIYC/qS6MAZDuJdF3WQSZVlOZHb8ozW9Ls3A3/l8/F5c+Le2A9NEdg
UoguI6jmjfYMojLD5JoiEc0I064gTYkA+6cu1RiZNASwXQ8TMszqm4j6O2cCdrQLrVVw5K86SPPb
0sVaI+0grg9PCY1JxV8zY2q6cbsW33eiz6hI3/HO1DX02DDGhdaF9FrkIw/763dQ970iAnIRqwDM
jMNmt/da6S76RrIlzs7Uc77i88PlExrcB6+LSGy9YSMU4mQlD62nhBHd0PO8vmq3kPklTbxNlrXz
gfJGB8zXV4YIqH3+RtsmD5G9OqDKnKmtRM+Z5JQXLvSaWirZaueL9Udv0uCtEqhxmv0O0MA7d9fP
jIOzfMY+MgSul6fer416ge9Sr3K3zkg6Zd1rJ/YIKsUvOSxDuSiEbqfNtg1hdtAPTeAtQmoEVj/s
JfJ4xtrFyvP+S83d0cObba9iIht3gzefwm5BFNYiK9aKATfPWzeOV1xm9G1kUVSAnKzIX1xZAzZS
YtW+IP8kTTfS0GEupV5JDkyuXv33H3E3r1j7QALDd8hOBuKa2EEHPRR/KbXDPWbAxXUVh+EPXJhY
L7jEaL0D8ww5EGPBUkXw9xlt8MnH/Gunk5vvruDb+YusIYjJjIwqsqtZTi2mBxcmUt0O9mmC9LTf
meW6YdpTomf4RX5pIyUWfH1Lo8KmPSOKCHWMhfHffHcvrW4cfKkE4qn9QmJcMLNP2rGxqRN/zPDp
OpOm2Ih0PcKL9TSphxTCAA8o39yNk4MnlbKrOBbPCejLOyUvkMZSc8sry5LRbmSpk3Ol0cSBMSsK
lpwn3z55H24tcsTcUlrhT5fB5emIZzFIi4P4xtI/fNTOTGEk/j4a4PQP8vIiC4VVXgxTN5WP5hQt
gXmefONu9J1XpcV5S+5nHdq4lZ/vnfCkk7X/+bY2Pny71Ye5zgGT9Q47O4jGz1BmhTPdDJVvHDz2
niLZnlgrhzsNKSgxhxGChMIiputhZO2Uky2b8p1C1MN088vc64vjRiqtMaSdRZkuXEIgrfftEUr3
ZlanebbRtb/jxfeuNuyNoZgk8UBxf8FtSfGWgT9rsQV2s6YbMS5XEEPh1C/UnIQGd69encrafXVo
DqCEA1pIIDDq1UErh+KrH7T5FHsTp+4nv2aLfhqBpf3Cjtv/OzJ6Ga58XMt+9yHLqJ8lGM7G+BJ5
Hbsc3RlQXtq6xg/9/p9Y/OAAjFL8/BJbzu0nYsLfw+Na0F3xEgNQpv6Ay580RrvSzt4Gq72X8HpS
f1p77/FWOls9RhasSBHQ2iO0LfQA3Ok1DWvuyOzcr/XkoaXU8s7ppxStvIllbQd+1uj+2H18v0bi
mfiSX0b2o9BhjAetT4ZNoME9Dl9HJWLtGX0e4v6yeK4e3YjT4XogaP9vSnjsf39UkBAOeipY982a
myGPEGkb8gzROw6Xdi6eIMaJihdlc/VtndKxYMAbOeBL8h4rE3cxw0GpTC4vjDeQyQN5Czd34rXX
eNtR1t3Nb2eemforKGrtuhpOe9+06LhLyB6NRsOi15RxHGpxr895C41a0a4Ra9/HBIMCeoR26mcd
I4muvX3ANyMNNDHEXIaZIkd2oJMiXa85N5y6CYAtzJbhzWOGL7x+tna1aN8CxIIsuikmQ9t8ikyF
CG5hohhzL53rlJpsiDHV1xIIVGqw/wYJe3+gcYChOLJYRP5tzb2yu18QtTticUc0WQ5L4nUeJEN8
/Prtvuq5CiVZnq1llNehMCx0Np7R9cEqABddZWqQi85MqnmBuQXypZSrAtXrPx+EwICvMZYnj2ct
1KrkXNKNcWIsA/U6M/refn4DYXh6kY1Iwo41cOyrTL4t+pKbhyTbW+U7KlXSsNOG5NOoqDQreBOs
ZpNqkfAKThezqFrXuxtCuSW5IiM2ZAQwqpsShq7XQRtTxEeTI93Uf7ggeLsGdnstYSj/L3AijHFV
WMiDSIzx2Lrkjln8j5tnk/XIyj3ntbWrIorWkrldYdMTb8FbtyG3Iv2VIW6Fn54o+6GIHcEDJM2L
i3k/GJvv289cwoH+KlhBp+/B8l0CUGxfQS2Pii2GuP1UcoDsZhc5zFTvGwY6gKNfcHLcVBNIWyst
ISTYziuezEakqxzro8IXRyigUxHz1pi39ahAQ3YQ+dIeqsPWkEHM+BQqHLfjhJuSCQuAxgAuPeHW
9t4T9Fx0spkMI+z9+O0YKPj6tg/+/zo+IIBylPyiIJwHziuHxlYM4FIlRQBh7U3DTK7t73gqPmgG
X41rOQg/PzumwSOMGFEeyc6D6nWuutXTCdqdGck/IzKpL2JOqMtJ9AsvA0UpmWZRXj4T/wS3f66W
b3yWaafSIS/reF1l05mBkN1k77HS1/i671nkfLFhyR55o2pNzNixaAnkHh1CelykXJT8n5ypIxPP
qiz2xj/5T4d0tWXLhjlRnmN2SrcqKkddN4ElxU0RJOC2RCG/v86jAivabRCIvYTRT6NzOiUqmr8z
lz+ZyJXL8bZi2cyvsR8Fk9zVww5kmiJ21FshT86RKYX8boT1Z964K/+Uw+pI7duijq6QSEdM0Ad8
85GJbQzGfdD7ETJVQ25BpXMRxfAnfo83T3/AOxb+iVnLrf+OpWd1Sl/w5OooJCbbTrJO+yubpKrH
vR8Mg2DggmABDAtR5SwhwUNXU9mcqOLXR63NMsvReYK1Q9o1bbOHSDWg7blfVYhmYbyRsVS1ajfI
ZOjMVcCxPCyXI6Xgt6dE6U+9MPrdC4N9Tn6T/q/CmVcuTIF2k8ecFGWDcqOTuT6qoe3jRrbRSm0Y
/WS1X7sFhp5E4GtTZRImtKhrfTu7ez0xsjs+weKLih/RYwn9ufQIBg2UHimT1c5qfWKUFzGeNlFV
UxOm5/CvHReSbQFRXf1CcjTCvzztZnpksnB5oMJIbCZ4SYoEHOXl3qp/AbsMTZ2/6ZwadwuUMoRh
P7Q2uwj10deN13iYsW8pV5Tbjwqif3amEO82+DrDK0r19Hc1a0SNEZqUxzmUXavtGZ2dgeYbvglw
0K9pSB6Ab9qRb9gTE8lr6AFOc9UIB/7jwgyX9v33lHYlVqhU7ESS+WjgYrv1fKstlcqTUyPKtvHF
9QhgfDCQ/wDh+nNUlXRk7c8NFN98Ct+CcJtqMVpDZT9CB7H6oyysWijGp/MAIgdNYZc+wQ56Smjj
2z6ft5kNvSwRKniDDUHGBU5L+vhxzDQC5Ru2x4F5BCU0RrVXcJK0VI5B7oqaFf5+ZW1YVgsyKcXI
D2Kwt8dV3SGrdFkOLi+OPKRdsa0KqLeuzNTRX7klcgMJJgFkUNf+1jSy594Lwp8pWyL8Z/+6HZf5
gtsQbbNROq5VEjOSwMR6S+s1KqkeGanYEtK9ADt4fcfn2nl+Ae6yPPqDtKoxniTfuqMZYu1Uj41v
zKWciHwyDCtVrFeDrRY4HiByPd4lM4m9cwFmCv6tCp4TYXxleToZ3crlU3u/Mt4jFbUDvjN1Of9L
JejnxTjYqfKPCZv27j2kVnNGUSxun4djDO13AwhTsPvqgMvjLGi//eKVNvUboOS4Lk6y09e7au/3
+tlMSFzHoptmfy7DsknylrRZIa6283+vVx5xpG1/x/fbmwkRKqRcjsEjnSEeQ6LR/F2lWe05GLoF
PVoVBoUSMzJWiaNbrM8Eg19xvGP9y3IRqjQwT2Nn9VqhRIu4b+Q4QpL/gzo8I1VxcZetIMGG7VIM
jhCaoYIuRlfyYzOZC7IKttjpqDeM1a0l66THcJAb0F8D4T8cXOMNAnhD/cxjadDZSzSTw15VePJu
EM9533qA+ZJ2q4SZQg3LtlEHS26dprAxzalmUv7r38qI2ow3f3q5FcF1gRn9e1qMgZACKLoD6899
EzzqUv56SNb2JWoo+w8XpggrQdfOFiqVNpcGudlbKsK7zEqNlzDPZFlKFl72aVXjb14zgJGwVZSs
JcDhbYTeGlUFYgk2qv38QIW7I5J3ziRIHEcCEbuKnrXUxyggYtmsS6/KV2edtubtxAf68keCvgmg
iqwXod9JB2RtC9l5C9+6ylerF6kBoSD8b0JnYh2hYA/iGLiChAWsxDN/WSqT64HC4EtJyJQh6AcP
FXABbIcBzj+lbNLsWz4X2R0Ch0HJ/Eno5T9YA31cgqewguOsJK2U04QwRmfXBh0ayyLzVkzEswai
vbI5V/GsucC5WBs6R6FOvmL/+6In9Qfg2fxa/8hhe+9c0i4M/nJQDdGwCAIysvYKETWtmWM4OO0R
81svvtEwM4G7UuDu+AdihC4/PhlxRo9a+fqT2VbZFoKuAnDYN/reGNy6VMf+dKlBZ9DCL1j8zuC2
uiTd5tyqIQnhKTSwreoG0IjM38VZd6Iht1+RlgRVw9QyBSxutYX1MZ/RA0mN4DwT3JMgT3G2QNt9
OOhwiWPU0cRw9VoS/jJiL+07saSFPSGnU4esG0cA0EX4Fc0GEumIs4UL0DQ6bj0WNwxxVn7r2nSR
jeVUcIcQRZE8nxlEP6K00HSom5aIIVSBycYuHV+cUWCu3wuUY1Xe7XEYgNkIdsfQkPPgVSFwG5tc
01fXQ3zV2GGYyCsKEQE3lxEPEKqUY2A0u/EZ5lhW8/YTiurHTN5OsKaqaOtNHhQvTv90AsmEYcg2
Q9qNwTkS5aiElV56TCgbaigRzEkTMC8q7KK1MBMCEyss/hiA5p8M/gsZdeMGoMWDodqXInzWl0Kf
oQBbyeAUSVLUZnLXAtz8WtZcGFj5joDTVtle6ePl6Ml+9rf7wP+wbh3+s/Sa54XQZv/4JvEOJZL/
JttGujYowilmeFipJ2IaKGm0g3Xm8/GNKhVhpKQ0cDzCXMokWrk/R5vGAd+HOftt/Zzy3UjP30/y
XFrbjkHjQ4q5kw8ameZBfP2/ZeZCU2ZXQ1GA9ZZ+S8gbdUK6D8T2yVeNjtW8Dg43M8QaV6dp9fm6
jtTRyNIMc87LWX1b76SuEnR429Un5XN6go2FQZjHPLcxpieJJTztOQ5sfbuJUoQCBRB19PwyHfIN
v7PvGN5UwcRUdYbxMMgUQ15ReGbrarGAGlJY07zln2As/Y2m4N4JTOJpMIj9Zqg/JvntsaqjzAdO
KDaknE+H5mIioN4C6/lPDtgSnP3mcMrKKfPNZD1CBrgPyKz81tUZEALP91YSTgGqTDt8Gs88mOaq
/Ow0fCzYZSioDdvfHJeTdTcSmPW4KIPmSd3A0NgtFBTrBAksvjGwGR6/5B7rFv3jsDyq1WmuVVhQ
mb1agMU5tnqCN5nb/x39+mzz6dcxVxcsEJqsSa62xiED/qrf1o9eUCC4F/h/8WRe2NuDBxEP7Eig
nyBbKrMS1mu1uqvIpXaWUkrcCwRaYs2rXJSynyBQf5RlJ/C9gtF5A2kqo23Vo3i7XEE/Jrlr/hEp
0/iJf6zAHcMz8HAxfpIrYIuYgn8Ey0uHyaYmWQhU2WSpKQ5h4K2Np4lECxVEdyM5kLSm0fZSD9+X
pCSSEfqXGvRp/HE47ft5rnpHzkeutb+sH/g3Ud//YmlbLfNOgfgowxReiQUcP2TtmxZwGSHSw1ds
IspV29ablb1ig3FynCU1e32oC10u5USeWYrC6YpyKCTea2HfxyshnG6hY+pk6qgbN+b2nqq3BRp1
2YTWDKrlB1tkt5YgqF6KCDLyVK77hNZgy6QlifGteb8cy6mjaxwRh/6xmZ++g20pFPLY1DTevbIT
TTp1nRIICB0KBHaEpCdDRQ7f24fi1Y3Qra7Cm6m9OL0K/AdYCujwhzBeYSNwgSZZrKmMT7Ea2SMm
hlrNaLxxUNemfyAFFu/v2vn9aSqVkeQKMMDd4C+HwiZN+KcGxfg/g/kepXrZwBIkD8UhTEL/XlGz
sjUV2S8WJisoxDihRyCo0vITVzYRKlKe4bkocWOyCnQmfnlrD17ZD46qrQe1FwnAlk6KeDEzxmOx
zalokYlp1SUBIwo7L9cZFw7SzfvWSrddx2wGtRKrTh+f+ehNi6gwtHTmsc9cXwzt04h0L/HtHF67
63DNcSnDsg6CmdkZPVsWR/3nfdnHrucipUD5PpCp5wFgXulX30czZ2PdnHB8H+a0+BO4OqaYIJBP
nQpzlhcFNYdGEbCCFD0BR6ZVyLmaZbEWIAZaihlds3F7iAkqWW7Y8KWHttZEE3ppgoQihyEs6CKr
FJ6CYmN6Hv7S1koN5YCY7b3jpbEVrIyO/NUkhlRbmB7TDmrl3gkvR/xSqAY2HLUdBGbVLIpmizTY
799VLvc8qEu7oBydsGcqnW/mNJqkrpgq0yr3cDCj2noTQKFBZmWZED6ejzsVHMsmtkzRrvnVVjWL
tIOVVei/LxQr7TTEW5oD/J+3gqsucPz+QISIO6DWwp+mylmrKSRGmHOGxH7JnY5WLxFTbYlbpbVD
yyw8vVVS1BrP6Z4WjWAcKZ05dBV2mp0mAa5J94RPh36WSe5Vfp2w5vte2SKsKBO+aqghtmTmtIyE
diMmFDW4sr/AAZmjDW3toXKjouAWWmoV5fHBTFIgA5MEwN68+9JAJu33LUq3+4JU/73Ynnq3sXgm
oiZ5Tl+ouGRLn0nJuliDSdfMJJm7iW/lktTU+3vocXnD8hV5AGmRxw86QqV3m29HfR74LtGJISoU
VSbJW3LISdFmFwz5iWTokZJMK66GBvJ2v824oq7Ze1ymHOSB4NefhDpKaK2z6Lr4RLmsjfVs84S6
43Ca/Hl9O9NNmv7PD9yvhL9UYMP1hq6zF1kmicnlkDPiyXfNbUdxZc+cy/ssTSDuC83t5KZHF1fL
qf2I3fX0rFSdN1UzOpey4Nr1rboIRVTEmZpnUeD72joNNHxjpjMtG00Cbi5im8Wi/ftP+e7raxVo
ERhK5yFCfDY0cLn7YfZu1Fom01mf+9v0AXs78V6Yq1DfIs1uUfrcCbyF6KlXWfpgGZJyTK4dw3lg
ZIdVYeLQBhqgaRarhRgE17EkPM74NrUpUIPUCCkgR6jZCdNsrpC81wt+lsYX2QONBAes+ZtUFjnS
AMyXNhaaflaWceuOrfT5V6DR8KXIdrZoSbLaJ9K60a5DTlWtw4B+U2DRpgcIjyolyBkG6qplEmw7
n63u/8KHnCGLywDFdrSBd6Id3Y3QuboRMC0f91+tgJjg0qTCsjoz5AQxIc/q9doKwQC3l2BvWAIe
qyvPlGxlo/kRy32eO3Fjv60ol3v3opnusrD2w/nuImXnve6hvBqGmT2DUw8r/sJ3/xDOTlZBZP/2
KIF9/PqgjFJ/hFyWgBEtozCvo3huIqodoy//j0CAix3YYldte0P167S4Sm68yyXXbOkDtR4L1yOq
pJC72zkaFRK8HM6ixQVNmKFU28iTHkyrQXTcDkigBCmS4h1ZX7lOx2jKQCAsti5bkLzH3UuNLOq+
NKLCc4dns58PyeTiKBGe+i2U9jb8uQEaFe/R7ALQf4y1Az91M/4dkU7vvw0+XNcR7ox4pUTO3dgK
3gr8ekz1uQzs+CVaAicVTrVzy266ofR/RuQWum/WpyVkJG+rBusLe7IK23+ECSnJEx4v/CtjpURZ
Bv1twnih/d4DBxTXFgx9iSnswQP5ouEEVROeV9YmBWNsSBOvtHBZ9kjlcIBaszlg3NYuLYTggGkl
WczSeF9gSM3t5M+3dYi2Oz6H/KMIYFzAYYuaBTwxKbrNTIEJt6E5IgUJEVNxZE2N5NDwkaFyxD1T
Zh0y3W62vtcCxwNKWGCZJIbpTNFcaymN8AFWN6hiuUNCF9AwWhqcs5KwVzoeqo2iviwm23QFgNyo
TmFmhcmp2GTdZCSwFGrCyIzhnQayCT5ACAYOJ+HY2MRJl1Tv3dRnCE/t848/Pep19Dz45yjRa4Pr
ZupcbcUayI0DXarRHezaq323y3BqqgoFCoQRk9DCNkVLD95Pln3sEb9yDV1t85qJQUifx14E0kOQ
vDD1ldAfbsmf3QKk+dG2fT+PVNSO5yqnP1F4q8lx4JC+mI7LarDiy2terVbpiDkkGezjxGOeLH4b
HeyXdOx7ULldo45B4A94p78oD2EFOc2Ijq8yt7E5hpi3zmr1mJlp7c15TOQLegmE8CqDPoLhUJXk
ui2iEqd8cDzxG0TWNxoVRp/iZ7Z3Zu+0T4acQMof4AL7FJIyErujmzZhqCHjAiOIF+ePkfcHq4q7
Aa3VW0PQ9EImAAe2ms72rybKM3I/aUpOSQcj4QdJXpxgBdwIh5rJemjxNyNvVbqRNTu5ujlG+T7e
hpPwXNQQVN77zXgIS6XfafhaPvx1V8XooqfCW5Bf8INQbOgxe1G9JTja93hOzsz+JlbphKX4/R2Q
hJ/WksbrWIMeHtCFGu5NvNcnqBJzLt5n+By03I509aZHmn9HwssuSFcYBHMXc7OaNuXtlvjXFnCz
Z1geEcTgLcbwGxHdK9Xvs9gGCj4NluDnohATcQJKXGr8QKp3FIpueBxpP2eMFVCqaI1ons9X016N
BPVx3rdgHhJPBGR4e/Qs4LaPH9Q8FPWwDONXbJ2RVIzssGDnMW2tl0cTZqp8BRRUcIGqwqvVWVZi
t94chRRCXrfwDVd4+On4qzOZysfkgFFQ3DrAnWSwF5fa5HdBSRxV3LZVDhSTeRZ/aXh+ObKXXLEZ
niylHPTyxKngAYvcKTqiTu4VKyS2Ttyi0VpXhaUbpQq50jj7Oee3C6YTsEk00xswqMvdQgEMCxUR
vh3+QGCHFrKwBUplk9xQVUPxc+ObigtfJ2GhOQQ1NToEP/xJ4dMYV1NkWUPau7/wNkgWTQqAJnbr
WVcMRMqziBI5ktzBxAEuyexjjXPlK8YBa0UwjEwbm9VbDVcB7ONzno7m41AYRM8yqXVSgeDkZzQK
UvMEbDbDMlysJwZCXZ5ZuoGnvB2EXTwe2M2Pp9nMB63SOaiD1S5SapyvLxn1F0SwiuOCZLiYp6bU
m2t2qU/dR/FLyVeROl9kSsQ8f0coAAa/QTxSMjtqnCDWoylbSX6LjShDW+wWITFvkLy4CgwQT08z
7+c3F8ti590/tBkWqyWjE5Sdboqw5VFqegLCD8E2KcSy6iMKMdVMrk9Au7oZLvc/6cgudgTpJXyc
KGEL/fpExX9G+c6uwP37fh2Z6LEunyOHz8h9KKbw0PjIE60v33K+ZYINRx/YEKJLmwAf7R0GM1RS
wXkpwHN+n0El7FW236qUY9kyBkzpj5zk6yjzxarMZ/uy6aUH7lqi8Pmnm1P7RK1iDKhr5JH1hAI6
qN70XrkHWm+6TL/gG0BUYKndw+PfHEHxBu1/Y+rq9x1Rr2/jHyiT7Mt2ZVH0riallRPsqWBNOZrU
bQljyAEKQ1Mo5DyXPGFgU5oZzpBzEAdzpNlrAk3ALV8hcAHa4o65g2f2LXn381fVrlz6P9Oi5nva
LkeFDLvmPhAlSKcVArrIahoLJWiqEBdw8eDwm5vuBW4rkftfisqeJi30yZ8CjgX5gqU67Dl5HdxV
SrxoQdcHUowcEbeRZlNSw9NS57pEYHmhS/RK0lSXxi7KW7xzyMR7PT43yUhE80HPHelkhcJlTo9V
tDjbX9gVPc8NZq1MzQt9e8KB9Xxq/scB0VMvtrmwfGOA4vhJlwYWTE8jauYdzZ5SmsVR9wDm3tba
Jo6Kbg5vKOUrb6D4QHgY5kwJgb7RgjU3HjTTyAD7VsyAJ7dSY1Oc0fZWh7G750FOc+5UyAVFG6K3
oC61/87Hl4gcWAtge2xMY10SAk/SBai5SEkZYkiCaT29IuWINwnzg6rhltvrlfc2WjClE5fd1pHL
rTRO//3RPCSaUKjvVlF300MCFRQJ92omB2YdADXLae9zFWE6nAVtLj/oQBtO99D24uHcRI9axrR2
xsSrbYs6bD2jibzKhnQIiCdaxImeZ6xCqhkRURNgZbzpQ63yZd80JyqFiob6KroT7kVtjj7g6pe7
HXG5JnvwUIYaRNG3gJeTMUj0vvK7woPOqdqDOXok0aF6tUDfp1/KCaxDSWACK8qUBNW8Wwynk8N9
//eU/MDGs/l0ryksF1bOgzXDYYtDNfmWvI1QrNibhCnE/5tfJ/HXIwc+YcZ87w/GM7ghEvYw1GaT
yh9c5d0zV6E4xvl6gAHMtbJPcBtHGfvT5c81alY7TNMTgFF7uZ96hb2/1IlgHHl3NEfAcD8i1xpR
SQ146cqRXpfH6bMXN4y0GlcBnopgEnkmnqJMC9DpL8pzoQXOWdqhwKfuJJDOC2FBbYBJjzo78NhE
WPh00Y+8bdV1ym0vx8IR4EMOsL8dlw2Mg1mB7nOb7Bjv5x2moOed0DsDFeOMmE/vxZeMDxjqv3jJ
d2enHPoUsE/nGfpvdQreNZT8G/0B0EKbNv1DhJuRdgHUnML6LCaDrutBo9UeDj+ce/taakzBA4Ic
VR2ZKipxdTsloTjuzffzIN0A0CpqYBvzbtFGCfgCJ6S6+FphBkyyCCcwmd5oMB3p30ZDatl/Je8H
wLh8fI+X0GX8gAgklvk9x2Bi0xsy5V5kFqO/kc7F8PFDQ1VVFWxLtO64/XmLnFCmQiQ8e1SufPNh
j1GON48rroJqE1R8OYoiYa43ZArxpgo8dmkToQwazhmSrmacvl2aX6Eaw2P9zoHmmq7LfxmEPBRA
CGEm6fqWbr6b3Cwk9ObqKNLJKQERfNqLf6/2gAOn40cB1zB7XIPDxlu6OoB4Z1aFOg79t94TeBsZ
vBRP1FL5bEqUzP/FSjhznfVtgkRyLkkuXyJ14h0bW6CzjpoFRNiP97vm2w5JPCGLiuGaX70bwGad
G9qkwE3d+t+hQoGLTeO5BkcN3zfNZa96ElYv9C6gAxCcaMT6gkHFRh2/mZT/6LqpDC4M2FJk3vl5
mnJGI9bkxQnA2qRAnkWXM9+zSajNh5sx1YcYFFY1FNJZqO/EAImA0oakvecpIAHu/G0aG8SOjFV0
fH4M0up0b4gCVsbUfA8Ksp9LK30RfgTnw8kq6LlwIHddP/yq5dYslZobiVhTB89sqokDxCkNSbAP
OrFQD1cTZFhqSlmLK8G9RUGTVujOYY3HcA3Nnh4FL0PvfkUvtCrcGVwQZf+bKLTgXSQ5Jt7YhOM9
iOYT/S6CNg9Pav9fRylALeZcQioR4wTRrNi2lxWO56LPtsSkuy+qi5vC8lhvI07nB+JGVpVMK4Cx
L7GfY93oY6ep2KOFIDMw6TbfOz3xalI69U/OT88WudKOMLq1HQw0/F6d1Op2wtWnZ3pZC/xIy/Qp
IWiBoM+OTHYy77gDRzno+Ihvynllx1SmQZ3JDqCgHBcCuYQIf+ax4sQ8yqRycVtivbJ5RC6xUMn6
hhMULlKYqSj1pH/Om0r5+ZiTqtskksB76M8+MHg2PnouMs7wqE2cpRaMqctkCOkN1lYAGAzx6eCN
WgZ+3pm3uHfSO0RkLtMtV5p27IJlnKjw/ywrdI/Atn/2n3FXfOyk7p+9fPV8kTamym4TpIqqJcNV
Cok0GFJ0gIxbWcU9CufwoDE+uU2P0yjAjPaZjRiFPwOPit2hBSThmYZ6ur74Mb2tB5m12riiV6vd
VNv/MSGBElPUGnbujK0AimXIXq6tozHrmlgExUJoYd+OATTDBFO5mBrU16YOlGDgFZumP3gv0QSE
dLpO0ZhvA0dbHcyn4JqdqVlXhwah7ymemg2W1MOteG4zNJw15QfeVAyUIbx2DxEjhMW+dXDINf6Q
YDnGh8pFnOMVgZkS+rjV2wbgQ2Y1snaWe0RNQEnxWBBCFzG4CNpybbhBomdhOZR3TxtZJ3A2VwHE
qmog4zRn5hrJ3SfdrLtteSa4JpAQLDkFmeHHPzp5DH8/aYxSBtAn+437KMtV+ccsHs9YpqdGTN3e
XeljmLfZNVk0BqmfBw9EVK4n8MmUNf8QztTHj8h9zXTF2uErn8oWGMYQct6mLyLJoiHQ+Jok0rmB
ufweFqW+fFRE28mF7NaqtLZYf460056ShEoWm8ZSBpESYSTfYa5ZE7OA2Sq+fyeF+5JiyPyHpcSw
o+qyBWpSZRRLCkyZbN4nNeLBojxzUyo/7FbBoYLbnAHrzMpvzzJ6VhTswedb5XSC1SYlwk7PODn8
0urnf63OwplN6nrxAbBF47926Ui7JK7ulX/8YIt8ltJQ6BSCXOe4WOtn2SHtv29wtKSPVEJzTkCg
HeW14K3yjmBIpk/GHeX5xv4+nMAtgPq8w8D47QIm/53m2nsG9cBt0562LzTgICIflHHhdkomdV3f
qXKr3SVJFSEg34fn2zODkLlosjPvltbzTFab33ztzhula7S6AQaUxZ36qrAL8laEzbdyfzDGom+j
ofOWWVyOBCczQ56PhNe+zsg3OoQkV1Txl7su/gRNOwcSF6Z8Ki5J7NAv/1B3idOQm4SAuPlKWyAi
SvuyTaWpL/Ao0WalE2H/UYPTVkBGkhgaI+3ZmmLrjxUAWFcO/Ggo5w6Yz9nu/l5uDRhjoAWwAUup
cYey25DjZdv0KKLCaY2snUBNqAxugPvjiGER+aZSRK9k2O0L2sMFY/H17ssBsEpn6OcB2lVG61df
NbUG4Tr3kVYuKc1VvQb9NlVqI/C+VoSqG8qg61PQBTEt++gCd/T7sMcPlREMlKekRKeRnx7y/74s
3Fes1Z4q1fvU6iXi5KSJqQ03JOtkE5SVu7R8Cqmrk7N6np93Oq/NhfoZBdgk9DeVR1AHMEpVG0OL
mA/UOeWJ0ySwmKxb/XNAmopLZZ5LFPetBef+UI44hGQ/F5sfLPNYtdtLVf/icjypvvXMZvC+o9io
+vkeueUy6fZjzeEO6y4y5gfwB+Zk1LmEg1xPdcexPdpdSE6NmrOl7CdbFqXNcQaFrG27y+Upwhpd
Sl9dDlETDyZ/JO6KMuYtFZcqA6F7rY3UxAG4RYGa4WP5q7UL/exBDEf8kq6k5EzGLi4jsllgYvRt
EMmUAoAptu1ApHt7R1rsIWVOn2DoQ6vxnc/CPZYX/P+t/WIOARIjLa3Q53u0panrXTiOTdBLxnb2
Bx6QcokOpqf5YdS5e2sXU2h60FVfengJV3YjFcHKVLm1d4hPQ0FYKnAO0QZuBiR8GUBuUqyxQ/V9
jROEjS9zTU/MufOL7+vkUBobEtAvi0vCI+1O8WfaXvgqLM6vtMAV+qw3tRnfJ8FPvt1Nn6ZjpDE2
j2xpE4lNd4nGGaMf93TItR2Lr9tIMmQ2VBJMuTmSLnT0gsd74ETsDou/ldsTtNSbP/FfI88Ge0tN
RfqzVJ1xCGEM0USlUAAtcu5ozLy02y4IdJ7uc+WZOaw3v/L+urhkNKoWb7w8/OKKdtABuQnHWaO+
PsZykR5liCmPyngxQwN0KXRaAAc4skA2DxvTC2O9Psa0bAQgV+C0tv1DYXVel3Yw4Eqtc2hxKKvj
amETp7IrOKOZHksF6psi6lboKmLGrs3b4RPp+SWbL26aN/JiRBMziM1rkWWeuLeqQGLWVReJrN8m
85jde1+ViiCHqg6vOYAyfB7j9sscb+LWgUQxVw0zuJhC+vtNSCpyYedjPAXf5vP2xL0QND8jjoFI
eRbe6fUaB7ObIYNThX0mRc8bYoHDZm9BtssZwl1RzF8onu0TknAerv/5xN5Vv4ZNhF2mhyOyppgD
eQ+m2Tz19meZ127lnDPckUAfdOgZ2RKvueTMJNK/epooVmcbZ5zCE4I2Fx07MjQcsSbTM0qN6llJ
gAuI+D4YMNB3oRpGExt28/s4PGZ1/8S2EBpSpy075wHj//jLzG4UUWGismKS/vTRqWbadjG7iKJe
/Ll86cP6BhFzg4q/pPOI+/RCXfbfeOddk7ocWexn1zIHcPqiJz3uw6YjBmqhjzzw0KtQAVa7Cwvf
W7hfI1ZF2v+B68EJFGx7jQqFwNpAdv1aBTAysYL8rbr6Ye6VTE7BoeZstzCSACrPxwOU04vE0iUI
c3nVe8YJM+nACJG5zOzyl6Kn3lX9jWEgGsIIA63aoZg9k2pGRP4ncJnc3J3D1BEE2rnCsaaAHhWD
K1WgPsQM73DGLsvNilSMiQmh6ygYZUGQ2CD5TLmjhjOcsNi/QKgJr/q+eUnyk5FUwmrWH0mwW6to
wioObHQdtH2/ADxU6aJfZn0JhgKu5MsdLhShnn+2ivEylH1ayqmHgKxX1Rsfp9wF8OW/vJWX82hn
lNeYfEiB8fbunQHH2tXipgb/vDIeQdDKBwROPsznlf7wE7SDPCaVCryYr5+kpT0dcUDuCe05hBHy
wvwYDZo0FAn3q/HfuZbIDm0fdA59S3ZbVmGa7O1cP7u2dP052Za2dtcr4euBqEC8adbzP282Gw5k
Ao1ufoms5Y4SyTeBdcT3qYSz52ZueXVJUdeP+uw4gteaNmCDRmy0yUJglpqjDXPHftP2TZoCUVQA
G/XSSXnc47sDUyZnkE93M/+QSZ7SffhOFTN3M2abi0Gm+mdqS5x28dCjAdYXTUqZYXp5w4MMO9gS
5koI3C12D1ez3YpRGGCDHA6dyBpgT6ZRRtGNBwmIx2UzJv93WBgKXv1rnojp2BjK/tWXwiv5XhF/
Kqxrt/d2LpPfQRKnf23jZg/usPqRoNyb9VvVhZBxXPSqEVXvGHKEMFGjR3csitxJgSI5wwXLbXy2
QJkmVdni8j33Yql1Kg9nPyX9Lpauj12ssN/M/R1HY797ySd0LZzoAMm5wfWQQN5wUBzXuX8Iiy+V
GioDxhObQPQRH8o23Y4xJY67J3UyOTltrc9fe/Ng/wi9ZBzwfZdOT65hqHXWfg2mp2U1U86qWwN2
jwmJJFoT1JPTiYywWd/uBVOtrfOK/HFEhktai+J+qUrkdvhDEjWasShzyIOxl6JGeZDrkbBo3sQ7
eM6ueySNR5VoVGvIlX9+MyRseEaUroNNPcv/p+xa18Ol1WiRxmlEHLZdzJ9CTSC/d65pkcS8lLnI
LuTy4UXm10naBStN77jzFoVSiV3qvgz95VFpPsSmxh1KLf7z4art963z/EW++mrX2MY2Zj9jeyFN
buD/VdAtglCoNcy7sIHkFnPBvpA73rCDTH6c7wOKV0R4G+FVIhacNAU8sazrhWtRjn0bLn98aX53
GMJ/p5+mXEnytiWXWdIZ1QoColvj2Brergc4AO3LWARQgNci56MYqSJtvOPU6olbsNGSKb9Rbk8o
TqxoKExBIJ0TZ0Oafaj10pL86BQR3nrnNemY9VeovOlRhMOOPoJ9EALAgKh4lNEGeB08jbk/rl2X
sU5duf+rWxUB7vfu+rJHfi6TFBS5hBnVAchtPdx4+UD31UMyUr9EFit1dbtO4nIx1j6KdkueNTPb
ie130Hn67MNwRzr6myBFxcA+k3T58qBTeoSdH4m/NPg6PnytiBNXLO65WVeM/Utfo55IRGGekWnG
u7BXg/4cIBaoQO5BxpO3uXvpY6A2UyEsBJ5Wx+ompUK6dKTazt1uXxl4ulq9AOdLweAXvSvK1BsT
Z4SvcTCI3rzM6cYSP68DJR0og/nL6C+dz54LPBby1u2iQSQ1ZqDRpO57mqEErYpcvcOATxk1+v52
nBYpSiGBJN2WS0FsLFI9WUtYJ3veupsnHOfWZeRu1XtMMiKpcEVbj8/ofzmcWIDbbvhQs2M5954j
OaIrHaEhWmknsa2oKAvvHTumq+GqwsvOje5n7Z95H+NViQXf2XwRir/28Za6mEm7Yu8cmpkUFZQq
f+OipUhaiKAl+sydGUxdx6MTJRSoErsQGs3Xbg8aKP+0o/Z75+q4uPd+hwBHLSShaFHkIxG5p8HW
mSCwAWiEA3M2BdMkYdBO889wjnJKlO3i5LfdjGQH2kmc7gwanJ8InNK1ygDoJGTHApJJWgksmyYb
u8SZAMpxQwEZ8/GIXEV9Bp+ggwnHefdLepCPR6YOd1BUqSo7S3ylwBEVV3sHB2lCWHHf+RpmBLfs
nr+dwtlyqJuqyzuTu45N/WvzHIw1zDWzvxCmmqBWdr9gGyvzAq3xeP7aIpw0TOJBHCGunm/p6EKT
zP4iniqtwErSLfQhdgeBibVoV6tYNfoqT75KXiIjjmj8MgelGxCOF3frCYZMl0edMctR3DuDNPUv
Ierd1y3ztDMfnleVB3Ps1xXskl8OdAlnrV2HKUdCeOITsGVVq7AD9R+jKK/9659F0V6zW5dpY2C8
xv/V7GKPdxzWwdswdC5zi07uXWo3uNDOQcOVZWP9Az02UWoHFbdeayXl2Q8aYy01PY3d/QYvmAhy
Aq9dZnSZQ5D5i78Fj/nnGPdFK4VnfjjnV7MFMLhDJsBdaWOXZq6K2lfzYX5XCnDZJJafYU00Q+Xc
pJ48PTU65kn3AMh9L9afpaKpZ6pQvKv/kRzPYKP2y3fF3MhIbtgueNGL90U6L3kuZTQWF6PutCtI
CNolH76Kg16k36FjL7eGSlo2Xx2cyZPCM6vJiUC0hrmS6E7aHQWp6LlPeYXbThFuELswFmarGhJZ
WyGOtot7zGcHIniWSUaX9M0IAJIa6J0S3MlH9Q3fYNwsDiya4Qjf3fdzz61PXOIAX9oWb8ZyV0PB
i9f7gEkWIKvBNLsnW6Vqjoyql72zbRujUS7LTue6RjLB/fiB1qzqpq7QEmm3cKSqtPf/YdT7Rt3L
tNgtjt/MfwEFraz9BctkQrBqcJKj/N/RnU0M1cds2QbUkNK1SfUeMV21ewEXAnHYwYisKmmthtvb
lxeLi9FwwH/lBYqBEofrZtXdQC7HMC1WPbUNCfZ8Xg9lhzmG0lGQt1V+XZMUBcQNVc1X7hENZlDK
2K7DYZxUDSvHkSVlO2MGo5+q3r879tORYaEfseU5au0Op7FyWVp6A0SDcIYeDSZnMBSr6s+RwuDQ
sDt3OCSyVrOL3FHIMGwDReBriUrvD/kTYnH0vLW39psCC4TzORyCRvrnvngPuhS9Se3ydkNfd7i8
AVrZH/khD50ulkQJoAYVDiVtYrXWF4qx21ornxDM/ZGKvD8uZoI3lfVPDJOZS7ueWm4sBsOCvgb4
DkFp68zZ9nZfpvYDs/f3svVRgHP7EuIypvPezdmm1oqEvdVjtCaOz/HD0XVttTburIJ2vr4SdJz2
u0em7HviplFh6o7Isn2LtlDaI7sGvpv3oq9RHDejaLyMSrs6Ov8YCmSLW5rdw0t/906t8UXZ3ZfL
/ZeIASSn1sBR0w+kyjQmEZHiqf0gnn87ZOFymu2ZzA82p2zTpyN/+JPR6wUWqi6hzZq0gTfHc4O2
s1KnICqj5I6R887HUFPS5djmmKkxsolA2Thoi+ANBzYOTDvyxeAitsSv6HNILPaJoWFwRLINxxf7
/yang10lWiHb5F96+QvgLgXpokXFq0cAHY2HdMERwCwzSfIpgdyf72GSJXVmtc6CcrvXRKTNjRWU
tLTuikLaOfy9SIBpBIME6wCXva62m7QgJ3RBOgDwcI7bINDGPBX/I/GKSchd4M+r7/h2ZocEDeSi
6u8FpNblbPio5at+xp8ZUo3Lhz1EJwvJMKfwJDH6KdDzsz9VICso8Su6OE+xpukBKtzf4CpIluAf
NtI+20JN61xWa1rwCfmi7douC9XUdOSzUKyfAubRIgRHVPJMdUXZ8bBh2e41xhO8UZ/kSd3wM4ar
JaCWbWV6eAddYI8dhDaW8880fkdxIlj8Lj9XxnpqvRH+hswwvVMV3UWApo4KCeFNXH+Zwgn7tZg4
THaQYijoFSJ9rvJ7NW3utMm2GGILAT04nfD1oWJhAGUEgYJszKZvJYOmbssZ7/YVRosqYS3NhO3a
ZY5FyoVFqSeIMiZVS/gQs5BiO0kaIBqs+oAe+dhkLnRKHic9WrkQU3Ebcgp4q8br5Z2L6Xr2hcSn
cv3feECUobPEZomE9AGaO+MUaVjxJEYRQmJezWEmN6AdBfZ/8PPyv9hdmHbk1+N2Es0VPVuTXhCI
dCqOLZ/Nq0/Jvw/gDy2MOLPNNqS0pFwR7khax21Ny/SEa1YRk/IKWfyYGAErWhA3eDIfdfGqW/Oy
FgTgjsZIewXFV9ELxELxEMFvzw/nM0zbcntPiyRMqjgHJ4stoKYRArSB3OsfeHogsAE98u7njJsM
6viZQB2hXjTMdERE5RuDz2wPwNXg/AjNT3F3gvm3UNIPEv1a/ygYsZIz2fGDWbxuRm9D4aVTw3R4
OqE2oM2zVknuLMnPqyk9W2SbqQ4bi0LDkoL6Jf2xTyj82xyhSH4EsHvTsuthYS9cibaK2U3ZyCjw
VPpHb5eIjtEyJ0DGaKx6JMR/8xBRxXcr1AQSaTsTbN54RJereOMZEp9JcIVcvDeCrwIQI1hseHi3
A0o03wrrQ248VmJrRRKS8cD+oWnCafDHsRE52++5+CtT5TlEeTMQIIvjqDCjGuw3gb0m6TICCDUT
8/qCcx6bB7E5kekIAa6vy2qYxfHdabJUzDeuFJ2E7Ca06PkoGOpdYyPLC6Ymfgyj/K5vYeSov7xM
IubllcWOX38PPedVtJ95CxWRtk7WCq7HAUFHdXwhFHqNpA7/no/dxKN2nj1y4UH74yGPZiwv3MwT
2hUMk0bzZUjqJpX1XAjgLFfcD1tWsnAhfr9J5oZDWF9I7nTFC+TY7ia748vgCVyvuDWRCzNS5CFB
vNwbpoUYS7pKflo5hbcqiyMhcPIoUmyuB0Nfd4q6JmE2LC4R8TAymF9yqV9n8O1KJC9vtCMQxfB0
Y/7stBP//3LtepypV+GsjDYJly+nTx9GXVdCBPg/6E3z8DcJO5sPoHWXRKp5AZK2Mjzty+yrj86a
b7TGbxiL/7QBmqd6/8NWwyujmV9AnG6zH65XwckAoFvlxdg064yRUDvPKo4oT4QZL3vESJ2NL2rK
q1rQ6/HAQ4/S59gjNNWRYXOFAC9d4QImPL/bVScEpOQ3zrBwfMpyhKEWToMsgPDNVgzG+Cu20XGb
6dcT8r+DfSZJ8LszEl0Ilpt9VS8BXx/G4M+JPztuI3JNJkBN1sMtMpULWScz8T41/w1Xy4ndhicr
h91BZX9XiuSFyD4Tnve3MSSs8dztivCxX26ViBZ4/8MG5mCzYpoogWN9XNIgTd9V56j7qz77PJax
6xydc717UT3mfaZjUf2oeo9NgdetK6Et127CE2Aze6zivoE+dUUXz7S1/VI4embrV4qbnnL5aa0n
TBRRIGDxmYvRvLBh/S22Gz7QHI/XPT8WGl3yC+TkXErO/EdiseD6eD1qv00qCNC8cm7NL+zVS+Om
c8qB8O017Cf7aeT53kSOkn7IiUZui7uzmG8eUUdkbGuEfokD2USSfIKIkqZAXgeWL/VGAW3rsHpr
+ztMo1btCUc5EREylAcjY9BclDO3jVZMB2CeWRLK3WLKNJjdyTNK2i0VJZYa7odzSYe1YB2ISHHv
frH94765afX6TNThAGskNw8u/wberVf46Vuh97koJPBJ4T5J5oc4C20qHJSjBX2eWlAr0xDjXK5M
0olryt6C6jtbqkmBOcBrdKTZfnVUk/BADJ6mljKzvScFeuMaHhOqU/f5uUUo0JabpyGDYb6F+QMc
W32GWpi03jFf94ybkolDdD9YyaRRI8Q1rTZpj/uKdt+5gJzN6ha2r+5tVav0DRVRyUdR7Rqu22sn
9hDkXnMFrSAAI6wB6Ym79uPkjdoddbsZUgx6Nf39ZsEMxFAY6deFAiPMCftNdofXL1QqO9dcnVmc
21QK6j+35vx07jao9jnkoL+6HPpmjCZG6rX57RbBblKRYB6AvULESUvLPWAgcgYlusysYRMUAbxT
AEP2xyTGG8X2BewvA5+MCPXe/HEdMQHfybq5pHwyZEWp2pw8Ok4jJWxg+UGZT/wT3p3e3KwmSinQ
5Zk/YUcPKlOAHfeFplwq8gZ3nvw6rJJoRgAhhvwo+4KMgd9zs422RS3w4KJUYOZtKg0Arm7urXov
qQbM8fSOjAb+95zvuLyVKWiIKO0LLfTOIqdxzx1BFIxBjWjjtmS6s9uRD/XLXllxXhs8JWa/OiDV
vivZyjGiA+DP84x7jCDM1wrnt4nNnjbYhP44gXiaOLMSPM4nZ6g8yXbZE2UEaQZH3q5uprjfJot2
CPDvQBzX9orCEJP0EfZMSllhRb+1cYV9rkQ/RwoKK0opDRkTV8T+/W7u5UZlyIUHoMsOS6AM1K1G
4fjJovpiwA7i5eGBXvGnW9VE/mzKFCReh2NPXNKpNssUgSFoGUUNfwbTEh/S0ehQCG8I/Wdzg5bg
phJvW3yW3R021oPRG6hQ/AWRn93k3IGhj85y5PbIQG4mWbxsFnCk/w6NNzAjllDVQ7sBUQ3kD4U+
Mgrvi5dqvI1G4+bTWcS7006bUNxvhzZIXZSdFCzO9S7k3FE1OQ2t7XsiONpL+4N1mOrHudo/ol1C
mqFD8ivOMrDGSj+R/Kushv/cuQChwT4OtUAxSFgMjJ1a61jtovQ/xZLO2tgZh3knvC26zM5Zn1VA
U72U96a41q66pgHXTceFri97nV1FU+4ZW7nFZH12/dBOU49YCFaRI/esqpH9zpkYP93+Pd3w8uJm
GpLYbKNyKRU15KiNK1/eNCmm0AgSQF1xJTDHx0f2YhfJIB7eqyg1DosB7YBIVUin0cyUbq6LFA2I
TFDOHuQ0jtkkSqS6jDSbmrJXc+lQ/HZSb9vllTT++lDIjDS7t73/RIJ8vI1W8Bx8LD6pKg15ie6o
ochk935lVLnk4XUjf0d23/IW0t+8/0SmjCAcfOle3AvVT1ywp/P22A8eXudxuR1rMnU1MinHXIoq
rlwtZhpfNDkyvLo/PTdQ9xjD6VkLk8PnjTiMbJdiRz3rGT5SNktivSVXktNPII6NEgK/lSb+OmFG
3YpPj5RcuVT30TjnNcrzoUVnn2wiBPZHAFcdHwvWq8AipPTnoAKpT+QKv9szI9WhCqt0BYcQU79h
hkDHeTIuyusqiDWgVPXnnPPMaisPgNZXdJaBmtlz8/qNfxh3Gqh+3aA90XkpSzrRgU/d8NcwXz2h
4KFJC0RzBFV4z6NnIg0G3yrKLv4zaPmorTAWZlU5b+YLvcXZQMGHVnXjd8q+W/e5FFpDVcKfSXTd
jRlE1VjcYabaaWZKSTy+sngnqZZ7iMYZyUDFbMSVMFIATdbS66oN6fz/H4T3cgN2NPTq5V07+qLs
tKNPmlBtinMtuDM8LDi++NnVUg1A/+6VxrAfEbH8E3MAcWhgYG7cI+qkrYXGYbjgfyx0wP0O9wpq
q5BDYEBvx6hSNKDBS8AqIwPwVosHBKd3JyOfmVhlBBzIi3TZg7aytmIMJGU4jX0ga5FtlFv1qQU2
/6iRCQMMrbF1wJ73GCsL2EwbajHoWuNAvJCl0+xX0A2p4sNwgXWpXWOBWi2DJmh0euhkxx1ZQUOC
TVf4qp8+JbPbe2cjmMRYMv4gqfeVcplcJ3LUDreHEudMtYJKnG4rIq1Arl3nqICJN0227LraHOJG
vb/UiI/v4MOelBH2kyXMH64+cu8pUYR2x3NqVHzEKFDNSGjpH2/kIO/tneyGDvSMojjbvpudtk25
zT6nyYRthfAM8SZo/5FdiiaOSeaf3gRCEgxfHxQ+FJfc9XOkwGFogU71ggzfBHGS5dsRL7YkNch7
ovfogxQPxslrV+cxCggjc3hGLMrr6Vi8DasXVLVNAIHUAdd215nEXL2DM7KJVgMiyDM2NkDRRf44
v464aQQc/+b7o1WV8I3Y9E5xT2rxI8j9Q5CejBvrqPMtEd3MWft1tS14D3z6ytV3vnT3TK4ZtW7b
hsdojQFIBIU4ZJ5vzbxuiayZc8zelzC43XG8gLWSqRrHfDpquu1q6Tt1WNW59KEt/PdAtEWtjO6o
uu6GiyrW2cHvb7BcnF/FIq4InUHcq60Wa6vENiDvrTW61JqEhOlHxqNCze6Q1J+pd/hoIUde/xM4
Eb6sCwdoaqbrFLMWuef0sA/HwNHzv/p8XlBBVdbqhLWI8dKvrhgYcfNuLoDGjWbXT054ZI6Au/uo
j+qzjwQTzUila4Yh29utgDAocwggAALcCHLUYycuB28sdAXiMySDDvr8HbMqA+sjeckDSIwBNTqj
vBxUh+PVxF0eBLS5RVPHeaVpDkMzBqC0a5ZCq6w109wp7WLbkawgE0qoI1xP/H+4d3+9htkkq+Oh
bCrTr5ymp2vQPfvAV/ejqNHLhoNVIdy9pHL195OTgLzgYIOIxfuCkWyf80rct5sMTIxIe6snMCNb
vn2FLigULO/hPSNjmMt2ICGSyswt3xhmzAG20pERF7Mr/cTpWd2kEwX+y6AN+LNfcJRo1a0KrNB/
FDCvt9O2KsZ6WjpNmFgL/7AKU9V2hM1SoUG8o/fH8DEkLSmhp8zkVjqpEZIpz7XRjr7v/CrYGto1
fnfJcrEThck66Bx0SzgphV6+6rluyH0allxpiHT0OO7zq9G/b8PEEU9YarGjuXnF62ro09SStFao
AdNj3A2+gzBxwh61LonbzXTJ/kauQCMS8MnS/2TtH5ftlf0BrXDDAta6ci2JC6N+hKciJBzuc/ga
8Zs4xqWZh3JMU6B03eit45i4SxdUi3h4GC8YMaKzuG6/3FHRmmq1WECW70bC94lqcT9qGjn7TUpX
4huny6kAtb8OWaM9LBv93TjCPCgf04eJes1OH0YXxwFRJyivIMKfE+ro5J+pk1x+IWUJ7WoZwo/z
O0x8pEgK40xkMvXpB8gCmOBXfP7qfeSqTPvb0Kl6t0rXsD9wJd+3syvLKQBs30tJwkhn3Kcwdm6C
p7ol3oVuMtSouvsCZppMqCzm4o/fZz/9/JShim7+XGqh2vDAetx+HI59bGf1hD9+QTVo98GyPhnE
VcRR0gHArDqEymr3J8UVD10zETkp62JHhR/TF/nD21hQTkg3njxMQIUW9vDw/o0mD5luu5uU+a6R
8MG1wFKDPFlsP3IofcHYFwWP6zLfYGvuDpTq2VxpiHmRyF18UUeU94KoYv0pse2Trigwu/aMF2gJ
mCntnzsNK95Cr7Vydc9HcIVudzEqvE2aKtsrmw8HD7S17Jzx4krKZtb2ar8kTew9Z7DdUKrBcUkx
1TQMT86AxoXoZQl7YdHaeJBy0grbld6su/7YSVNGB4uWZzlgCoFrcFP3LRaqVwQDp7wTkuAEEBYm
1C4HSgPxGQu7jQfZYnuh8mTz6leShm6PLKJ0w0XOTUwsIZ+344uLMCqwZkJ2WFuXBectXlqDPteu
bCukhfII9D2AQQaxoOXslWYLXNnmoMhUkcuomDD4BBUtt3VwxjrZhhr5nym4BvfU796AR5OzIuwz
0Hc40ztkGAu245noEOq8Tc0M2ARXu2puy+oqjzRbZp15lG1wOlLFjmNHJBX+nMqpvF5VLsZHfBZd
rW3eZT/rDZfMvonS7C9clM4gxeLje/A0aK2KkxfiPvG5mByYH799FQ4gZrPgfBm9zHdq1Cx2LyIy
WmFqGergZrQ356RpzZyCuU6ikhXdkSn6hD56quROd2+1TOjBCNTfw69cRMhg5V8ZnVpM+Uz0vMwY
rI4Vt5IHdoMyjKjwg+Qvx9iParKvYiYE9OF2HivzN4pXZSKHNY6Z/wtdLUj6Bk5HXeoxfPNgvy0x
g47snZ5t/kDZ5Md2k7v0nHAl2RhNzCdvWcCnGRDTNTsTmbOFIDOh0WK/wBK4arDX1QtX2Q1rgmQA
E++Qvyka/AisSX7mRY7FS8PMtnsbBs3GtS4AXlv3oviSfW4m3KdTBzn0jQPxZVF3JuqDQ7/nuZzA
w1fBVjmO1bCyCmxgCbW+79zQ4J8dM83p/N9yLVYeXW3TvOUAMnySs/X2WP+0QQP5EgQO6/DqMjRl
duM5catfur5gnswDCCm3fZWk1JI3QErB8Q9jfV41Q6qmkHCOw4zupWbZnsdyQvtijvogiTzUvETp
uSb9YjsMyaOR3YUdK8U+6HRn4ry0k7hn0BL/txuJ1bXb/NSI3GR28Jf0xuhpuNLctrkq7ZqrWYRg
Q3YmZzIggMeJueOP2FZmL3dyUbF5xPG66V0ff2VZ0YRm71L/ZeTPZpFKT4/kp6wi2WXzGGFObroK
oogFcfaaM7eOs0E8rYVdBlm8AKdMuq7aAB7p5Jyq8nPUXiGNn4/qF1EBU5SRGQOicKPZj7IS08ly
GZMYOmISv+zZgUyY8v6JDFOhHLDe92b5ci9p01gh39y0Re/I/R6i9LzMKO220XEgeomshcJFk4EH
se+ASd9AZF9rCLU5jOR8W2VZku2nRtt7KIEuCjLib2K5XFASDWMl5D06vyyOH+RCm1Lc8MyBzZDH
mNEL1GioQTFe87271bR/rVd/ikxIE7p/tTP2oIlzTWhRJ2gnO4WolDqJ/qvXZpxGCFbE2xEjbFdW
bKic1wQYBu2k+sb8FR0xv7IylqxcE3YldKflHkOvxll3yZR+36FUK4TdiB8+xzB/siS7xAisiFYA
C88+phPLrcugVFyodMI2VB+7kG3bcwCtaYvBcLtAYvGYVjSCL/+wel8ged9aITVYA3qYaUxjEXDq
Hn9fVnStw02W6kuE5L05kBHXolswdtod74fqgHknErMXgMgMjN/MAF2sjJDDwKx0OjS9R9r2IriT
mny6mgLFDd5QRoUykCGuE7EVOKE8aCjR4D+TwjyiMhrmawRQv9GRNcXOF6dn/Vn7RMJN7b7767aY
Xbm1qd5xvHUyBlkRvX/1+mcw1DlfZGSkW+llpgynZh0HbqQD37mwDklqE+X2kzhigJW3bOBpxKjb
AovtnoIHmGAOrZOwQYNGU3lIHzrR3ab3nt6BmHtRh52V7jbBYETHF4hkZamZKhhY/6xbO1Nv+Be3
FfbZFZAz7NCnXVG+2h8slB3kpydg32HOciR/Sot9Vbbl45Ft7JtZQHpWL1hqprHU9ZO9qoOSW80M
DYPF7FQ4RvoPslbiKGrXcddo3e3OYXpgpeBIOKBDclrHQhmG5/KFWYFT39sb8SSP6Mswwvlq8spR
Pqe5yJx0BbUKeUYRdzEpeIr5eq9qQzJmC27tQFfBcIU5g6XAZaKuhNx0yrHitVsppnLptlFMlMWB
hSseoXARP7q9UJtqdtFH7YYgwLqeQbCPSs7IShqVqBgQQgvnqpnFnXB+NmGnHqQHZJTu9lJYifem
pCdayLSArU1KBB5eoYcYfbe30MwT5kJR8sddUGXI/7+GjZVDG4QssdnQkQVWHVPJkkjVO6hza8al
jz1CxMA2XRjWHPXsMvyJiRNT1AGzXlejMEkDHbaWDNW/hEXhOX8NDhnPd5MaogWeXfCs+2s2ewzR
8yzKlCb3ESfwkpVSEdCUqszK3AggEPDWz8+5o/WepKhcHOp7Yhv7gmS/VEWYjNjCVPb9q0fTzmqJ
1u3mjZdFjxP+upYynOMU4SDXFdB20aJmoubIQfi+T2XS+ayhkZGVZ9e8JaMvgRUIW9VWxdAMZhXg
60N6CFBwKNGF+e6Ja4x+dRg9NhmP5FGyl2RU063nCG9lTIKotNCb+bDu6TewMAfTcFOZA2M1fcn5
q4paA8Qeemg1DnGZr6yI2yqtopTp0DeiWh9++h5+5fdhrzTiphAyX08JxT1NIm0AH9zApKBTK+ox
ZdTmDQfoqHPRR8sclQgEieoWrrGv6g/LjavAUoq0yU1pxE1/0Jf8terWDbaIYnodV2PJdRQzNXxJ
1PAFdyBA5Sisn1z2M5yRy1jNCa7CLCON1RptcAkhmJIH9eUPvieM4BUKos/vZj8qEuq4PgSpGQ8H
+CE1YbKBVTkgumKnhMca+r88DAVx9ZAaGpa3yoM49qkVI9XNsqhAM+fvDnZyLrEUFgTKF2T63L0J
q8wPH6qGcYwQO8bfme0N1U4QGeKRzaE7rZvSKRPtMfyxnbBfb1lBgZEuh9ukQTk4ikQm34ahVjgJ
AV+UgYRbkbnRRg2l2OEpMfvs4pu9Nj4IpabMR22KroE/GSj/6jXEHe8nlF1uHL4cAY+9i7qrq/S8
q8bftD+2ko37mELsqQ0s6eW5ZFL3Sz1BO1dh7z0X51KAnKjUtA8rBtqSu8dtbcbWajZUssox6AjQ
Wlw8zmRYQjzLpUIu4mWaJqBXmdssMzx2z3NOPOFoDxamuXZm7SQnchNZOA1rZymaCPzzRRhaF7Nc
FM0MQEIzu/WgkVQcpHkDvzlAPRREXAU2Nunpw+w3/45FjXltgyc6zC+VF2biBew0pPC/JLOUOlt6
xhQPtMDLWUFdIa+y7XqUww6bSHvQ38uPEt9ghWB4QIxgpWhmjtglOsdXtiSohYoeiJL/HO3JrcAi
NvcocQoT22hKA4kzybfz0Pulbs63lKVQV189EEcP6gSOp2pyxO930fKLry9HzLHpeKg54eLcq3iG
/r7FuxAg/8VerqvFKTGAyn0Gg7+AcUMnav8txUT7VYdXrzVRCud7/G/iwsyRYnqjTKOLnaEO3Ued
OCf9uxVLMzOgpj+MdQrCZjmH6/rIWfIF6r0N3hyxsxv03fv6g1dO5JLkADBjRq2CjYanIwXgvMfM
0SNX+2Hfoob7r3SuOn+BcKzIed6/ZZ034+kDfwNyaMWMF+BknSuObf2+qzYPWvLB7iXwhHlBKPqn
xpI17MuzStY3MkOvG8H4gcrZvTxFoexwbdg4CuiRSwM3zBM1CM+sR68y3Pto0ZpuTUuhD7Xjpd8p
PuPrOl/hQ+Hdr5ZVAqC6Spree2STKS+ZfT9KzZQVIhDuIuIh1vVT2YQCTXgKVEExnvR0Y6AyI4Ue
M/MkWzXVObvjle84SMnqSfADnULEEpoUMXrjC+n3LqMZrYAC/0/wtJAK2yredMbWwkzhlLgwkEnQ
s99/nqk42Xxj4mivg50UgO/02DkWMNGsJkJnnnZoRIFzvNi6uRcEfvta4UDXqC1ctlv/os4+uAIA
dZFzUe4CJCEl7FsikqJwPw9RY9Rq6aYx3tFuj/jmjjn+x0UoEKX/iTIOezEj62eMXA/ZMSmO2SmI
j2PpwMLv2CqOosVR56tF7MvcMTpQ3SyRBgil07P0Yvhm5LPMBFb6q31xp8pvBTV2LNRRLgwqG74s
LS0LItXLZB1qJ4Fp1wIjs30wQXD1HltssaOXA7F1jVmnECscLpaknT4AjwrzoMEe4wuUAqVkPqTF
6khLiok9zR95184i9KKh5HhFcCqX9YkwsSl/2bi1wbiGxiJ1lNR6XrfyBqLzPHE3HFctMJt/VrOu
gQUbnzqEvzi6ftKaHjxa/GbV03WJPG6+oV/UFdlxqWhfs9nKSnXliVcy6qhbIeQp1XAt62SW70ai
pL3i3ovvZGhp4VyOKhDEOcaUG5njyeQ60FhYMH/rH1ENlL+GchzOAEva9biOqLsHZZUUYzHw9mMK
Ea62uO0ZoKQGV+SEEAKBxgCGAaW9/4UdDQJ3+LRHbKLZqe+9t8W53x1afE/863bTHOkqaLDT6B2B
Z2N2VQlQ5ZQkNAOkIRAIJ/tpwoXNGZSOZ8TVeEbjJfgpdDnSe2PanxrkfSKCtdFEn8Urf5vZvgoL
9YmEcwsdmjZjrauZ3cCVu17Iok3tE0szXCjff8GRetr0fibZMIwQ49X4ncLNGaOSDQl8xjgSCUHn
v3igVG8yQhtKaYyVRGeAsZXsQbz3E+I0fGIMHI8vg83/QmTE0CSOqn7zMO50D0QQ+qkJEJtJwaAN
a7u/ykVPJ8/h/d8AZMCVC7lM+gP7nhqWT7jz/+LaUZWLuh2NqL6txKvC2ivrBmSiJIA7o/ocFE/E
NiC6TXbV2+DNlz3HMc2wtQZg+nxga0xZtZ9xg+R0olXgtlzfnPX0WaG10kCdYTEKlCh/ux6eiVQx
vmsYahevsufLsRTj9KH2m0HzfpkqgXs07S6Qr3iN7leO2ajPH/kmKAgXvC0Kgoj6SCGGxWRX/BwH
8kuClC28R+Tahgob7xGT4PH86WCXMlFmhS79WkcKfgFneIRvucJ+8F9We+jvJUtaVzcI1mVO4Ebr
HD3uzKxOjH/xtVBUXfpOrp664QQ4JdkNloLDlhTWfNU8FUMwvA9S+JkUo4EFA8Shkg7buJqtuUAI
q1mlC8hu2rDUujEP2PjFZMlliyRMBxQre8r5IfUc15sfBdPgQHoJM14wjeFvAr0pRCWn0PpOYBLX
ISYeXpB6bIm/0QfRsKw5/RcCVfZnzNVasE/fEZQAjgteygA+xMIhGFLiupwi1fsZUauw+QBhXa9A
+ekU2LJMvlGfEUTXBdpD21khVOpKpTCFjf/TM1Iy6iuf43IWDGiom+nzpjwU2fYyFA1fuatCOu7u
cEYJLAYGnO6bfLT2Kal2EBuOkusHOSQJ/i1aEPTIJIGKIkOAVayndnb4XDSLrtsxvZKq0ZhHmgT+
+3WeKVtrlfKWaUbmIu63DRXtUuP2OIojArmDlrRjI/6cxA0bpy70J85TvQCB63iWypfEYrTJg8oF
90A71zrlru56P6ze6iblw40MTzq7/xvax1KTbFcaUogrNeKKTspq68WSQBxvs19RknD12JZR6jhL
vqvhTp8rDL3+++BK2gEv8u3O26yaDSBNUAqOfs84DXpErdK1vhCQ/za32gQ9n81bsTqmM0Ziv6e7
ivf68lBanSZZTZk6J+g34CwBWD11dLUEJoo/TYhbdVy8ARVUaRVIym3zRPFn1DzKjmydCAhwmpNq
SB6FZ+iHfOYCWdut2jzfiKMydjfme0i8RDgSbldv13OgLmCcYT13oRuMCfAcAD3z2T1z5sQlKE2q
zcerus/St37z5OAjkkuVww7GaJgZEnx2xuopEVi3NpK/9F/+127D3ecsRwIAj39In4Invuc92UtV
yxY65dbbG1z93vaXzbWJGoRXgArf8oER7clsM6W/4deHoZp76RAS6OLmgHt8iun69uhEV776DeEs
SxCJjuaaA34ePnE4wjlBBGcHG/NjrwgqFxDPKtsB5OcfetFmv78PqXZgCUcH8ilAKtjQrt5GO7g/
nRA+5mOki2ZobqQG6ecXDjkj3zvJjaEwbeMaCGk/vxlJipa3xXSKM32g6IPGiuFnch0yuJc9PbDw
S0cwhZAkGXOIPeQeognsBxX3RLToCDVJFtTTgKBDTuD8npIlNuyhqVqbvc8fjwOM+BUGVlI5tWaV
uoSYuMaqb2f3OfcGqlGyoHN4lsDnPSLtx8SGXg1fojym9j/5kU8Xf0WglMvGsVhWpyF7fecaNwhn
ostQc1SeOGqmigkISPBO/W8c5lWf04WxQ/2XvboAub7wJuzi13TeVoB/3rMKVRS+45ItWfAXTIjA
bPMkYUAhFxhaqMX/6aJp5U8IwdRUcnG+JU1SW1E9IWw3sSsKxtUSIK+Pjz/cLx8xJgGPqstWmWZV
wymKKW+bZ5ZHF5ASU3DFsS0aqCL9V7TIosq8QnYTFboJg7m8XSzGwduZfthyTFkZ18l5yQPGw8lM
XWuzJSC02R0bkbNd8jdPIjWsp9glos/pICe4nGRciwGKeL7oSHP8YXvvdl4jbnR2021++Z+egHaj
CxXQlXQFGEBDgv3lMYiz9MrpHbPoZsY7m6Ho5ss4TUym7eN0crc+xMtc9BmWlv+MHhotogcWfY1X
nt1x7q9wVe2C5R5oDDewdRrvqsMoBfMsI6pfuSlAqLmI44SSMQkIv0gAa3WX4YEmm9U6/k3u4V8/
bhCLgI5C0QJZBgt29JIUwYNu4dvu1R2p9H4TNClRWgNQ7vabF1zq9GiNfNw502yWXYBkR+d1ymbc
jsvmTo6INI+yg0L8XFTR1ACVJryV5eKv+EiefywbMErfBklyAVAe+mRpLmm0Ko4JjrAmB2ck9/uB
U/2ybjmv0LFvU3wa59Br66apjzpId0f/y6gEvuMG8emDrpVEfU2hKYvRhgrc1kwDk5MH0nqoXPO2
xak+IGcIWaQ27GXyLFG0iKusP19IazJX0G9VEpmgabCfIDKsOXMa3S6cnuYtnOYiLvNKd/qRjf2m
Hs922lbx3Zg11+LZXB4Kwm7VEf8KsQbFZ3XJhK93gCsaJZ9Y8jC5h1z21LP/qeWR61Zje33nJ3q/
FdZ62FctENobwhXbv/SaVWq6NoBBXERGrrPS8BVYFtByMBA9TDmEOU88naubdUEoBihSm0E6m5fW
Pku/uX/tHVwUk5zsBoS7MPEv3qvTUNm8hM3FcF584ihyT3yEcu8BRel4mrjtwJFq9J28b+vkLC8a
SjW/s1rMWokEsYGZiZExlW3nCMhzvqt9z/aNegV1zi/W5m0e2+yw3Y8BjvqJ22nbZ26QlxSF1eRM
jxNjLEWD22cZKeUQkG5k0q2ehvTpD6N0VQTaloO8mizQF8nZ/k94uEzCuJ4yH4u4zgkqXVApl0/9
AlxskiYjubmumnqowgilWLXdj+ZGqNQIebHes2BQRr/XuC4vdYOqSd5TZ4K+LccqWSdunLk3KOpR
gHiTql8qkL0VMknT5esCSHhcxByJIEF7G5Ixte56ZNtZJ8Q8l+yzJ/fYqpp9iyA31SHYj3HLbZ4S
1d8qvQDxms+4gpYL9AhJZzu61RUI4BKrjrjejSizPxFI03fw/r5N6kX4v/AK5RSsEaycvV21mw+v
rsz7P9miKqrexmxfl8Bbnahm2SdiKpQvGiX5njfawi0naxEUzRNVj8V3oVRsCfsYImOqzw646WEe
EE4riC6MANBQudimeE76nqx5NOuE5nNMxtYO5mGTH0uRiIXu7I+Ghitm03Oi3/EbAHkUx2pAS7Aq
rO6usOt+4gw/LmfKu6mgP6oQLooT9WxnEDefk5jdMFpyCBu1ocJoA5Vsk2K3wkWE70QamisPdQc9
Qv5B//a1bZFCDCbF1v+YyKy/97wnUGm5AnqpcInxPavcEQCg4OQxhbQQP194thm0MHB7zjyTMagQ
y6DWDQw99pFoEW8G0E9g1ac/WOPKVxYYIltKaRzpAAhh1GPfVaUmUKASAxFQXHWOqWW7FRZhifgF
++4vLgDkVc9dUUHcPG6moPe3SOoz5wcV+1qq+unlz267awpVvWM7sZUe7vKyWU2p2zLMvU5nDHlU
OVKRUf5MhaDAY78Ko18TNWlugsVYgG7r+y9FKV9LJX1oiCUF3QcZ+QHbPuKFmz8TUVlRMfBkZSGK
MXdpNCkD6WNeqpfQ1Gw+iNkH94yZp5Pptq389jNQzcb7xmSevMDF8pa29bB0PRpzMVAI1M/3k45u
f13FJsDtfg05x3FwcLb3BHFKW6971IGqS9XzR+vqVo7pS/fRWfmWF1TIAt+JotxE1iV0/YXgpWnW
zgzDIhzYoFvQk8FSh3m+mPJk6UTdiItPd7rrQHyT3ovuBX6IAH/bTVZvnPJh1pIRUiIGEzidBANy
v1nX8tNwC5jW3Cgw84UaviqZjngNHH++fwQzk1fVQCS7UJqhhaRLQGsasYAu+H7Y23DBEphDbGol
BBoeUzcQ7FokKiTKzNjCkU4W/OYY4Wk9baa3RKGYOCin8Nmu1cN1SmKcjZBG//d9Q1C7u95GdnHM
luyfU8U3Y1YpiFGanxA8GCXDRDh3JtpLIDPDC2vHZcBAk+WkSI2/1SRLRMdoLc9E4moDjCD9zAYb
wT15bE3S7giyXi9jysKmtBvzQQozforPLmQjc+h0F2YjRz7T2yvAmCc3UiocpqKQ8o/89mMjmnCK
Szr1XporuBVTT4HTqBblE7ZSqnDHRuQXIj+AWzZ21hkJDSeAKR3lUnBZJwaoLME7pmYU+FNh4cTY
MJjHg7+Kec1p0lrE/p4EZ9XlZqyb6C6/oaZuf9+hlXcvAwyJII4vS8jwvixKHoMvt4SuvHaIdiEk
fgQ81R09qCRM7cV9CQO+Kzwtukp7ddd6Mok9vmjKeB2JxX0W3II6p9b3pKq5djyCgeYWA5KJnzLq
c/yQScE7rG4SHEShZ2O/hpxzBtWB0lsStWLUaiOvGyVyVrUUvS5myotEieOJncrHVlC+AJBIh5o3
i8yb8h5zHW93lck7IO1RKqpK4m7G0r915CqMl05b6O7qiDMO0mKyvTusCEQCy3W9o4N9Ga7in1Lw
VJrxsYZ/RwHYbr0CLS7O5IfLvY+d2qZ8FV8SBc/Q+yVTJiA/TSCEtRu9a+cq1oMMaAnd/1MBMUhN
nAY8iCXRFwNfi+J2FYpmbVys+De3EWpS5duKiCWXyv8Plc4GpsJcCHLmgZvIAxyM2H6QtX2E+yT7
V+7ZFq2tbU848nQ3c9kep2X55YplzcHBiniuHm8rVgtQ/5W9jgbapjpYA6h9UXt5y1RiCSmXVcWP
bWTsZTz6lGo/vIAio9A36KTUhZ+M4+dhLYupKjxXAMr/PJ1u+6k0c9g7kugssl1L/SNst1VqtAQx
3mvNBaa4YVzSsA5wfVIcQvief6j+Jh/QBjDoxCWUOFXOHdzD7hngyqfoRGNUrReInC19zouMVBuj
hK7g6drgkIwvq5NhRdvAMdz9zylDCKDNxsRdbe2rhH+NNq7WvrkmfmaEI7lYucuocR6mNW6WghCf
bcGqctVAbwg7JcijrUCBVfa0J2Tw2VvP1gddteVteIY9ke2FZUjemtgQyPSHe570x0kAu3P3BZBb
quwYmEBLqRtAoNzeel4HCZNQwJRIf4JrpPRIuB9OeLkUJULj4RVjFCUHLD3ynMf4HcNYZCELJLa9
jjKn+rcnqOjbgC2vAzYGsNjzi9wGUHm05WGC8CWT2UTjJqTj860qA/SHZf1sPI3m5OBRZgAtK9f8
fNaXb8Buuuzsh5DrAP6ui882EHz57aW5SvrS/aTMYcwYWLR7T8bHDCuLyrBvGL8k9nEiVf8UHZ7y
IzXrS3goL1wQb/gpq7plTqno3B0KCIl1evPWxA9xDI1cs8xzZS/FuslECxvsraRHClYu0XhRsPFX
IR7U20bAP+s/CYqvK8D3OptQoWnFTmnzFsZh0k7YJeclXKKNkfZ6u+gXcWB6NgAe3geJip5CFAcE
9ht8iVrx4GGRS4TztI7n0fpwaOLucAD5VhjU60IlErP12vW9A8sahF6KWvjTAkCMsLJ3Kvj3K5Mb
uj3Yz7+wbL40XsiVn83vI/GOyLMy7GDoKtlzk7KfGgNRWg6y1MK0i9cteLn+lI/OakbRxsNASjxb
XAgnmbLnhCbw1ukzRZLoVio6/JxgKLHyuzinw+19cwgLEu0OtAX+c0H0DQ6/cCldyI5p6mifNYfN
owSGvAjU+JnVMNolOHObAf+KYmMsLkpbRM2DM1rt7grJp3bW60WB+xBIe05+9jiumx/PK5DDP4A2
WKtb9VDZRRvTClZ0le+utlx7SfbA5inmTrEC3yG5pB02REhk3vccgBcYf/dS92eTFO6NSGVQLJTN
rf161x682KNrqCHm0ZV87h0MNvGNDY0JOaUakgC2YHJ+UT/31Vpsn/oPfpu9VfnnK1LcGk+wZX0J
WEI4w8pBGn5P75Nj9uAQhqhwueQ73SClF7MH28GJZQLpeG87NBuxCRlDIKT4L6T+UV2/w45Azbhj
u5R2ePYwr9xb+Z62RG5lrG2xYQr8I3Gu6WVC0YJrTGkazVQcTqNSUQekYpMb8l7eNyyq8jC+Bnvg
rhw02KOSEYl+pMDIXcm6wuvecMkEYZeRN5qNJC4DD2lSGmR2utVIbzXRXtDKfolxw78WleZa2k77
u119BVyixz0duemXq5LUQA57dAX7M0zIn/Pgy9h/CA0hvwOU6o7Wc4KnOonzAT5PYLUzfoLemQrg
oDQeQZ4bEI4+Ug6RQyU6LQTPnUDKCbwmN8L1QLlLNMSDOE3bDowu3hM6HMFaCAN8iSgGKXEW07qd
fhxufylntgL1VEghuA186xRWuFCk9aPCWyOI3NjnZ/4PxDTwCHaEpnDv6HIW91AqARAuZY2y5pwe
x0wlyANpsxDyU8ukZpX8xwCHESfzM7s+lOaGkqToy5QxDQN589YAPaahFUaTwdEeMBO+kJMv6eGE
FnFFP0xhoC/sm3HZhinWLXFKbtiHVreo6BuwCVOSCA4roNstlhEhnZZ0VSHfCbTCtapzMyNXhSMY
lpPKdFVTQj4gSfxwLod4lIgPmDHdrWtuNHt3I3SNP+zWC089wDokp7J3xqIa5cGlLn4AWNnZMR2Q
h8nwKxP4NdF60xYmJEEqEkRjhXjey4W0RULml3zBPLavZNNhttmjXRpSy/2OH5AmkTS9PI8Dq65+
s3hHJYcHAqzk+IeeGu3AvxKJYOYlEmYUUo4jv1WXbV3wCRqYOynxOFkWyj+aff4QPQvFvnT/OZDM
yytIrkZZTKMYGSSM3zsjj6gLM+RdcmUWvWVbw9YGOW6By6PXCo7VhNF0xWv9imEK09Qn1MXmAHAd
eygCVuaGhE3+eP2TujitXzh65QB3JndSNNXv+RLAbWBah7B5R0gtF0ivbZlkGHBpUV9X6up+BJEF
yDN9rHg+vgjsxsizp+ZW6hV+s+7Kt2umOpR9macaOo7oJvlV3ee3R7MI8y7HBKY8zETyxkcOOH4E
iML21qRDUf11am6YOAntMQs+TpMgxAJKWeWGvB2s3wZoM3DWsBno0lnIgUIGFJz04xrmJXk7xWFD
JEhwMlUYKnKO6BIZCS3++7eI+HtN6TGsDBp3yjt7v0LMarpOdL2B0LHVt5uSI+jzilCtqG8cIzx7
ZIuYq8yx9oI26gqseb5U3ucOErvLhCj+s0UnT5L7laKvie29MVSaznAmSCmFk+txuXE78wcQwhz9
8tBDqQG+38n2JODWNubLotkFHTpKs78ICDfsoGICwfmT98nsW2EIsaB3A4VSf2K/vOLYl8VFbGYV
AqKHTA02PC9oh57/lbKkH+HP8yZSf5o6k05u6NbZb7PyzFQZk8SxkwRN9jAu+35NvVoenglViwO2
M3f58/tBLCOVgIDNw/63o0QXJzE7oIiRzKh/J+PjRWJkfnHrUL5J7a562JMedxHSTVvNhwAkvnGR
B9iaH0Pt0zwSqLWVaR7rmD9qnJtTNJWrOu3u+74px0qoesonJxfYOGZ+zwfbt98Fwleo8/MlaBBY
E8Na6tSVP2dyQcU/RuyD4iaWyXl6q8RBk42V+XRQ9AmSc7XzVj5NkumacpTNYKGLb4wcRDiq25V/
OiZ7Nc5agot6AR4XE8CA04LCtqBVYbid1JhmuDYkvqXjjS+tgzMdZ9aAxM1VJplKuJpSeMnly6qf
lCXp8XvhBYSbbn6ZZsdHqkZRIvL6s7fbaEaL2dhn2ZSZr2wjswBnGiXLzfUaKXpGXJr6nc/CCJWy
oQEXFEauFaiUKobD7rXMSysBl8GbuktlK/SNeAcoJ33At+xXDKj+gS+m4Z+hsEObp8KFqWsnRGZI
Pa/PJyF8lmr/djBASUGF3gAXduZSaGw9vTFzGhKMXEjhhEJDTsp1SNLBVa5wMyknQHH1KIY1p6iX
OQzRMqrSVZK2KKysn2L+vag5tEtxsRMuIVkh3TUsMHu1XgS+1bmDF/oWj3r0SJ6PcTldpu0W58Ec
d+rtXmb1EMU00dveuDYNfFc8kuHKwhv0+uxtWZDv8NOn3WWzLSdvoy/BoHDrRJR0VNWmIYbr9QTX
VR3i4eXv5J6GCTPOnRXdqeS2ld6t69l58pFRAZ8rdleheKCtkPwqKHyHu5x/VRibQJRAlCFZe10y
RLqdn4k/AOEH1bLH5HYXnLA/yWkbNGXzXCbFmeOw2d9Xuy9W3WfOytcGmUHwRD5B1BqmvbqFqOcI
BSgbVM9A4g2IxoFTbvwTGoCG3uYE2H2kJi1INKKPV1cVjn/2bFJZP8rBOVqzLMRYP7I2i2ybu9Yu
Vcn+NAE5+XNCle/40ATO6FqHSmIm615rFrHCq68mZt8Hopon1WsN8xkPOj4Jigdf5yiefUnQ1mhj
M+Qn1m5MxKqXpuxPa7/CKCjgiGzy7oaKBle75adqge3f328qn8SOceLAylMjYfW+YIEjnWLJf3ov
gX8L5lHn796Hl2A+xSsS3xfduBedZvoBhzGd8lXeT3p504eXSq9TIQj4Ap8kfK9X99gIKwXLNhZP
YKZtmNRFYvQVWzTUxY0hQ1hmGsHiY+bsG+SsN4GH6BUVGqzzLC4lrDXMIWLsAXfzRNktlBR4/P7d
QBBB+cQz6xc3NSlKjqv+mzdYQZ1WfHcaUfDhze3ZSo5qXWDgk5YYis6Zbg2/Wapt+PLTeGlPDA5k
oxP/ZfP0NvWwvMhWjj8aMBe0GTBAEwE48zT7r07bQrRCsVK7vrE8eZnBW7sEsgPE/hTKoFnwNSDu
c8f9sGtL4Ckb8ZggjPKAOqs5kx0wMukEqKXv7+VYsrXO4j594VHNaCbRgy5oa/99b3In03YkUcMr
sIQFQYcgNPMobH42CrC0Vi+pCTP00aAU8RjYfRXUYgVtaDEymKL24cIbCWOcNt4FhK5E4tCzznXd
KQUYKTN3N/BuGreOsELS3KLuWRf2E06QbAQ8J1rTMpRWYKoHIkTt34WzwF01KWTl0ms+mRvwUj7J
CDqvn1s0UV5LwV7SPuUHl23Fi70DdOu6yIV2U8Dn+aMPZ6zBkk+4OfltjAt/qLh7Z0G33GFqLVoG
TNSn19CRc2Sf9jFZSSlLsYSSBPyvtNs79+AQB3DtkWZXrA82kxQ4s0X17mk3LPIblyE+kr/f1Cla
71EGKxsGX0ViMmYyb2LTnGo2N2xFqQxPKNZjPYWcPeDPBK8KV+NEmVl2VwBI0uUjqiZ7WpNBgQNa
EBleZRD4FgdBqUK+51ON53BAHjrrC4NJvfE8fLLOWBI3hs6ei78XrWwpByzrOz2ZiNhHJ7gw/aw0
Pf0wXolKn4q5fM155m+oqo1P22CpMyNnGP3Tntlr87T/cjMcxz6MWuicnEVgOelUQPSLWNbttwoJ
dS3F51AKcsJtuFLSkGNHQfXsywUAXPF1ODLGcnzMgrLo4ehOFWyGaisRQeYxsihBvSCy/U5XgeXZ
KDc7vbroM7vSZDTPWD4ePrkJeN3wmnol9EyscI7TQEXuWZY+UI+dZsKtDrcdemWt2bD9Maih0+mb
AfPworcmp9cymkZmk1OwO519kreokIRgs4njSySxnKIl8gUH3Fls2OtjKEAz1EULBuSAtcgZyGCC
gT1SPj446399durK4Rp8HAluq8xkvbJnO96+6hdaXPzueP8K1nfs44l4piKuO7t2N1OAstpcvRA/
TzBu/zQWwK89ThKeuHacva8EZaGKoAXxQq57G2RkkUXA2GPX/Ct7OhBTQ9ldsY53yWyubIQ8ytR5
YoCVNgvATH//ycd6iAflxVIJquO4u0VyvWakrvI82w0uj5ZARR4QryUD2/zUlYnM36/18A6wfwSq
/KdYp25oYgqspea4e0Yko5CDlBW9IlAA4OEjNf5Zk6ORYB7DHxYkf7+N7EN3MJ9phoKwbm43TDb/
XItskv6f2vtk8mzrvs2/9nI52DHX4772U0UArzSDHeu5qUcyvYek4NxOL/ri3/DuBmB2LEFV+IbJ
ZIxvPpYGUTSx1xKSWXCheHQrQHeHTtdZG5gPkiodL/9lk/5tO8KcwWLb3VPrr8tJPqKlL9piN2De
dGjeLHoIsVKa9aZDOjN5uJOeUZLVef8We7IiGx6qVxTNv+GigiTuYykaZgZk1m/vHd80tGvzZ9av
7QcDCcZAdy4BuVuEjy73fN4bClXrOSWW4Tf81996A/GF+DMaXbN4ihYaALCqqBIznXBH9ZDDqUnP
Q/tbuYywwrOBwCH29S32VTLEWq1OpQlPQ16Fwo/fsKRwiT+2hJurGZjQMfjsquOnPuFX0RHHcx/F
3ydvNqaY9jx9Vq6RjeNABv02PsGNQKAeEWSyyapl9oWNJF9jPIkKUAtmDQCwwd8wb+H288eoFSOf
JCwa79hqxOaY1wIvFHIMdy+K8TQvazFjvoENhe0TfUIlsbCyrtQNdP6WkDv1RympDnnvCaFyiYJ2
AWxIc44jskyDoQCmIW2pgkCmg3KRtkKvkgXpelfzHDcKavg73fDG+OWKGbFdTK2kUurfq10dP3HU
fYxvwSM/CYlgEP4klI0Cb+Crge/4I1iSZVWtTdc+8O40Zh0L66Rcg9o/tAGMi1IbSNAHiZ+K0aLd
ywMEOHrSRb19WrinVBWOxLb/1jjAVMdj0xbzAgh2hz5g99uBWg88a24CgHrRE0AIeuqysu6reYkU
5+LVZ8/wJfRJxgJdpr9UpkjhmxvhGVmlTf178LfxXawNJc6g3V1OdMcxq3iNrm2GCoPw9AiQc5W8
49vmR3f2+wT2cawhyCYVUNSCr/+MpHIV3T/VVv0TC+jrSSIQG2yLd83a0GXExyFaJN0BQxBHPtO6
4Bbadyheennmr2THDTKTmAzXQwY37Umq8OKhSQt5n8sAIxOjSlVLoF6xLV6BGlu47TZFhNZuDba3
OtepJo9iuiSPrnvrIqL6RdeYZO5/atucVu2AzXSxrz50/3zN9ehZ/YgoRRzZZXMqexGz4S5KJLT8
9IfBkP9rcEOqgqqI3ibEvOx15U0RUMaeTmCftDQwcVEhY0QJlhv44/QQ5wonA9v5rRhP+GE7qU2f
nsCPuT7B+PfgWGZrMyS9KdVzb4bJE5ZdY8l6OdHzU4iBH0Zaah20pLpjUWYPhfIVB8o/Dt4jE57p
NgD1XlE5zBCkW4j5ct+eS2cYjGav9BMBJdzQfVyR6bIsLOJE+O7Zsc5m4ezHnXX+e2TYp13i3Grv
cTKWxDjzB8ec9pVAnBKbDLt6TzsiALrQtfSsXSeZWMKdHS+uhJMXVtJGnMmwQdZIHPRsOtUzLPAq
B8osJzcMOng+fepFNjQ57BQmI3XXzY0nB6NjL5vUMZVsKar8y6HS6W4dTmldG/Ir05T0L5crZzKy
lsmtvIYwjsSLcDXL0FvuSEccUXBqeR2wb5CEZzt6kZ+jNR8s6vALs+xdDZwm3l8vKCdukw1cW2Ja
5rR6bQiOKvlWxtvRZQ3bEp2eg5CYmL0ipeNMl6X9odL2HYMpsMfnt3JkjnrpIZvcz90cAoROx3+x
Auwl96A+cyclcZf7HzOVfkmOKW/BSblAyu7wVa6nPRtfdH2dljk0VNSS5rqciYmhsa3TmDfna1Ox
opmloc3mZVPLfV+DHEhANdFXRajhYcPfcH13qFZLCdiarRvJ23/k9rhJsRL7UFOaVIe0YMTyEkv2
M180tiz+ibhQoBY+VhtS7oSOgiI1rJLdDFXRvkRI8kMx8VzIB6C5ib/yKdopb5vv18IOxtjdA1Qk
ktZklxoWvwoE08+8c0A/2it58O4Y/V0j540W03jK1o8cyCuv+CyM+XQuiGQmhRguEnYLOU5genGn
7cFdtJ/HuK3p5wTgnC/9LjDQF6btToRcE8EnIYYkWD8x+gV26N8G4cYyByiFmGukk2OadxKR0gfK
kPJZ33FuPYlYAdmV++uQQyn7hDRIgJqlAF2NrXI/yFPV1VVTSG3xaVXGPYYnHgngRprd1PopFdmE
8FViCLmKBgolfLmT3sSWnpWrqAYNDO0ktCg6sTewCPd5Rm7h9V21E5T+mHnogdVXo/KI3+NUKXNZ
IEzL7IuRjdyMbCA3nhRDl5t2IbvRSP8ee2Lviusbzafn494RghyJTxNBLw6aNs7wMTC/UjAJoKyn
AqfG88x5mQ3ImOJODfHtYLO3EOsWMGEwC2X/FM8hat2Rr2hTNEct1pek/xpSIBUpSjqoFUfWtSMC
xiFdlngH/axT8O2pRh3zehGEJrleXvcU0YccWNENDLDI/WaPXwItD0p6LSLGXY++V0enhFEGjs43
/ify+5EA2Hp+JFjrIBEYUPCYYVtYER19mkgctmAqYilc+RO21Aal5xnHWto4NGa/7L3M6PIKOJka
B/itO6ZcxonU7JP0cetHU54+LUAwl+r2j6CZSfOTSmFMfO/f0JbjmikbzGCxiXSo07UO4k5J5Kyn
DuShFrSEQrvEb8wqDSS1v/ev2WKxd6pgCJCMW+7HV5/4Sq5meC/VNAVpNVScrCnSYaXXbVtQRMlp
yfX8p+uTani8xKY4I3owLQlgHwZee8Yv/AA3hc4xW4OhlYhD3LtRdD2ikEAhk+U3+lPJFlW+SkTb
MeS8p15XIHw1OQiuwAOW6Ly35lFPLvrsP7TjbQoV0PyREozdvnVPpgF8rlsMgNwWiRyWBswSXpvz
bxwvL50Atc8Fnz6B9rnZyTcg2/8IrIaZ1HSz9i/H2J9+WOAYhsXI0R10irKu3JvdFzNxko+kEH/E
iNBpP90MeYcX/tRM33SMECAHDj8jcqwXU8M13BfTKlVzELC83J2Nflktq+uEj2xdJ6a0uao9z3wu
RigBhmOJkHNU7od+fQ3KPa26kvwly1q0TDZiJ/zLG63BcKEnK+pNUsfLVGqcAMl37+m0sLn5D2Wh
udKnEMVKLrZ+v3z5acOf06J9gKAiJSAYmgYAkGrGKjbf2juynhmojnCk1U3dg4jwDpnGjOCL3CcK
zdYFfNpZAoQfsNLhZR4PxIwk94NgpfcN+09Et6stmzwjjftwYxzlVZLQ4sAloMEYu0wqQo5owbKq
bs1Zs6WNCviw+CEassIx0OpvlCXGVt9CQn4ClPxKnREK7VxFoMRc3FxhMz4zlXjmjfmR7V6ki6of
rxTAahNxZMvn5AVY/aIlSD5ZfmHoYbPPEAjIJMZtGWV+o7MiyO5+6Xwx3TLYNCpRMGqGZYdKOVDt
8be6PUSnz68rL5SzwNKTYLyg1lnziL8prLHFGgqH1b0pDhdoW01jUN9Il8DjPwjp01I98qF9oDZW
flVnwwxNYWytL/2EV4OTAVgJTfhQNZkzrEoaFYe9Iu2qO214VNfo0iqZG7OEya6nYMYkbEyTzb38
vmL101dB1whidjKkyZk1xDKyUezAG7PDWZ0Tv+atkD9tWsYJXU4eOMmYckvOF/DN3WJvCT97oMpk
zOx84uELxW2z5np1vSRMEjVjCzx42CAle3NGtZhZCr++OPRRwjuVEje7gWLla/7ACNSUPwFf0uz4
+jlDXujRlVsLppBW6YU/QgglTgO5QrhrFMe/7FmuVf+JKp9QZ90HHZcLVirQRul/CmSfG4r+yEij
ALwfb7eWm7QTIV0NUIAGXrRtnmH1ega8eR8iBwPKHISjZxpqTFLqXDf+myWorDCAxG/x306bs1nh
43KDs6MplRTKXaZmhWcGNdAqXx4OEV/Pct1JzaZzk8jLmYHz+fjbZvIST+c45lOqne6H/+Ne1dO9
u7rSF5zeC5UPY/pH1IMb/8Ntodo4WLbOK5K+zu7q5rh8MWRP/sOCQTXzVJLKaRrzKyhsNh4QHnIz
DRajCynVQoTY98iCvxlqwERs7vpU4m8jOQM/Ab5kRd7oydDHBjSiip2P5ehdMc+fDHSzju5bLhNn
qlAoEVS2kAsqR1mpxy2Nh8TXnhYB/o+nUlW49kiCOTcoiOcLMx/njvKOWUD8kljrBhooy7H4nucY
WlntcF2mjfD1mIEw43RUyNqOqVBHDKXoeK5npfKLXdRL4vDTT42r7rR+6KC9kae7k6FYmJQ1ufoJ
f0Olg7uO2UOIllImlRZz7bSh5h48rVsqAt+3naj37o/MHKdTBlGbXTOs+OWCYMbNiQIs8rDCHyU7
DJwRAUe0NZetAHMDp7lJaiFUpU8w5ZqwPU5CXbKHbtuwKy49YSTzV+qXrCk3VqgXWyzb1+8WviKi
9avW683YrGA1EIIX5+bnEKW1HpW7Fot8AQlfAKP19sJrXyy/lrhosF+1hj3a+2ifTDiBKP+UXmkS
JQR2aH+qfWFJfbyx6UWjQ4qHoKVoVJ+QTouvEoO7lbmRJAAxaTdHn/g4t9AAtuY6sVDcT3w2e7JA
lktkXqgo71gHIW9u22u9SfQuriruingNe2CdSfYKGOvgUbf5g/wEy6oOHDB1NHw9jNNjNT1vtPsr
vS1+aogLHWl78STI0Djou269jj1oiDTvIYPCnrK5kIjuEmk0gy5YxULKRraRriyZ3Xd1rxXyE9gN
hrEE6mZ0ukye4grJWbhxJ56RJ96XbWmZo6APtZj4eWkKrXaJvllClHHkOYjk2PwXdVARJ97i1mqw
RsGnHq9GFp+/T0dlSkcov3lQpWf843Tg06RmgBBItMK42Q20J+ZU/8yX6n7HS9Hxi5cZA+5KrSaM
MOTqPnjfCPLJwsKyJsNQJS1iJacNq0LmZ2u5DnGYlMIaK8AIjIDUTACMMWbNt2HMJpjsVFINfcSe
pTzlwdM/meNQR5I0PLwvMeOcOOvjXTSjiUeY9QyHVKr1PX0UU0UvcgRn9tG/CnGAZsQjenIeNICH
Yp7OuCRt9JyKaD4o+Nc0/EFnw8D71VpXA8eiNJ3iBe4M/Tb6Zf92eUDzbfPe3naXN/A4NMXkoN3G
icsyMJs6dVjy9e0Cu//aH0o6aNHJ79Uq6Xm/ilqqnsjFeJlnC+T+wfqX5zjsIi2XaO8JSS3gMDjB
qofgZTLWk5jvCU55JBBKB+ZQNq2rNtTE9IBE+2sQgBs0FfRbH3PC2zBe4K2FSjmf+EXIggESLr8j
DHtjpcrS6JNnAXyCNy1ISRXtOdrLS2Mp6ul6IBsQpKXP79zrkeKXS2bIrVRN3m/1tFJxmtG15Owe
D4GnsU0O6KaJvyACZkDZfjwjIRJVu+3l/3djBJ9iZSS8jwaOCPNuYffIaFcQsWyXuVSbKLWycvmD
8RM9mFMaXpRSlMkvaUAL/uBuzv+ZQWayEns6Ud7LX8niV8YwbVg9lcQw5osEP5Brp2HyrIfAPQge
lE9nOaV0r9KeEUtjr7ohwOl45pacgBPtjHzMOERL/iW8K8lD6/MYSBwS34t7ae0NbTokDIhCjCen
1ZaLYIjqKCu4ZT4i9qE4ry03t3bV/7HbJHVKjhr0TB/ZPfqzFyb0nC0NbRpZMM3qLAgZvNWMjvu1
vlHLjKH0iU9eMWDEvPYpc96Edw/H9jyOOUd2UIZmDHgReirIzNynN1gaLrMzG2ls8tuxyFf3GS6o
h+7UNjhu3IfRHLFEWeokxw0gDgbnIaeft3+ACUChJoubrFVDBkihEqxfj581eSjupmWRynonIwhw
l+oVEF3+A5U9Ts++97UxxsjgLoZ/9/ypG8PqPoSj77P3b/Pllbkze/3H8peh2QTSst3xd2n0m8dB
WWDVM/TivtFHxWSkTn7iADSmfXS3bEcE5JPr8FOmngJGglR3LKloLiuvw1DLrNz8JBHe5zpIa8FU
mfeaEMU6bmHQCqH1jSS2wd864sAF4PKRwN/gK67C9z+rOVNO0+PFnDduqEef1flD8UflaXyjv1pn
1BPdovCGWS69FbIcQEPZhuNbpSMyaOXD6v0W3LI/sK1FofmFuYfFdRRiQMW0WUx+BsVkwfmPDkOV
IPvGSRj335Mg8eO4mvo14IDY1JFN1YKHVbSY1IarEOw++fIu2r+V/F+cpxSZClly4Zn6e6mT9W+g
IFms89MrSzobLN4t57Qxofhm/+EHALPJwQzHSu65CMJeEFkdAgzO2+fMp6GSzw+h2kg6s8pC69Uw
i5O2enZVFBtUfcstoSn93jS67oI9DN/nUsK3uUWK0QXs+7aI5b3qT+IubY4p1ifA6LgoLAnkkeQR
FD9sg/4azfLfr6Ass2b4lPPLkRfWhv/dj8FMgw3fMI8uIeoAhUX2DE4LjiayXy0GquGUBymr+ZcU
+Nh3cn+mYMwGlRUcdT3y5geTjPVxWjGw5pu8bA02p8QShG0TdBmgQspdUNIvIbgKgio4VU7QL6qy
+yLGfpDISPgmiV2JZxX1Y9fa0MaY7pW3m+4RL3Xo64OlUooUICrcD5fZT7xq60FMEuQjXN31Qof2
JWUtCozvNhKuWEZDOM/jHSdtg/4SDaep+F3s8gmOVfYozhAvW2aaNk7V3reY/MpssXtDwQENbmM9
tweCclPAaW8/6+jBsvGh2QJp9ofQ9dJTSLe/EKyhZAIuAtJRI4zZtZTmxA8hxo5JDh6Qz8mR/Cls
4xVHxDOdQ0aSEyt4GLtoZNQfBppEZ5JVGZiiBZiv3dPti9p/KH2Amrs5i2pOS/JNx7JjUJ6Qrcnv
9Pzo+OEdMH7E16ENcTYAlQex+RJwc1uWw1b+E/Wbmsa1A2r57JKnXO5MPBWfqOeynwt6vU6UKOl/
JkJAqfNoysBPljSY3YxtqU0tVq9u4o+tcuUgF+mXSBkKh3DH2+4cXE/OABjiNbfDL30KkM+4OsUe
ae0FAd5MvArULAZRLje0GNGTXGeK/YxhSBusVsHVY4tWkVOR8iJiv8QWJ92jgdyjCpeXsECyJINV
bc4qt/uVcUxF+JyvVGmRFYzibSroCL2HIbcs45relworh121SoY+iPkLHSskty6xhy9iWNzaHi+F
Ox2iEwoRmUmO9mDDhUa/kWf58aBm+aNNLiBLYb9MAeU+p9UvgUvL45pBVwcen5M+CucaNBokYxmp
Q8ZHpLk0pF40Rjqxg1OgFBzzL6xj9Q3cfgSsf3KOyVk1Bzg8awuTAHeof8vSaDQp7RBZuP2P9/Wo
n2rMVM/DOYfCUe+1o8Fo3ylri4NlvCHnRuS+VJkO9xyDaCnpZj8Cse3E6wzNU4c3SOTbhHzPFVF5
dmhHlNLXR5rRC0nd+Qte/Csv3ZBqvwN8RiZeWq1Az78qpiA7piHWtXixl2w60hvVz+o2MWGPeeGS
Qibjp4gKxWh5/9PzfciCmg9SUq/4R7moqN5gV997Ap/z842AAYNeS1slolJFJQpQKWB0Pq8yTDBK
yNAIdi2XLADVph/+cNrBpsOkkIKecQHsQDs2kXt3l5gT+DRfrA+9EEsHbLLJ7zQN0Nmqj8NIZ9A8
ZteZUEIUvtXsZGStT26LXzd1W4fWl3mjEePo+emxmpFLWde0sg4em2x45qj8w9pnwl+d0+S3VSvF
E6zQdkXbWBefoLgHsGPcbKBvbg67CctzZ5LqiMzC8i7S0XUuK+C/IEQ9Vn4RB/6UhHloNldn6exG
FWHN5b87hmRYQw6yxrI8PElJ5zCHjx/pPNOFQJcD9f3ZNogWOfJBNaGVjF2kR0deLzZRGDfMU32v
x8qzCCZbwWqIli1DXcvYvpZndD7OEfbYFTKiwaJ9/HzcqpolfRZQXxd6sQP3I6gDefVpq9Fp9s2H
JCQ5htWxFAAQvLVPykqmoOz8Np3SVCk56JwPSzZWRLBGDgBHivXVCDJhCLSx6qkR37NwFUdPQYZc
uz6T4OdsLM0Yyzw+E+5L7ww+fh5bC9G7c+pANgZyi+JLs5+SVltpT03CJ7AasggzmFE3h6k5GfvM
TPZVdQs5JC3N86qbMn2qgGvziEuIWQ19ZgU3HyaE1qLoLvELYffZ6Fo2GwivTH98l6Rf6xTNkv4n
XCjqg1AUetctUfTfXXx3ox7iIlY1WMI8iXvwX1HhUBp/zXchjwVmS+RuxS59wsrk1y48WFxzh7Sl
Qih4TXtRvWrqmENRWtA8aZrA1jBqoyS8BRLGBxS4sUPVAgFrKOvlZYa6qlgC1HhxaxMGhrbiQQAP
ecliY3SqTLvvihjf89D9TT1kLFqRNdZxmoTcyYi5exTGp9ApzU3lqzn4zQ/b7onde8XaiISFpKqn
8Ocfql00xVLBGSdR5k4mCGZqPHLVFSqdRIX/8ISKTmAvliH+Q0L94wRXTlhRiWDhZhwee2IgwbaG
5aEuHmxuZE6HUB7PBbCJHiapcU9dJAGIbGbYQR0iPWOgY/gjhJU3/bs/GGeMEuJme9LpLVu6m90s
lima/KumZKHi9gCKEq6btg9VeqeiWEYwl/GPE5DP8Qzja+ruuPtZKYeTRIJrTLSgN6ZOvod7dMxJ
bcqgdOLf8Zh3XZXQ8nlJgG42FkMbHHdOyYzMMyQ37++7rr1rt4mAy+6qFuHZnqcJVTcwHSgSVJns
EgT3W0WKB46AcFJ4cWeMRjs0tZEmQuiqBcCo7uBVdmXv9X7u3Cf3XZ+9jY5PdYelPzG+X34LVvQX
LaLiMwaXHIK41ibnf/omywjtdtkEnbFVk9Ln899XnGcnI9Set/jbcNQkLeSRWtkcOTl/5zIYHsLA
QavqGC80U96fP9AXTj4XFt3T24/8+XXDTLrsItuC5We77MCc4Yp3VXXuv8UUxOvlz4FC8bHLkSRR
C3n0DQAmBYG8lydDEAmhXxDcP8AFHCcrZMAyNkfDHhObkis44tMTDuRrwzyX0NleJzkz1PXw8nVD
3Ccl/CcvXozBsp2eo12vPjgYS33U0Uu30Av+9jkLLV80n2FQW+ZmKtF9Xf4v+0HFoJL18BKwruOk
ZoOGBsTGewDuFPtab6WUWWELoPwYMMqhsIlOePkghXLsACaqqEwStSxk7zezAjzfgp+hUkhc+K8m
fl5SV6kT1DN+hN+dlNvL1+1N9ix5ANSJOAKUYz+W86+xcDmwr54wVm2rubMFTWDkn2qu5y1183y5
U5opV6umU2pIaRkog+2H3BLyPSHiiHSzoW1WrL/XdwqQp2dLwmPZFqfO4ihuGJBfVrOLifCIHHlu
A0fhbulMPckQC6528qNPQ8VPiEyt05D2MKPsM5aYnkOME6t0PKdGcEuGvBzwrMQwbu12czcWBDAK
vjp2/pundT+UVzY/g2LG0KdHAsrh03AwvkqHQ5IOmMZIG57KNQlvYcJMG5j6aNYae17J9Btedcs+
Ra9MArrvi3HPM8EbjBpYEI6RV9sOk4UDy1B+Cd2vkSvN67sKVRBTROhu8TWRPRumP8taYFl7+dls
TFS7OTOocoOgyIf1jnDTmXkN3hwsN+zrzMRZCk+609pciV+hTm0uS/Ao0fAdBVr8rJi8OQm5XxSq
16jnKLXTY3zsYRFhl6Aj4JZWxKilbadCRpoGNPAnHRzlQ7HHhxyzukmseY2mCnUmuMtV/awVhAuF
EYQdgKHbSORaEsFdu1JBo+fwcFQpfDTHZ09kaFaGpVoBV9UrSrrdHorVCuNXrXHTf3hXPVlHLcas
mYyqeYUccIKnnewPWoMn0trpK3shRNnWIDs5moRXepU7SQqbbLCaYiBAi45V/LMKi0qoRVL/y5FH
1OPD0QoSIKzEM/TA6O5aAvXO8gmX6bMMv9NQkvX3TPTDAVhFIN9OPVRttJ/RTagTgYt+HEhoLRD2
l7mJwfv817G2BecxvDtHs6V4KWOytieO0PndaiCtORh9MypIvElBc48/2JIQ4+pJCIESrQr4lPgp
GSo+nwOmfhOLxMtZAZxHRsy5/vuDD5mpr8pAOgl9LzLP/8KR9Me5j4Cf17qkCbXG2nFDtln8OFbo
a1nRdPsZTiyaDVCi32Wga0vb13I4EihrO9kUcuSiwglKyQ2iaKc8ZwalsdFoS5UGWQWxxoCoph4w
XoS8GgSEgDoBTT0ANzMCv1zGyhQWefIdpgY9gjMCOYEcFdmTOXHAG+7WgT4oIEoTuQpI3lsCtIsn
5DomZdblDAQgtwXtHfyObNfiytDjHNsWjcswcjmLiQS7328uNbf0Bl/f6BagiEkshnCJ9SilOsqh
NhgcuHvKOnJgOSuGlX6peIbVQLPSf1J+F6x+/lxmoz3tBmHYty0pCS5eC3ls8MniyLlZ4WGOv2+l
L7y7rPoYdqaP1A5VwJtHBYHgQV5R91ZA9G9O3XLc/zfKD++30LUSPnCAInHkT8jB+8OoYnxqyRYm
YPLimdj9gKtTUC3tnTeXn5x0h2VtphQ8NukM9Pr7Etkumm9bpJF81waHEYgdtITWG3YcJbFUmCk0
md2iyjujCXLk4tw6w9/pr/cg8fA2Ov2MEphhiRNCNM05V0HS+YUQso6g6E8JcAZN9qaQuNqYSoJX
xtPheFcG1OBy9LUQj/QKYPqZFhmGKCPVQqGdqdA9mM+ivab+RNwdYXOERR9+k4jxAX+NgECfZ2qK
TysnwUgyxwCE3qCaJxfWoGPy4WQwBaQNzQDnV9PUWkG8eicns/HE8ILc0ftwgFgETMGCvNgSRHR+
kk5R+ZEUs3pwQNyzGCdMy20lmcd4bdE7pqjcX97lK8bJ+Dq1fGMWlslXL6UV8W86Cq/i8S7DnqLC
QJeVdDg9e7yHzwGeEX5f6y3CRdJUFd29n5aTkSpD6kVLXtvJf4xQp0BeAbR1lTshAtGiBnBLYahO
OCKPO3PQ6dIp2CHQUzvozg5Ey4GP6IfbMQggoj5HFULFnzNzJTftZUVmhd2dlZpP7ic9az9Y3hF9
txKgvVxxNrt6ICJuzPGi2C4Fn8nki6n/fCkeQTeu2m3u/WBDWcLY3MbzKf/ouh8aDmUcMFj+tSX/
PbS1++VWpm2WWsGEh4tnpOsDcXer2ILTKwdtQKKkCk2U2hlA4kArMlMkO22QK74BV+aW4zk7JK3D
pVv4D4j3jL2EuHO6LgyTQGkdgdX99ma98jP4TQZonDWZchG1TyJRDjJaywfnGBL8YO8CSGug0rnq
hCzVFJaNQPlESIcydU70qyv0cvqHfNeUeKqM5XgeSUMrr3ZUa6snpoH9EmhhjGwrNms8OP031TZZ
Z4sCymG/fUrQ3GiUNStDrcbF56upGXgH/XRgNRBPvpb4gKHCLDOFzdyWf/Q3c2iWVMSpFMxzl6pi
D23ydYBv7pJh4EOqBXIJhhg5yRh4JGVCE3MeL6BELFEGWaXoy3B8v5a8Nburk1IacxFmQVBS/409
zonozMUZcTmjFbT3qKtImryAfAFJFp0lU9jugc+Ift5BewQ0wQt26TSE1iM4UOp8qlW70j5gxzSF
pXndZXS3wZIwSJmirkuS2oFGkN5/NyHyvZVIM6eJ5sqpGOajw5/6L1XfzZcB9L7oXq8BVTrxWZk8
oZtDc8HaiQd+jqnYEAH4ndJqJsIfbTE+TElG4HfcL6/iHXQkjpXRzj18Y5oRyI0bVRYRj857Pn2D
KbHM56J+bOUCk+M2yD9memIJhFflRi1hOfAjMGfaf9UBsscsKmRhjXDSwwvpsm8YDG3o+D8+cmOY
tDWXIPklW8RPvWfoYzb+L3MmotKOrXsYPrMEOFt8tW9qcnMhB52rmzSYVMVDdv12z5Rgcb1AXe2Y
v4XURNkZ2gc56v3hjr3ZFrc9x0uwbXhxQRxCoxZHG97C+F7dLnjcpV2V3PBW37tV+3+bUkwE2V3C
AFbWt9EjJ4Qf2isld8b8X1hYA2Io5SpN1bUiJmrdlm2r4kJH+CQVqj73GzbgvcJ3yfUR0xxFwNsV
bF43Zzk3uQNtD1MoZ+84OaSSr4YKxSUSbXEwBDYY4HmfjjdMKAq3ujK6SISy+djENqF5j8d2sNgh
k9yZgKWyzWcBksgMoNPkD7WY4JDmdRO0ZBN8gw6zjIAx84Rt/2aZs+bn3V4pPS5Tw9gkybFm39YD
pZDw74zGy5N2F6eA1yR0ZxbauIPbTAmMdCuqqfi2Q9r46EaADxzflCGH3e6+Y40nIbabpSLunSMg
B0LOQoeBL3bDhoGKvwrBBIPyzk+59ouKrYP8iZo0PMEhCI9C1ZpnxZ1zNJkGRQef5C5Kb3R7/vsx
459Xv9pK1ZjKmfPPoV1jakPfkJEO4EWmyuUPuTIefZAkZraNASCQAXx4D2pnz9rRz+tZVrgfclde
VVUaw5yoN268+NXzvsLgw8WPi15Ax0NFVRyzHNyD4mNz28tZIfaMEvhYEndV4fIOtGK2puORwHm3
tpD1lSRBVkjyErBX9O6jhI30KlpJWUd3Znzsi+Xzdfkm9RG69T9U4zbi7KXMSe2v8deJ1wxlR9ru
VsIxFRLx1nF5M3HIOAldmSrPwj8bxdY+8e1v82kEMchfrXWRDS1aiAeqvGEjTMAixMCcAsHrPQ97
PXYLMKhqu47UDdEJMXUXTR109dL9eRnVXz5zD6ZUnL50LZ2asFwHMNcUj1hl5b80ShIpKmm3jETP
8LsuQwdh1gTH9ZTs7EXGc0xmSPyqE/MDB6jgIuQry712IdQD+vIpFdbn6JlfeAFm5N7tneSzTZ49
3+IEyU62eTqsCJuDN3BEVAJHQEdfdky+7nAV+nuRQqyFXlPWUEHZb+NF+JSjS8rmwcbbvfiE8bPA
M6Lvafkm6hg6X+q8ySndzr5XTaq6Dey+68510+ENd2mWv0cuCsuj4x5Lkt1yIdy4bI0gLzlaVgQq
bz0SII16QwbS92HhULt66UbjAoXuTHaqlpxoiSxzrjHuHjy39VTmRM+jerPbovyQfNQ8KEVoJVyI
s9vxZ7K1g6HzaMOxjrQqaHZawkgtHGkF94Z04MXNa/3FsRLCnzwVgvnRcDOwgWK6JZaQv0EVCh2T
JlLFg/2lx6AXeBTz7u8Td/BD2s2Fyhr2atd7mp/g/BvN0L3t/uQXfZDoWCSWf44hrcng89HiZ9I8
ecbqe0VryCunUx419msYp+rhlzxzUuRgF6/pMdQwqAFnFmaQNy5m2e4fE+lCxTcKzgaVXIrrmy4K
pB0g0ehqQsaRE2vsYFz2S1OCMpVmbYdnFc2v6e0yJyyGnjOFhwQGgPsCeGFmTQsB6wHMp9NIoJLh
Z/XFuN+doFBX76XghLtykKT9H+woBwaA/7VC/za0TU9VCn2jQzY+4ltRbua8aOTmsaA0oqnWv9PB
ZrUUJczospn3W8+p3qlk+qcupIxBqzjrOanN18kFixa/cNYoR714OvQRmgNR2EG59sgHgXAv8FE4
ecEW70Bv2Soqio/mEhF9hTYNEJkuRazDuGr0iBTyoNefyzeiCBA+mN7HHgr/jJ74e7OTZZGsUnzr
3ss6H80kR/TXy7iQp/9mii6+wIzcn3lP4Jqinak3qzk1An98/ECGQL9QYosMvbNc/FTlnqpM5Czp
ByJeC+/KTMfXGjnMvqx7cgU00RUIca5AwXAsmYD7bFYOwxvRDL+NX8iNccg49q/j6NuIktDLHhWb
xVptUWJnczdlCVX5pScK0TXffLuCcaVUkItpkbLTGktBtS0iJeUXHkHCrdgZbDcWmaZIobT8a4zh
gxKAMYLzjN8+7vVUlSndg91DBluIo2WF2VKpNpUuw9a3fAS/LL/1KhjOWFabXZhYskNIVu5mA7hY
SCHFRAC4oerW5QDPBdifWJjKV68n9TDASekWWxaX5B3IcIsFGtA0B7nud8dkMh0nOcQpqofe1cHT
t5gEhyN0vKXaOJLxaA2w9hrfj7M1dxlXdvXUF07pRRCboKazAdQTbSVIY6nwD6knYPOyqs1HJqKV
/rwaV1xXG7WdgylyE9sKhLgdAwYETlyVF9pjF8hnBK7H7sxKsw+fX49pcg6rabHbFDkXtHfVXKzT
+aE87EzD5qXAGJhtYLcOyMVwYRhQF3+eAJDgmyQbK8OhVQtgPTIkr3ujuURAaKpNoo9WgLhPUPjz
C8tO/ynklk+73Rp4CYjIUF2q+B+8qyb8aLPlnMciBMpeFRziUeohbUArwxYGfPA99uNqXmstVmkm
MCGtspFJm0B6Yaqu3yAb/VdbXwfCb+EyvqKMAE3iFSaeWcKu0OgVEYprSuPpOxhWPoMSa6KAuxIu
rVE1y+wBDP35g2esyS6ArEqSv/Xu4i1MidFnA3/cty/A/9hTeiwHYXEJMzUnjHcVdjcap0VWT2Ef
MxgqHf5Hkr6h86Rwqig1+X62/2i4jnG/YNWuOOZEdfyAXP6Bzvg8riZvRBcaI2gmO7jkznqCKmed
nyH4vnE88X5sCi16i753pG7AaEs8IwS0W6rVxcSEBvu0LHvNVDwLcBoFPBflZ0Hk8Ol6OkvwJksw
+/qxlqozGc2PryVPtxF9vt3b/8v1mfDpOwl3MOJuG38vjAMIKp13jFTZCcSUWlsKKb6XAmEsk96f
TAEFCj+08ET6eswfEu0aXZyS6jju5pUzz4dSwAEUg3XEhL1xfgB71mW4dj1orBKRasKjSpeToIA5
Gdx4CcDPlN2IH42RScfnHoChaHX0j5P7hz35kz30/u/WY/cHge6alJnAvCgAkMatgcNJEYOq2kL1
FKz46yQud79bN+akRSNhPYHW/LMKDTfW/ol4HeO8RVHuUPy1UMefK4IKWSQIzdSVmKwDBZkGnC/a
HvaToj2haBIU4Z9dQK67ONQwoLNVzFROwVuQ81BqTq+NZGjB7LjubijLxjHobAvxyN5Bsa0ZMDNV
5JX+pV9ixGcPfPd9DUiyAcIcc5ayW6GORSA/IxhobVPxDYP8ur6YRQxasdj+5DBqs4vvFfuuOaBI
T6c+ItxGPhtTGPZtmcB+lm7bHB/2TZiymjWMufk5LApfHf5IFlc/F4C7dxJ3ic2onB1H1pP+Isle
0wdTqpvXulELa1jTpOZzsMzFzPsbr5u+i6fGNm1NEyoha4vJOwVn0ZcnZXYyylMjTGRLgALtENUE
sMSVUqxzXGWLDDGyDOvSNjom7FkYC2cS169aP/Cu4blz/s5lD1kUYw2B7aFcxoDNWzvJTBlYm5Hk
SdpVLOpyGnQp7qgZqR5IdoMSpQGS9Fp2oqXewpKf7K6Il9S7j4w1lkyuiny7wCyo81WYhXD57Fs9
Vdq2gedcQRf3+6QP4vZM0FcK+4y/04dpcmVkmlcvre3GfDbYxiQZP8VxpOLEb6K+EgeZ3sHCAHG7
Gu2cPwguxos/KLSorltk9U2ufMHl3V6RVeR02Md1pOsJmYNE0Xcg2jvmA2FSGH6PKEofZHRewxuw
O2hHPTO2xl/3AdNPEw3CJJNhW8F7rzhBcjmJq/omxKfPSJO7/uLr6fJyTWpvEzAwcsBEE3rAu+84
sGXHZ2zWJln1GzMtCL6t5GMe1U5hN9AGQB4TI0qSHMtbmv/yMciWtZU/9SM4SR6lVHEXjFMf/l92
RTxvcPdzTDU6lWm3OSeIGMJcLVAJQ/OSAUv909EhCNOffcb824dNIgsl3zvM2jtbfNtSqO30LnzN
qzrsucKQZsqpYjjZFCHb4kc1Mzxg6Wkw+1wYSinr2H9SBVu1AxTpRHeGWue4nciE1oqDpi9ZUKGL
j+JxxxfAa3nKCmcU4fL7MTA0/4r5E6WAkovuIz5fLGS+S2j3ruHrYegLWboivlzqwNRK9ZJDY85B
ztDtpEuGg5RCKaxK+hOeS20zXpwgkbn+Nf/qJfK36W//vlPXHORj9pW2WCdByFyKWKv8/3hsBbdC
5yqD11DVmRCoJTkjW/qcRTj/YeeanvuOlk/OGlcQfkpgPMjZsILNjK7d1W/2n/84zGDZHadsYifp
sesW55hISsXUqjySWnh7JeBGK+V22V+63GwNlOAdr+wvAwSfUa3u2vRAlzfYeiFK6lr2qMmaejH3
i7yTXUqK2fBJVH+riDpb7iWQEUKMHs3UJU+W0XSJpgI0qEmKpuxPuTbLlGov1pqtaAI6Ma6txjDP
jPcQyEMn8wzV8stDpvPDzCcGcYauc3/yZrGiETn1X5CirdL9TboNl1bZuKTkynktsw0j2vp+U8td
pvAODz30F/JjNBQHUeBxvuHGv42TlzuM3P2CgUXQXAKLW24C30ADWU3os8OkiyDMnjVBN5YTwS57
p0Y/oWApywyXPuMWn9ulrikL4W+Ssm7ccBPruFPkOgDGPpCrPC3TKBrtTHf+7LCpww/mCe/qR1Y3
poMSxTtvGecSgpk5GtI8YHdRItPCQMaLVSMmhPmpzlUN/z2rdXwGjyacM7Gze8a7hkwRqK+VFp3b
QJ7GmjrW3/XF8ZjHyazm2S76fXI+WYGZS0nHgyzEHm2xaa0zU/Cn91EQH/llSfvxTUj+6ixjE77B
qNKKlNJ8xe1Hky5ebDdbXCt5YwTSbcwZ6Iwp1V3kbEds0jsZ3w8UUTWlFUbQyMjqe9hO4/3/DGOK
B7n8SuRnyzAF1smBxaCraufO23FlfJU+shOFj0s74HQg6TKxGHXTKjo13BLQao2nYM6wGadVwu8Z
9NVQA5wqCRkwZNWAbWzKoKC9LS79FCLIg2bj22rSS4XvRfcwLOaFDaHRkpzylRR3115vv0Vi2YOd
0qY61FubJ/ZN2B/bcmOjaoW7veBxVVb95Q+G8Zs62VKpV1vn0XrlN1tearRhh65iLxmXSnxsE5ku
2dn9TbhNBaUJCN9OFirrK+ehENWcVw7lXLM9hCBmVag9HK/PqblK9r5LssnhmrAXPJMLilmz7rpG
9IpPCF2m7vva9iDGmQ53RJlaHAIY6yRpgpzRJ8J2h79er/rdrwpo9YTWqkFiT2JL1ymN3f9wJ9P3
8hBRe1QMci4mKAVoIhq06GwuFiwWP/NryPoYFgx8LXS5CAjAv8Nl1NSaThodmYI42TTuMVLQCsaQ
HfTfFu9mvhFO+yY2TRHo7FQt1ThgWsB0tick3Yg5zdK34NlIwHzNAY3IJrukd2PPo9s/IuqSmruc
zMqebukUOIutZgeskKtKl+Auwsv6cdVAPUks4XORG57ox2zoM/mhssu71jQZvkotc2RRBLO3DI7N
4AWcDnMSCo/4GxVdn4lRtV1a2L5A7UrCivuflr5FNdXy6qMjlVTPN+4RxPXzgO5wLDq+T3Qa2m5g
nCJff2g7kUGiTRfJibgLQI1v3+4v08bsrqTjEyLYjCUiZFL6F4/SZ6mTf41g1DyLRXO+hMVfhRXm
m7SNMO0o6yn4ze6Po3BmA2U9A9plcFnk2upNKeLY51Q+EL/qidEo3sKK44N9YtNoOFjB8Q2/EsmE
3yA9TOaDrDpWmc9NRd6qH6bUmveOMVj03PErk8UMTpx2HQiQg5GtUB9YClAvWP91TR/CiYHgWjm7
sBiBHlTOM7L7Nwavno0fhwRD5JowLigk2MrjkQ64qB/cpmDi3xWY6Zsk6FS7w/WOHAvBftfXgNMU
44qFgdHEZfD/7GkRN+FusSQ/eJu75LY9SJKr4XVuwuDVRZl7ETuk7/969HwFSyyEPgtTD+Y5tWiI
e1Phv02mgVTk1HsxzOkrGDr25aQtZ28stAjaI19JyhsgBAUcc89Pw2eQN7uZx/SDjN+7i66Fs8/k
5K+KU9cRXa99bAc/UEbaXcT+hBVwQCyrQ33sKxlH3OkS2s7uNI6U+BXgKYzTByGN4d2ueEAbkQMf
5BxHvUXzt9oa6DXDEJGKK+sQMQO7hu5/NdAyyPnON5mSFcb81oTpmKdbPehJ5vyCKxhhf6sHe4S/
ErpQkxY0DYMy/BSLIxx7fd2BVcD9ITbwV/njVfZghIz0c6ZsLfStbreVOjEp4DHFuNVrvUSM6ahd
EFvjb2ip22jXIXEn+WHJ5li0rnF6FJB9OF5XvXzxnGCpH2xzFR8JY5tH02tP/afWBMtu8489xgq6
1aM9VtyRfdbxheealdmoaem9/N/bOI1DC52ApQXuF2ugDMOvN007c4MQqKi6KhOfUuWTH2wgFMcV
fXuhuyrYN+Qr7/npZ+cQUNgr6QCBHYDB/7XW8nc+hV9uq1kjAZhzsHU4uVhm41hGF7rsn+LBwwIk
NGkM7kRRuuvqCXOLO+g+ZD+92Nyz1ELgNxLH2s33oxyfVff7ex98/C7iHQp/xy3s8ypV1nw7tFxr
HhjOT4J+uGoTrCeFGdIqWBXstM7N/E7fJ4K9wFMH0TD+ZYu2eBY4kozZ5RobH8xF1/czA8JN/RQn
IdjAgRmFYQWwTo6uRwlZtCfiTK3xVunKMXjPpXnRW8rt4o2AnZgJQP9SMOcimzSLVu21wrUOd2nt
ph65zZchGCfF1yYG7Ih2rxQPPdZ/tCMNpOuV7SUHooAy7zd9iYQceReMnb6e7TtifKE2WlhCHHVO
ovv6A2f/DdzOa1LMEEo1+QYj2o4p+LGvu09pgWtHyXRNJSD+yzNzOzTMQ8AX8czvaA4HWOiTndCm
ZN39hMRI2ObuIXngJo0lHiylMpMlVFEPV/vUe9gOsbyGQqtW5eyw8QvnJRStkMAtSIf7fKZGFW6x
NtBtOgRGOgKJNM+nPWGGU+s+3Ef51g58w9WKOU9VDH38VEM8vW/zDyTSrJxvfhg+lAytpj7sButx
6ysB0pVs4aoC5gYjjbWYufy16EJJEecuLMIbBl+ASUZFqv5TwMKFfkvJ9UcHlP2PBQwF6XvojaHe
GLZoO7sS8X42flMSuLUKqwKBwpe49tb38je4MM4WTseI8Fr4nhkpXdyZbVWHK0/gFpTLGqVNla62
QdpYj+GOFTOZgq0vV/75JguPHjhDrp472RRmiuvbnGFEJWwqrB6RI/jaoSmk4rWwsqfGhpkZTKbM
rEEOC40KJ7L7a4vllBatlS2XEwvgMrGckyFGTbc2S5GbOrbXYdnlt7XG+AxXM/XdsRXe+QpaU+jz
MmEG1CXMOC4nykpXp34LX4JPuFgfgtKLAPcj2HyEVKi8LvyDwMAfkfd6UY0qMynzM501Kqt4JfQJ
Vx+fYxeQJB7hKnqoyext+xrFg4KSBwAQNnwjHwJcaWafvAQgTTsxPnMzkwmsAitWqyWlRLEKKLPl
fLPt0NV7LlZvvSzNlNB1MKzd47DVHbvIR3Pc06+QujYEmiUJguJzCk6+Ydg/l+guW+8G3MQg58ZU
ho8jYXfUDiJS7HRCxs1O0U8E0iHNJ+2zPI8oBKlwzqudDVVBIgdN4cBoG6uc2NVrrGYgpm0VOA+n
gZS83gQPxX52bnLx6nSbyM7fermVm3A74dqVhhnKlUrKLVodvaG4a5+iT+c7BJvO1u8IQoH9Uzro
S/GkQhdQPDsY8fZo/OLtJuK/EQWLDGkJPv7U6Rm+wuo6bRN3mqU20e1rV5fYXMdXlORY+NxDzJFp
m2bV0i2fchq/EcbKuzkHWCHSGwKUXUPAqrHebOhTTDBB2sGMWuxro4VcDQYzENTb/WKSlWNhCVjS
V2lrRuncIuKw+QLeG3Kwq19HamBS/FXt6jm8Y40rLQ5wuJyqWrJyzmcJW5rXk3r3Quuia/uHKPS+
uNDAKorwNZ+SeRZAmTaUlip+MKgV+7ECox9E4ePzCZsE+zdhP7tUVzHy4Gj6FmroQ6L0nxztj7lH
QQqrP92gINoY6Mk8xKnLrwQ19hOL9rZ45ms7iBV+p4hHK5GcSYdIwhBp0Pc0o8sSE5/uCd9XzeFl
It2x8NCizgLm2B6tC1Gkzw==
`protect end_protected
