
module ds3231_inikey (
	probe,
	source_clk,
	source,
	source_ena);	

	input	[0:0]	probe;
	input		source_clk;
	output	[0:0]	source;
	input		source_ena;
endmodule
