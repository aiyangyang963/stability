
module Qsys_system (
	clk_clk,
	pio_key_export,
	pio_led0_export,
	reset_reset_n);	

	input		clk_clk;
	input		pio_key_export;
	output		pio_led0_export;
	input		reset_reset_n;
endmodule
