-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QQMw8v8hVGZYDk0/YjHI0dekfmVblDXNyAtVkzc0Vt/dzzav4xd7dvi737Fh0K2w0rZ5OSyF873s
s6zIT/m7jQG0LiIa3LXeL2CswafqqjGtXOb6nSrR7DuDEdJUEPcdkAUdHT1CtSDB/Mg3rrBoIQ+i
LDwMHK6UkAmIAFSEbBGj1sxSv85/JUroaAbOZFOBuvE464v9roU7ZX80K74y4Lt+l2AQtEUopKjc
FdjSzxIbfQ5kpz6qjdIqvfw79N1lxN1s8lBjPB6Ri8RHqtANRPzpDLnb42t9VvGKyor49ramZL/s
Lza0JLQS442+/g0QmZP6UsMpFMpsV8QOxT2FzA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
7IKGnBVkc7wf7K4Sul/Q+AcxF2AMLAhcH+xiDXau61ewH82Hs7hX48kWAEOIlEHG/cmv7Ycz4jmu
a/K1bcJzcP1hQabFzYy/uvVtLGFkZbf/MSH17LpeGCAkgPNDXBgAQZnudMHiC/hQKMpzYPB44Vyh
CBAjHrarVfFrqBp932/RZAhDnyhC65r1jGqwApkgvqMfbF4b6NCjG+ee5fUxCGBH0Zj8ixDuTiiw
qcHtIzeUq49sF+zEFdd2XjniBGanKewyEoAAeUI8DWHTAxbwMxsSECP/wOvWA/PATWK6ISDsctm0
hwzsyP09p55eQs7AEpFDDwOpKhS0t6IO0bz8o0EKzDwnk8i8cKKBimxYYFA/85PDLJi0R6Q1SrDq
HmnnukYkmpCFDpxpyHizxChsa+I0fwHRUP2x21i+FULD9Z75PVIAJRh9s098OZdRx4XkaQa2V36W
JsaRM74QAUR25suunoGwuES4jjCuudiNad6yNl4tzKAnD+xOT9mdv5qKAEx8p++d+92Rw2gV0rrF
K9l86RB0GNI264Er/BTI9jFroxKr9oA/sMXZSwA7K0uzhzOo6i0h8OaBtNgy9Pzxjr+G4NWZHyUP
ws/o8SdwAYMQlLAIL3GNygURIzJEECEe1XtXbVBK0IXhqHn2d/n7tACzmymIvmFctAeveeSIU43z
+/nYCnt9dQVVxgRtT1HlEoxynaPoZl4bmlRrSMz3VTpycY8OIa4kK5eb7QtSWnYC9jJMnwTk60y2
/ot0EECMv2ePXeBxi2Lnd+38h51wjowsjd18c928tWstjPsQSDDdMi2C0+xxGmgXah69DGx5b4q0
A7JusgBnganL+iiYOeEvHkAWduFDI5MCtTzEPyoAJJzU8d9KbF3LUUQIIaxQnDnieN1lNzq5KKO9
d+te8mCbb4yQTtowW40gjFtfSQG2L5iOxloS2f6BmKC2p3sFbAm5zyUEBi3z6PIzZ+TaCSVjTuXk
sbt0PHwnQqChDIfsaXnN1G7iEKCt/8oX2aWbS6BrnUzkGsaz9b2XdKaWuIXT9IEcPWfWr3u89H9I
X1cHiuCFewrEAiw3cgtwi/qJACmYFJXYy0Tp5B6fO+2SuChv/MZlBvSCKxjoLi6TXjZc2ogk+K79
7Yo5lFjziiTxciK9MAs3qksiHou5i6OlHkPqocL2ie1cY/lUBY1klzQVsyzYcrk3j1a9jzKzq2hA
iuj0S7Mj/GSRXLLuZYqHr/Jk+sbCEZuo3QplQVBZvxMVU9T3JIPBCTlNv497v4HaYs0CLx7pQigk
8xH5aEFmMN5tFkKjAfpw2Epdbls+e5Q6Z4BESNd0Dleb2w9waA9apWLma/UP1ZtVu8nWE9KRCdIA
Zhb+L520hmJ0KCUuazzy0IsamgD4u4IcSomMe7du7HioIqCTuNRnrZwbJe1DMnhmnBYTv1wNC7xS
DUH/GdeDY52KbxGM0bPCF4p2Kk6v2Ec0mjFF75z3Cx14SJ04gDlOqsMoa4vfzs1spovhV52KvtPO
yZ4/JbzBQ4/jjFHUthJco9K6h3LU7rx67cLTx0E+xdeeloIaYe679aOj1xVIYdQNpPWDETpnXtHk
pVqxkOQn2r07ntD/B04Ur5YzfQ02XDYYL2bChFdAYrDEp8TMfmphEvk6Wk3+aUk1KMKovQa2Mq2H
9ds5om0d9Eylf2mSb+8AMtqpXGWNIMd8w7Jkq2KD0dSSOA0aNXyRK5SMp92fqBk0u5OZAY+SW61r
t5fFYfILAnTPUIUwgeLDn0VNEVlMAxFUryiqot00jNVOv2oId+jrQpMIdoAv760iOslPE75r3/7P
myYvz0brIXRsVQbWRs7yD4jgr6q3MURVenAZYWXn4b/9MZIVgP/VhhEmnTF+HFAjHhgz9+Fk9s7P
GZrykd76LWv4LCxl54KRmiQddQGErvOVULaA0or2l/WJYI24taTkvePbyDyGmO1wJaKe7cP8BcYc
n+VLhCjmvADhbgd4MyUfj+7sSWqmiqelcxnw2todu46QHGVYUzVid+IGLKlNLrxCctlS2LJdNU1X
ptgU5qpTMP/azeTkumUQLs9j6N22HiYoH9cIcfsIEWgOYjbtHSGGBhMJWt8VTbziVE3UNbFDc9+a
ioZgZh8hxBZMw6a+fmtRaRDLFxuYn5sZsP3Lsk5wDkbvMSgVgEXpUnKXM9o+9m7cYTFCnDpMaiLg
j98vWRaXvIQmCD4auWE/O1JLj3RTaD5SCLSi6g/pA5gtrSXlsZ4JnTNSNLBRfWFCv4CZlxC08yDr
/q07Fv5hRphj3qk44KGxkF94OOHLLGVSeirAxw7BramRy8elbnJgdIsw/MPD2tvwDOqwr3N6jRPK
H/WJyl3JaOnmG0KId/cqcySLWOwQqBZN/sJsV1yeWRlFMSjtYKJhContwT8CQKTNCWiEHP8URf1L
CDVAcYRsw+87HXpF07IdU1SASO5tRHeTsJU20T+RXVnUlrmspWI6s3OCMeFB+U5UCic9hGMWJ0si
6U0IvEEMu54hBMgzJv7QvDRwyYFIBFtHikdFWNBUE8d4zjE806X+geQdVCFWj3lozm6Ve3hXgGYI
Uf4OS2KAh5cAsU9oTrBzakKIMaC197k+T130qYgjreHMncoKKtxyvIrFnDVUhA17tQT7Myvups+W
dpf54dizj/ROImkoa+XUV0zN0ux11QjMGf+j1rqbS0uCvKr4/6pr7/iDTIWR3U0W0CBZxP8UWBCz
GflkgTJGfhMDsLc7LZ+G0CsOcrnIvbTz3JUasBYQRM0z7RCn6f8KfFjrzF7alWNR7YzzqiuxRRfe
tkmYS5LjrCyG8naDJMH06j7vyp/8GOrT31wgw/Otl+sIN7QAro4cUi4+4mWSu5mkYnVnnL6tVZ1B
zmT9buNC238bz1iyzRXxlRVX7l+jaH/CESHPIQh1u8/16J1Zt1ud37mgoLJVDgNtdYDZcj5xXV3W
IMzg/hcTK1ZycYEfH/0+4pNubaHvwSQztu7C5SoH5UQiRJA7bn6VJfcVRFRLYPDd26d+UkuBlZcw
bV5e5NE5LWLylIl4TNZtzAWDpv3Wr6C7GLAVGasF5jilZDIa4wqHN8O3Aj2yoVKICRcoyBv4WQsN
qm+RiBTCGmQ5ogZ+vAuNTo9gSj253PZkPZ3BJFTQrOCoGFP01aDN1YeDU8c+ExOK+j7Q/8lY01RR
UF3Y+VbW4/MXvlhzF5M1SCJsFtguAkfLnbgr31rWTAs/R4yXB0TpqSQQ8z+Cd1M91SHw6AD8m+nf
sal6Zlds4K1f2+Wnw+4ryUWo9+F0jFtTeh0VTmMHQmzvCJTX+w1q07USZpEQpgDth/MsS7DK4EAO
gSQJvIPHF2G/Sbue9tu9gqI42fsPjZv5gDojSWRVUlJZr2nGrIpJoqt90nH6HwDhuU4UE6SyUO+F
jSczz/pgh4fA8vVKJSpjpE0akxiFdR0kqje2G449R1CCiAOIAH1tP+EKhGgcAQfSLJcExXJXiOLX
uPgOwpQyz+2bJBeSpsuTD+Tspc/7iY4tI4EvJafu9IP/qS7KFN9aiwiw5H0XES3ZPVN5ioTM+0J4
eupcp2iKlfveBOxIF2XP3+U+SkapwH2NXgZ6r2nbZnV9QmMhh/nTdKKEb5A17I+zVotOVLGsGVT5
Wkjcwy6eLHwRFi9oZGJPpTWi9HUsvQQdROSFnQ+IGLz5Q6Lo2bY0l+Gj/B8RMrFRONrHEjqaOtvk
2KJUsxykuVIDydfmIfblhOinX0r9ljggHnhyYFN1gGFdn7jIFR3c373OdF7lMp9U+ZIEYS02D8Gx
iK50Ob0Um3WGmoo3biyE9b15ukuwcYnptPkXjjrbcI82cIqBmMwc+UwI8g2TzxFpEKdgnrOs8B+M
V6OvM5sSsgZ9fESTe+rqtRlBG89ieGu5nRAaTclO5fuUMHbG7Z/T3SND9B0jbbvxMqoHcmOX+IhT
bZFUj2taNRBqYaCFVyuGRn0nR5mdCFYSECnw0eAJVDWIR5wxLiP8pAOBqN4gxFoxwr7rT2xSmbmW
2pV1owXdLat8dyv0U3mQBVkxLMcMHIEWHzFM29yloio4oeA6ohK3a3TJtnJKyJCE73xLyBHGQpLx
K6Gdct0V0VSRWpZrJch0BP1+rbaWOXopK6LwOmszm4gmFlLEmcpUALtf7koOb13YBjTWlkEzUnEV
s3disli6V7Vps4RvB/apkd+or1t5kD55MxxzWKZ9QJCHr3Y1zsN0QqQkFbT7uqMBCgtA3wEoIVH+
AX2+Rwjgm+PVMIr/7aMpPuioU+l3K6AugmtYaFPomL8sLGx/xkjjQa6eyDIIgOMm6G1IvJIXB1Ac
G50sphdPigQCM4RNF9BichgNlqgYeiQESEd+4LuZwLOPYwOKT0JbZenO6c6wu9PstEKelKpWNXqv
AXAx67ARTjz6grKSTy0LbP8YsP1WfcAcMCWXejO0YuNST0owDf3xYrkQUi15e0Bqdow0xpI/tUBz
eAZPNWZmP8kI2A8C4Ewlseat/rmoMdFJE4xC5LhT8FG8p6DFrU3wTjIjt1m9zki/lHacd2DCsNMc
DuAEzytMxRXRTKrfqVeBlya1Q87fNbeyfnyeCRc08lRGU1X6fatsHJ9n/c6JlV/2HwJoh7yn8GaZ
TDXcIrGl5OTLE4orqN5Ko5fSZ12QSCUgd7Oh3TP7n2FzaaI6Tv6mRdNJQjn5trrBT7EgG0OBx41s
i5qaekydEB1SSB4HNMoubiz1ENfgjkHXGkcUcf1lpmxfTHdDcSWw1MyinAG6tmD1Z3dNgzLnQS0C
T1keDslXavkqZ/WiWqpT5ulE8Yur6upIL1Jm97dpnpRe9o1ERBSVLfVCRRwyKH1kpVyVOJRldpWm
J3hk8MgMs5VToPF2dNSDXhaMlzxRIPIyYu3cGUQCa2AlyJIXGZ3jealwDrYMUtBqzFibdNmyWZU5
y7MnLXx7fwidtQHbj7iUC14VK82VIlQoXG0GQIUoCUzK5xeizNtV8QSEdwVWC7sDDqGa74WmR8KB
5sxJg2xwrNrUhkNgS2SYPpCnYaY9hP63npiqGdIZClGt41ilK6xVVX0UTllMQ/5v6GUmewVfXyLq
D8cR51HxYjiCXo0eujQaVfIJD1KwKQQPBZhidrUtsv+J45qgjc2r9s10zAzvjMh29XgXR0ZIxd7k
JqtMlxR5KfXWQ1DQYazrCZDudA2eK2sx0RVyRDfPISd+WCJ2iPjB4n1rWyV6dRlA7lFgbcSSrQn9
jBFFSQV4fU+Fi0yBH9jc0nXuOYoS2cRrxs/f5yxIUN+rQcqud4J3wZqOP+BZ2pkrZaJ7P95Q0Mz0
HhAv6GOIugeSwbicxxZEmJ1IrSo20EBmEKjN+bEjyAmvwUN9SZSahPR24rlogDU6TLzrGzQ/LJ8S
aFos7S5ELCReYUu0V9Mh7u4BQYwaiWj9uK1LE353BQ0h0hmtbSXEzELREwJra/5xBuyZ9cA167R4
OQtxoEC7uzE/lZBsf+gCdmE1F6D6CXlS5wNeotMhZg+gJSjbdtPqkdrKmv7e91G+sejwKXuKfVs5
f1u+thQJO+ahnSOidLWcKQDyhFnrxK/MtgS/YENF7EdXWvE3AkTnsdXU/9PO50QoaUKVBhsjQmb2
Q8xinaNkg8y+o1qdI172NC0PY6sYd+PyRxxSy2abm3uXM/Dw2T4hgxUnF2O/W5Lu3RdX+voeu+Ix
QYrT6O09oNPYxtM/itGtC+fgjGJMVOIGm/YrqwfoHbzMoZCd3chlhpD5rRcz4AEEcWeYP322RbBq
KzZQscNVJJyvrwgbdTaKLyB04GoYiuevRO1Z+RiKZ45TanIsMBRQRzIOKdPMGi/oy2CvPByWvCKw
DuQYCIzWraRVRebXOLRRlV7FiVh4npBlpdQlIxdV0u6lF0PKx3TJclUwjwmuhsXfDOXdckZlM3FM
qYt3KPd/C2OztIqrOlVj+F7+yFn4UtRZPbslpHjYiY/cgFr9EBG3O7GupdwSpKmW3rlylmW0ZDrO
drG6u1USChqKjucefVxUj//GVOI3O5/VDd9rP0Yuq0tkZyqDYahNQLs4vzFqVvuZOXcyLh/UHVWt
RG0X6Qo5bqoC189c5ECqDznqfUzVw6+Z0M34gWDy3ydefl/TQViAooAa0R4BVJt7q0rC+ypbt0+9
+LCEOYEFUrrswoAfqI0m3xyrAUh3K/KhWMvdj7+8Faoyz4XwUtxCNz5jLK0fxj+GpwKOx9BUrdhG
rvdagJA5IWFLHJBoQoNLhtqwIARg/l5z2MijlT0sR3i6C4oholgxtBt280Zmf0N5CrPtQpS9QyEk
OERcHMRpTcJe+tn0RYLjsuahcfZJmcKx7eecTI7vVk/nxqKjNyL1DICRTPDQr9Wo0u5h7QADB79N
ePS9ijSWbKCc6+OjvPE0dHNv0sICxmeoGK+C2E5pPmz+rbH0n+9l4dOJMxWRwZssGZ/VCgJZymZr
Lqc9VnRKVw/ymUyWL7DeFPJB27qqFViZi4GJb6lzjVNuvblgb3Itlym/vGKMkN4JkOGgTNhc77Qo
IFUr+BK5veyYi59rm/R4CfUFQqgPxZiBJIGF/CgkFkSYmRYye7ZfXUmreJTeFpJOt+nkxap/eEda
uJAyHs5OQ+S9KpfP+7SOsXEMHg2hcNsUX550Mn2cbMzxrPFzK1qqW/VGAgdFizp+vppeLo2cYGA+
XaW+bxTaRCsagMYLyPddJeNfJePuSLzsBfErWP7+sceBJq9d0C7YQE9TcETf5kmeykhnB2UadO0M
pB2eM3ltbX32+7vEq9W6YNtQf5AZUGEBNCf+bsPvYnZxVJWrj8ZW+xC4LjVDNONuye6FqNJQdkA8
uHIdYwq4pk97EVsYcRTLWxFyMUZhxIqch3UOWX2Lm0bx4tG49J1GjvIbDOd4QBEWio6jF/H2eJHs
APW7OgQSHl5IAsEWLRxv0U+K5uRBxkul74k4BapJkopIgU5P51zU68jyzkwZCbWzpBnMXeiOPlFY
trtWg02oiNww96Y+f4SacY2OeRMoTN98YbIY+ESLTdthSC+AS7C4baFBYXDddATfGk9W5A20yf+K
yD0F1jwCcoyZAnzpiU+b8h/Kt7un7EJTfsEdnjNy6bQUQhS2NarFT/gO7SHXTW+BTdEB/9fbZSUE
zIXmK1+MPQRl1wuDbtf0h7kw/U53QyiuNjaOHJnWm6wld+0zzKMc1zUm8Ily5u1dUpGh3iS5EPX0
Kzw9t7R1XtTy74SlHvbp0Apa5pLhkDI9YEUvv4zqHlYbYiOK8PPCqE+Zo5+I7k0efeFocRiFEsKp
g0mhZuWQ2noiWCpD9qqJY8OzbDu8yy8nrcpLWZEHFYABWmNeeg5DHFT+h2OtfV4HzJYryDK6qbMo
fSx4F+KUXe+YO9boiGPAls755/Fnkp8qGh5uNDk33XWB5+aM7Q3j2NkF72QLyo7XhQEkdUmj8xtg
G9+Q395pqo8WPQMe03RHptEY7hQfmIbSmxvf35teknP0NPlbiBId+tUvezNZXFj2HSP5da00Fnx8
9q2e9xp4Oy7/aq50QryaCu3JSIJjObfo3ruCGl1KrRSM1G1LBgmHYMCNZ7Myky+VxW0+YPpsAgmR
2TyjYg0Tc1Dh9L8yA9krxm92LZDV89jVBzn4p2XjupqtDIEv2BY7jjqixQWWIZrfLMifY6MIi8wa
I/ulNuIqHX1XkpzlUErnfeJyT/qkdolV9ozCboXxBJN06XQi3DEKjj9iquDhp8Pc2dFXnaJD+noS
kp4q/2I9qG2uoRJh3CRTT1db7XMrjaX2yad4DGOIZLheCz65p51Z4/fkiL9BwQWHpZ0ZYMx/o3mt
pu3W8EKgeHkeYbUBwDzzUHTUSm4ZlBPqOYRfbQTxA4YlMBiKPkCaDOlEkd/43moYU+Avywo3g0Zz
5a81nuS7IpROJttos7WQm/OCYi4YGyMhRjuccoH9IkT84l3b/+KlO4gxofvP92yK6dIp22hz/7pW
8S9LLN2Z0+vqyDRsU6tuBDucwy6KwNbGE2klnPEWbjrMYTzRb/a12XmF1glxY+wS25D4JqLx8O64
xbDN1nRtl8ZDdqSh1X/ZGr8ZGXMcFTLyc/xzpIVTpmkFRaXJPicAf5/oEF5k1DwIIr1UrpcMCMLU
MloDin5lPDFwhnarzpb9rPJ2n/rfh91cNREKuqfZ+PqjQoZNpA19oLfmvxokAY2AYcwE7mTnv0Oi
DOKaiIjwRVJcPvdpV0kJ7/EWmuxUpNBITRHqpT6xIN8Z6kIxsiCP4zpyBjnGSvN7VB8rAH2RXQwy
+80AJ1dz4K0i8FKPrejntcoqsCz9XUqH7LlDmQOAX7s4zq2u1EWJNvcjfOk5sLZWcf3UTaWAy3vf
wwnw2Gu/Iys7J4uHSlBzXGzEBBWPmPbx5RKgvCzDFKPO0zuvCsqJCpMNQB+ufj26cls7fnskwXdk
1smYrwUJNW2mqpK20dsxL+HrlhemHi9fmoB8KP/1mIGquZ8Q8kAx6hJ45b+PHZPbZmqF17UfMltS
DljHMg7+sGrf1wAVZd0g0N5g02OSsqONBu3D2WeVlS48TXHmm3bPAx6Ee4a8Gnd52ycC4rRZ3peC
EPA7FCVp17W5lx5dMCKBkqV7xbIGUflGvlOkSiTosE49GifHtVdmsVFkuXaVe3B/MXxtnk9kpOFp
0bl0vxqxVD1IFiW640zShm/pnG2wclXSKAjDcETkhr9SWb4m4DVj/3oVtipuLnI68/dYd8O/HWUE
tgD5dyfe/gfdi0KUI4SpPlsqM20mVGkxASEClm6yuwckNVezUV0oqlS3G3Yx3J94hsQvoOebaEWz
9Ul8XRJ9FQKqnV0Zf+jX5Ltg6oN4wjrnZT3nyFjLCPpBc0d3/qOEba0PJRKqMBHtecmr5MDHBG7o
wO8eHv7YjESIWjRfLnwXFC1sY+UmYlpqggVyyfXiN7rqdueajSnA+iVAnTJw/2aRGEttIAdCslLl
BvRZwNeMbllJ4YdxcmSnxoBGH+xGHiI9aOMGz52NfLKrI0xJTOzRyXFsdYj97zON4/ykfJVUGITu
ZeI7uYf+lJVfOtIMFLolmlplqudskU36UUED3vwyPMKzOAJ7hjpXv2UfexxUHuw4pz+lF+T3BZ5a
grz9Fw8oZcCtM9mQtn5XI/eLeNBpqetSiFJ834C3nnJQH13HsUua9eQrYIuLj6V7OtnsjjL52BnB
T3OMtx6HPte7nd8Jw73SxNHK+tevzFZ2ygLkwIWXuxskjrNLjtloyhZ5LinodEvLCi1Qv49Am+jA
sYGGsOVArBdcSpfn6M0kprSEHo0b+ZInRxhoNTlOt2Cm18/Ac6O657MMpgmaKH2mazFTx02dYg8l
QBpUzS9QY2IxPtXI5L8w/x9wb5weOQkqZVQc26KU4R0X5rsbbLSJGD/7uCQ9zJZjFaI6Lav8/N99
j1qsx4mJjGf1HugWKII9OVtQ4z356SXzYnLlJMYUue3WApQ0LS5ypNKyMbAW6fKl77CxPnm2bkT/
k6BKf7gpFa4iushoHufepXQiW6on2MQ5TtHxcQlPuW7/0M9P2oTmPqA6+HTe+Uyw4aec4ZauYRdA
Cerh3S41v9P8ao2H2irZENOSF6lgx1pI0FVpE4OWOTJaqqDIy7OvYP08qf0/R+a4KhXhuF+ZjrQO
YBIcKm0qiVL1XNmsmljoMMZKrvh2NI0yiD8jrgy+b6DFgwD02NHWcRtqnY3LRN+1gRGgnDiDvml5
zVTb7/oDYZoJI9lrm069wmz4Bfy0extIsWoMWGQIbFcjsdT5SoGTFfuc3/kwP6d8WvK8d0qTRCFq
jhyD1pmk+mPsttP7TsC8i0fuIerAsQvlqiUZMpK8iLbCY7OuNZumN0hMTQqsnrM9uzTqSoyQYjun
gV3qO8my+0oyryH2v1S6iSjPmts7YnAbtuYsq/5jxMpcurCZbGnSVlxBvWz9AIWHI7pWEyjnX8d1
oUU64/cPiYWJE2gbIc79KMBglrjAEfXwoOtWcSDOr+dH7DrQmA9BV/6tMGIgXk7p7PmrBbHjf/s4
DLlV7OZ2xONuF/ciih5EUuuxFIjPJankI9bpnbfSW129GqCehQkbJUYJ6UDCYQRS7PxFJ3Bu3RUs
Cv4sgeQb88gciahHbqe0+9GTbfSGf0pfPUE+NRLai2Usjo3zGy7Lu8ww0fA83UzTwgpEchAqzQwd
AX2n0u8oj0C9n7G1FOwFUXL/15lrJzih1yQw2DMwAKhnInHEJ+BcTCz+nzxFfyWOdvkgSjtxxTCq
PErk1OtIbjMcdgI3e4Bem3WoQLJ1VvBFvDvKs7JBhHi4xYcRH8oDQUmO9E+pHAGDHZx4WTb+5mnm
XCaXInb1qvlQtaCeliV4xLgceLQtabxiWWWjcgg2D2h4tKtwWo5zOBJBQvFgYA8LnjQLrBefP/Kg
IGmjR3/vQu64Wxqt6cfzbu2kB6rlYtixNIN6pD1/SeQ17GXuz2J1MLyj3/2bWPLHeMri3OYHWfZ2
e3MlcfWS+g9CQyq1sVBu9swH4DL01qf6lEHSTetBiQCWVt4gjMYAmf/nKzZN4mdOFSISRKDAKctW
r4yf9Z53xzBUUCf47LL0alrqph4Or59uLr1Y7d7u3s9IymPc7MhBDzKCm+GAwbRPbrpIkbGSOwSM
vqC/jI8p0v0YLJp5HpOgVf8jeMMJnu9puogEyIDwaw2nz368hmCTnfXIF0K8FsTGCNyz71aU6rLw
atzo7MJgDe9YxtHFgXjdzLuR5VMpoOv70QRWwft43Srtxx5up72Hm8ePGiNKjj8UofuJDx28gHZg
JQqU9fBzJuwwkUhDc0PmJa8etV6ybdRexyDhTi+Yw6Ia91FAGdQMQzlxQcB3fi5/1MqX3k55O+qx
CfhnQa6czOA/hs4trzvArj9gGc6TxycxMrxf9nAiwVmx47Qz/WzKJ1xpzeGf1/zOWSqOpGU8YC4l
riaD7SdBizvEhQYqNqrxbFHxmU/3OusO2nQKNAcMYcXvmQPhff1Tn9vzs2GiAZniZo7r0vCXQC4V
4hIdyvHCsJnWXc4nkJakJrwEInOrYURXb126pqy5slARyjo70t6o4SyC7nlN4O6RMsqlbficOsvz
d8mt9Lt+bdtT5v09xiEDfyXuzZVsWuk9g7Yto8P/FSPQRSunsXCl6w1G6WGthoox/ZV27bbprC6A
x484Fbf4SE7hF8llzURm6kg/uGiBgY++lEW0S//YaAzQkEuEuADQIfJzis51E0OnCuUz388vH7mA
uH2eT0d4N+/aTn52i6pGvJmMrKjWHi4ngGQbDpCrsgJIL9o/cuH9/GeyeZ9Mt/7VtRq3jLKIx8tw
QdVz0a2bmSpHdGDtbrK0F0pC4XBr79N1w3UHZfwBrQeWpq+35jqIW8V6ENPusA28B7nSk0l27+Ah
mtjczGyLmn/twhFufakvpbrQpbYK1pnpT33bJK4I2A7Xja3PS4XejcDYbWEUivva2avlqSl8y1Hp
FmGvUbR39+PhDO8TP0wBZG4BmaTABdsUAgs9/TAvfpXYQbwFvJZgbtvZ1nZG8P90YqhZHjKTZzW7
dkktac7urngnbsmU/o7CVlVoqs+Pu8sK0iXr6HzAdpJG5PCPmIpPij8mku2NC9ZCCkoq37trjGqs
ttHTh7Fwf0WDeRV7t9RmJ/sTy1JlKsa7pyXSZonShkmGPNfJttypFhNLap60F3U2DrLkVNzkz9Bu
EzIBFYJ/r7OcW1ZV1yT9p2/0sjRxc4bI/3VYEBcr6Pt98nNqaTUU7lBZdNn+Zoe1jTUMG/USV03t
RKnzVhueWTmVvdI9D+SYQ21n66Ff8cyTwCUgIOWPkWYuCpX5hgmDaURdTJWJwwKUfeg4RGoc9JTY
T8/YekGC1GMIVLOY3WQL/Rmis0I72h2msq5pKx0TbliOA3zHSw3eKHsg5cDu/ssdmvzl9ITu+Ckc
S0CVS98hwrP+jhT63ZS6bF1vvn/45CZO0ddE2vKKYwu240pGhQNwyTNULr2485Zign2upseqFkf1
O3PzMC9egHLyqjHm3dTjhmLZGTVrY7O31MzlBX2tVI9oITp2pD768PFAt1+Jc8xLcMolEDh3SNrx
X6F74U8nG78MmqWEqpFtXYaVFSfEjIbPpUFc75TeBuecORT6+3FNz6St4XBONenN0S9KDlYzeyus
gAUJVkWV6glZVE/9KpI5R69c6S68I0FJ9IREUPP5WAFSelTYCQWXJpNJJZI1XGy0HjOkisxdklU1
Hkkw35ZKW8oPP254aJvZJiiD8NWQSWTYTUbFXRh06Lz5V7jV7cGs4/qeyOVMgwo2vi/cH05oarvA
PugfPppHOYkzQxWCN/HYzBE0dfT3ZvwCU2VclvScBV1Wt8F0t6IbuoqbReok5NaCBH1WmcA+VD4+
mC9KhZAGm8ucthN1CsMQW5aK/DfAacEMFnIyVvwDeUVgwN1zPh1amjzK3FZ/axx0hiUbzlf3ha06
6VsylB8UIJEXSJL/0fpK5Jma6MpYAOJPkeyPgS+38sSlADt0AmhxEqF96KBcCEuac+Av9FgpslBH
6TUXqJ/bbcKMXOuJpeWOXsZpNk4UT7TxwDGwfr30Z+E1PULyIkoAgfUKaCblu6ti9QrtP4vHXT+x
5skaJz+JhAylmCNBetbDSSxNl0lPGAmYL5xXEj/jaqd9gz7ModKNgCdLX6FY5UWvro9RVehhxlDB
qquddVGw0+SIt84Y+4XWGsl/asfQF5B2pwrFAKZw86qHKreMCSNeuuACRCE5WPNdd9SG506HeF+y
8JmtFM3ueOyPwZZuN7fno59y/Ltn4OG1Yjhd/zsnyvOmnuZc9xFaAR+KmdjV7H2rvfD/XinI5PEl
eJZXdKxiRiqS3b8CvzQdLiHBtgLvBNbZiq7pb3ece+hx+L5aJpwnRM+L+bXWQCzTUQRWLdVT7ovL
zg5ZePO0KIfxH9h5cTX13EIEtHlHPkP1LZRVDX9aR19WYdV5zo4ksZbEhpwC3YHQACNQuG9JESxe
/LbrhOuyVluplhEzy1tI+qfiRs1qxkdW5/go31itPaBYpeFyz/kiWzAglpa1CY2GK14+F6tXN3li
S2yCsiQFDo7KFhdQOg3N5XMV8GkxPOrgrrWFHWZT7SML1CE4BHb7kc5Pd16SRXsTy9VlIX39JCM+
yHStxDZdj+23rkXtWVk4s1rzs8JoB7axJ521yvT3zd3VpRDOugRMkE/eCGXZsHvhZExcdQuOgRDp
irKBZv+NbJ/tip/0q8x/K9tMsrE1plwyplV8ZKioY02FPiupUzvbgWIvlRbiRPeSCRvFiEXgbPSe
VDYtntju66Mer3HPj8HT5oiJeDDIqBHp0PdfVUMjmvXSwn8vl3EsREYFYBnx3HR+zzu6Gblon9uZ
VDGnZ6eARSU3/wKk7NHoMwavV/4oYd7yjySkg/5dat/McPJoy9nAQoKlChXiCRrvZlvQa3tdDYZf
DYGo+vzF6l+MYd5Dik+A9ItfGlkSw+Q5kUQSKVKOHvg6J5JNZ9vUgA51ZVPrXpO2PU+hiHmS9grH
TqXuwen/DZ+WpmuGDqPq5GZoDOBeQxPBRa/DRMews0SgOTRMbSTxYzDgPves6RsNbJ1WEPVkMQ68
Z4iuktiPsUmHSnutHZLnIiwhStbCPsuFIN5bGQfdm1Lxu7XA1USgNG31XwWdur5V2NeR5xVQgr/p
y4qSboSh/eUb/a0j7t746KMGQrji5E0Rpdv4unNIgzcDfNL4oKW+TD4hcFzYIAfmxWnXHzE0DysI
mnZmyN10t/+Th0J1BZDSfJ4EbSrcGyRnB0vFywdVgXs0lCjySjVy0YL/cSIOAZPbId+2X5fDmXDE
KLA9DW9Chp2f7CFurYEvfJlXHz6bj4FYpfiO41pbZWcKcJzDMEyfaZI6kHuwZAz9s48khO9KI0hV
2yACjU06aHMgrC8fs4BJsPcQtx5f6Fx3s+EndVN/lsliZxatjTGQe0o+qGZnH3/6yC9tTzHy0HDf
tpk5m6eJltTs2nBVefjKTqUc+PNTmjuto6RY0sc0gBNXw2SpIHovmT7C1KFTzA3Fi5Rhn0jXo7/g
rkznnlshi/PSR7Kn/bg/Fs7NBjdeOD5YJIHA/l6My+AR7kH2E0S6o1T28vTpaa8GnDb1Ix35KfyK
bQvdxNzrz3pksPhShneLQ2hMPL5RrtDosvaX6j1E8Bqtup5DUIXljdMxsGmXgqTkrTio3z04E+S6
jef88uhi5xgxEc7dJ0q53RavXcN90+3EnvvbwEwvt2MXaeHrFMreExVtBeco6DM9+O7s3g1HvzJu
lrt7HhoiguJR6zX5XPTy8PKV0S5vyWqJwYweZ3Xsd4XW9ei6qz5zCzOYqL9m3AOov2cXn4iNYXOS
JZ9sp1WtZjBPF81ikmTeBHNWNftOmFDKrA6ZVowqhQXB3FwLnHacdu56dOQwRfl8GI1Q6fZYsGId
95yXr70XWlddafHD1/2V1fc+y/IxI0zrvoFe8b1gO9d7EzM++crftv3j9XAhfUS4knPO+BbFQ/ZD
M0ErWIhX9ys2zMZyOS8Ldq9gyq5cizXBaNDEdm+GrksRlYN3xmYvux8xM7RzNH1PBLhcF3BzWb4R
jlFmRAbEOnDftw5mwcr/E0SMGPxHcQtbSr8bm3OWgZAZeoAyg6cXfCJDRgGpF0BPga8CnvFA+R+i
E0P7pl8w3eZJjTs09TEhJZ0pvUp2LN8YHwx+GqMHbMNZzDdRyrDlo9aRhDA40kcmFlfrL+OILLAy
VBElPHi5+Hlw32G7tBPBkCebt0bLDr1ZMn5l3e82w0aTbvNee7Gp/sy/lnoHWCWssIfZrZxe84/0
URXXgMVhcrJi/8zKHgzbeSNB7CUClleie5bw1r1+9WrULVrO1Ptnx0t6mH6ocAcDD7DckhEzRIfA
/d1IrPWBFsJn0YRRmq1F/oAA2MrTh3Xv73+nafCKO63hxasKw4BlTnMcvRTlW5GsTXv8bzyx2j81
j6Miv4bc7xhAYyIkDcZdR2KktdXVzN4GiIN9owOS8lb3ahbR6/CJMuTSoTgyLggXSAl1SrOdXFpJ
uDPuqVszvIzjVdBY+WVLpe7Hppo0zopNrx9dU7tyxZQaZBrxfsKa2bBUxJGAmLz/96Ee7n9OVo4a
VHdaB/qwe3UGIhTxDn0GalrkKxv65NWd9y/MgflDRJqJH+i0WwdHWiy3h5AOjki4hRpXAbKWBLIH
UZvH+3z11+ReCyycz/bTD5/BM5n71jo42TboKBy8d1UNazKNhKpS5hrGqIdA2ojhRwr3aBB2Dhke
QXz0ZRvnv2MNuKYm4eMB7jmDeWil9nYa2ehaWcVgFq2j8laYn+48N9qJPSj1ZC6r+5UL7Gnbqlj2
f/MBJQLJYVdm46yoq3kC2y3m90G6ABGjQU2byOgUX0cQ/iSGV2vZHVkMd2wcKv5iJ9e3bsOSwPlO
MesC+K3Ey1tfl5f8d0Yy/ZHztgcxCRgZCIOEcnvnHLVbBcmBxzNhNCAOP8tSzf225nHgGWCEEy7m
MIhxvVkfZF+gQwVNDH8jxHDvtKVyqaBG3SGo2hMFFAr0tkU+GXS7zqzP4CVKw0mhPD+FmaullwYE
jRLBB5vDIEUqU0GpjP5NHaYPlVhaBakFrORVVZ5rQcH03nbq9H5kbwzZp4YkS0wI/QsuZzDoSveB
ZMUlG53vReiybspoluhdk6mdMAKP5EwivhaMEZT5BCVlVYUMV745o/Zu2y/D63hzGDgyMUBsWlLj
BC06c0PPSYm2MwfdrPxAZ4lng8pfO3o6sINHQuKVxH1A2ZXuFvvoqK5h/CFjcnaedZS4pgsZhi0B
2y8+QHxjQVYAWxlC6+ZBhlHUC6RxNJlqsgfxGdN2gG1Iabn8lnCgh13DMqFN7p1XNwXJcDB+Da1/
apliB6wzYYRviCcmMxwdgpcAkDzAnyXqzsXgb9dUtyo5dT/P73PhTrytuZVW49FDUyO2vRdjNgZP
B/fmrzC5KYviUox3tF8uCVWY4oO/4PnF0PpFGrCUjuD29HYWi/Krz5IL7+S1maR+Ayp23e1i7XJi
RmPuOy81+gL4VY3aMXXGH5BGyvcPvOA1rdfNdqgBNF5zpr6c6xZMW/ngxMU/Cf9HHMSQZvVDY0/m
nxUvbSB7CtNZxFMR23Hvs/GDMx5rK6b+/hpwKdzCvGR01cECHb3TPPsVsO5/6qe4Leb4yuhUO4yk
Kqe9Kwl8e3yRYbcO/6f4l5KKN/PEO0VCHn9Fi5bJuPzu/At0JxLYe1VroC8ik941YRoUnD0eX8NN
rgk8Kuk21G+ezFo7MIaiJuxaSDo8M3MB5botx4HFw9XvlOyEa4wK4XugN1pMnsXg9RJ6P9qgDBJ4
WH/0XN0/OOypVnsl2yDgS8PFnVmP4KKuvit0DW7MyuBh07CoLuRgMLPTib++8uJH/+IG8psUOQ8k
V+Je6cI3Z+yjepo5ksOFPk0MbZT4ORQWHRKrYafe2W6TFkFZVjzcOY/quEtpZozfBTwJqnsJolSD
+AXiV3DjyYmpgFDyR7TFGnsL+lCJtt3ATv+O47P8RzAvF9Tpkrr8gz3ceAoIGE+LU9/dISnK90Kz
7azJGAeSxVXo2svCdOkZWTKCHUTUal5i7Pp/BzisVSz6G/mRfylvogErSb5HeQ8iAeip79/rbJdI
2LP4CfF0TtUPAgKz6d4A5wo0jiuEJCDC7NKO8IscyoKs/tBx3pP7kvNptWT8QHLXJl2WAwdP8Kpa
jD59g2PLM3C3nR7FRRJ/HNPyIRf+tnt62TZQlmpRDtSjOFLXC/uZEk03CHHuoBIKMT1Y7P1SIIHb
/5YLur/k/Z++hOIljWX5O6/vHPA37vthDoadkGKKfBfyx4XXmmfn1US106sp7O9uEFTN8tfdiuhe
GU3OXpSDd4pX+QKfyZx0wz8+7U17DUV7Yfqqo2rPsZpddVxzFds6NqGBc43ySEZhhGgKbH+bU1pr
ZvS4zyi3PugyXOygKpNK/yvcc28co0oYcTsK8IgnYEnzK5JUBHdCYCoJoXLegCi5SZyQB+2N5y70
bJWy6H1VUz/UQ1UgQ2LNcosMwLdFvVY28D6AC4INp4B7zJQ9iJ48BxeJvJzl/mPQQobo/JMn/NOC
oEttrKaVzA4Vegy3tNzWfMbMTDJhbfGiqCiCc7FmLw1yVtQnWak63NuPXbl44qkm7lcXUnaliNoq
q4KzM7yAS6iO23d8I9OWsVJ2iJ9C9jKEs7ID9twyJ5NpOsyySfE7NipDPSIAiC8Hd5K6GAL85PhK
V0bx9z65zDzWaxzIwAZpzTsT9yf5SYKiExbjn6wtEiZufYQnzS5iIuy4wx5bsRtH18snp0qBIPVr
xbhnCJynSnj0VIWu9nXEXVg5lvDlhkl+8vFiSsvkTiETu1qGrf7QOaAtuIUfrsfLsoh+NiJryI6x
cymE5iB2Ue7h7pLStJi8tqny1pVYoVUpwCJZnKBJsYNjql6HqUyLz9EDmPN8r1tKK0UD72fejXNL
jkCi2vioK6bp1kpA9WTr0ClB5c8DXJ6u/SfYrGtaswBtNaVGVfzVLfhpR4g9PCFQSiuTfZOcKGwl
clhud83Zj++npNKCixko1292Qhc11VpTgxGM+61ahED8eDLyWC39DSBSsNtbrQ+7A/n+raMAHLna
m2FL/G/L3dW/WJozsmREs0BtRL4wEc9PZDnTOObOyyZmion0O9FxRg6VL7scxYOgX9qSSbcrilO0
H4wO4FeuT+OMehDeo+blBR0ppRMDuBTRzg4VZkVgfHQQefHf/blEE4wEbjYS/fh0qUMWadxRXdj4
RLw8z+wZHhyWU7PnY7Tmw9P3RdgPxpzmt+VvZOIKCg98sEcO8IVOW653c6Vi6vgoG+E8/3oMLD65
U4Ro2wZLq6WuuChB61UcNASd6KgYC4oxZgAwrbQLQsdp/br7E/Q06MVDE+K9U/8bT2VDE9BUbEfP
kmLWM8NElsDKBnbin7l1yI666BVXTJ/KciXCWkex7F4VvNRMnRd8pojpj4D1MrqMDHM6GwOBnaqj
o3pOWm6suLBAHA92glPWpzktDR7E+sOcXNW/grCzM7HEKUmEZJXl70bXMT5VJIp2cw1VNbLBe5FC
3Cp0hPgqVYFA1GjjrLJ+Cd4vXyjUI9NzQak3PvCalDMcZ1VIPiRbaZqLqnQ+uJCE+8D/fUJfEl4p
KB0pAxWbZ7ilr9w9uCf3LOsh+90ZPEnPAjXF80pAhG08LGiEt20zFQg9CZniuyIaYTKwm91BcO8C
QzdnczM4feq4ePxt44VFEL35b56P0FyRbCB67mIICJqQ5YIetwj7XVL+nscTIrnS/KzsBzV8ixVv
crcYEws5C6iLvaL4tgaKUHtxWoBj7IuNB7sxkCHRslJSW+v3sT2ILiYSgpmjyYH6Cypq4B1JxBJi
Bg4K6GegtSg6pA9OmHEFamcehRQVfgP1c54pzTe28lscnq0L5as5fmlSrCdEHZBSo2ujahg3MC8n
qrl5pwVcmYrkEh5hBIbaScNYYsNze7nKryyAJS4yzNtHcwdvuyKIZMMpmVpMrab6KylPxOZYstGG
JqMOkavC3JYJQd7PG+Hacpc13vIrUr1rh70aBsjWsefWVN5dU+nMf3JUouZlsojL/4nivks+liGu
ZjcBiT2R4qokXR02PAR2/wDIow74nblvNEXcpXqPQsWVeuqsE/2yAWC8TBFz21i0Bh0iIB7t/40h
3lE8CJHc9c09eHO3Z4N+Q1z4rrxiJAba4sXVY3LCP6V7s3vaJGK4B/tB+Wq7yCDcUGNRVGhutmRe
/f/d7PlqfWLner/LHr6PocU1gVkERqMRUe5reGI3xfzdJ9zNOwKqWzpc+SAcBsp1Is+4JvT+uq6Q
At0biujUrJ7UA2od1XFnEwfdLhwo/uLmSiR7/Cp3MJTcyrkAOzj4QZK07jFu6DWt5W+QVXymIhvr
R9/s0Q4pUIiddtnDqvSW+NG7Nlg9KlhKsMizLWQO9EtL6Ez5FQ1l6qMDY6IstIi1vpIghlJHN8b+
bjDi8UusV1Guv6VOyNoO8Y06XaXZv8fPGlvQtOVCvwMDneWjDBWr1ccCEfZcRPt/wbMHMnHbvzOv
kWOgJg0ALmrgXU/vtbHHi00c79GjwT7sYUi9dLpHg6Eq3Yzq9arVQDLFki2dCuvA8D6ayC4a4V0O
qauxc9FugcsV9+DR/c71caHTJHkNjZf4w74zzAe4ZzcitN6yxkqG4BjrcyNXGHcEVPJNXKFJd3rd
dQxJsCOY/tFlUci88/EmuGDVd1TLk3k9g/GjJLzjCjlxTSn5JydKukhknS08wEsNWf9QCIEIIBtr
yGCFaal0GTcj5LNW1HucWCmy2+CmBahLA7RkiiGoVCzG++3lU+T2IekVa09Gq3Gp/4TglMKNzCQy
r20xJ9+Dk/ILR2awDPwHfM09sFFkvBnot/QFoZ4KpT3UZeBtITu0E2uS5/DsxDrGGsoksGMmF6Vo
vWVkZc5MU+52Vtr+xpaV0hpM9ZM8kSExk5GexLBwgGTrjWGTKvrXIG5jhd18tXKPgqYAlyc8fzHs
/W3HbROtqtN6ulHSQT8CI7ILeuiqOO8DvT8reum8ygJ0WXf5+//VxOzYVNn6YFSyDjfWnk397A8J
+tBG8ueSagTF4jPOuUoSfNfPQ13nPu1h3bIXWnY96IjcLglL964tv1zkOkF4TWETp+kloH3lGGbZ
sfWa+lcWpWL979lFdnHV247X+ynmWjjzmI67VsR+uz/4zRvcxHQLR5VJ0zDDktcHF4YegpS9W8cI
T6jXoPAIbGpdr0BzmF13qFySFyiB5Fy2V1QAaj4hP6MJ84at5XEjw+6q2KoyJdFxT3RLTKVT6Yn4
50sO2dQ/hXrypcshez7aALf2764KHosoLjpZEutvCIFS55SrUAnNan7YyCVAT402HeBwcVaUBxOA
TJ/Iztt/IWwG51ATJPlwA2Yf+6In7FPVeZBjHY+REoaU9Ve5JliPx+hLoJ2aPIbnHh4dIWeeZEIJ
zMeJPrzGPMnVTsKAxrdjTHJ4q9TBwXxV7h/WFM2Y/MytAfZJFTmFo+Q30n3Rg+iKjueIrvmUACN1
QpJjaNH4X72kMHfM5ZtpfBO1sm11Yahvctx7FgV4rs8dwGTEce6FdDqjPq4yTUFqnaBcoashsVxX
hfiHMJ4kOxnnKthlqDZapOrQu02mQfM/Fc+tiBKm/PlHGsheXp9NnbmotOdWvO/NGOkjd6Jf+Aj1
//flzRAZEu1OJF0ShuqpoXXrxYzWIT8jud3xQST4N1u/hYuHe8tqIlQ22zR27+EFmYlresajADOu
xyhQ4t1UvM/fQrXMOuTtJ8MPcHl4Q3W05WhmfXMUMyV0Leg5D06S7aXfo2h4nwqlJLQWDgMv6S8m
jL5B0U1j/1olTgtTOd6KhLh/b1EWD1ybLGxqdz7fDF33wkir7Hl6YOeqXF267ZVJe1gPMtGAW6ne
ZlK8ywQv14P3hadwZLJrEgz+RDSWf/me1/Z8OsiQY7fUnwrRgyHeOLTLVdTxcoIM4vVBN/bEgrVT
9IzlefbdFazaB6yPc2x8nzsaTwZGjZNCrxqJRMsZPRFh9CQu2+FLIU9KEAuxyOKJ7tnn9CUozc3Q
oYICUKaqtMbq4ltjTwzybOZK0TESsSqctcEhwUEhsMTj+4W2YQbqQtxLyB9SBE1ReBCNb+PaAUj2
touhkRoxPbzqthP2hE4J9skLrkKwJk1okUVPbdHTdYy9zS3am9sblpr6D5DmhLpdKf+xQX3jFVGi
qUAhDmYYyOIRcOWzUQj9iL+rcxy61uYuSkZ7UUrP0Vh/fQZdtkvek4fXdnKGG5ZBjqZKDyMP6JYt
Xabn0gWhgXufMoCJI8K/t/5p5HgH9eJJHdpVsBtPG/Wk806m6qCLKPjUQ7379C4mrMclIK9KaXVL
LIT9uG8JcDVwykTBndEQSB7QlaPpufnXISUqB+3Enifr/KqRTzx5ltE6fTxInInkKl3sG3GvqFzm
3ECGwHJvAfaG7l+Vo2SmE7dtXmM0FNZqMnYShXAv/aVYYOgZ7Qg+AhWiWPUodBMoC8pkCcxYqBOI
2WTYqnUlZ+s0ZEtDMtISkQnz1KaTC+h0BDgKkbkKxCC+E2hVkyECi3nUfkz4xrYkOvZgovVzCIu4
UjNM/1l94RHq2uNbpALZdSzTsi4F2hsS89LMdDpZmTJTDXdLVn58AZcpj4a/JWNcAhLhiKrq64Rr
4w4SIaGA6gdgKcp7Je6TkNMe0vcoL+ejfW//JmXdomGL4uQ0DnJeMjYMcymUi85gO3X3CGOYZURX
xa1wlXs+I7Fn8r62GZCgVcs5FcgMrF462cOVGcEEZeFdJVl+2Zn1BPPoMK/2zir0BOvwtToBb+Rv
tj73GsQUEyJ73BV8ykpRf2Fp+3O6UM7C02aBFKop4Xm5i47wT6lXXRJVzxAxKjjFrFkdY2CbbuGR
ncbxrHNDQGQpeZ9qSsMTq2qnkVq8B7eX1M3cBAED+ljWrpkO/xjDqM7l+peCGIAWBkGMD3le9kPM
NQCsOZwin8lE+SFZ9V9BZhPeeaFBxr6ra5Gs5QPreFOTa9HMy1xU5lPFdT/0u8ASQsqFyTZTLEj4
q2381clByQ3zpJUvfo3GbDlnpqsRuH71rVc8vKRozlwVdy6GE783IoIAesVwF7cP8RZXnLf/Gb5T
acERBjE1C2T9vaIz4FIt+w3M/du/x2unp2dgo9QweYxrIBdZFEffeubNrsgGsu7JY3XJ/eLM7Yha
BfR2j9H96wp3hvW33wkSSEKJWvH65KoMCAL59mfJNQIBFqR3hAnQfUA5N9wF/BCtkYP3acXrDILo
0hPavR3aqZ1oMQKinRZZwsZf/pCUlkOw7Iuzu3K4o9kh6f6di/LKJsZ/GPA8ygC4wTMrmpQFfkqp
PcK/anHknbjWTx2P7RDmDUP5yOP4d5Bg1zmjfYbWr+zWt+vSEyo7DYdS2MGIVQ3khOM7QvNEgftt
6QA3BLg4Z0GlfqNtJiVtj4cZJglBDZ7BN8F75+Dsh2UC2wACE69RjjawLQV2y83r3kOalbZnWQv5
EG2Z509DAIZLi6s/Jek9NkGZHgaczcOPaenkOCk5qYhMcJP9YGae9LWaXS8NaRgv8fxlDoe1ax3X
7jfuVxW3ucgyPzsRVo7PxOZ2PcfTHi/sfRpcu1NJzeIxXBz9Aq2cr2lF43iskT6CU5iRkRGiDsPA
1kYvFAl9nmCYMX41SAoXvC35Uy0fWzcimjpkBlZqDJo8eMsUxMSsgUox7iN3rfgClhS1T6HY48u0
kr0HfbLYNg0S6MO9Ar9pXkV7AauV8pGZfrB+FuTIkueg+pktkqYNHQQ58naFSgng3BS3Xm35YVBD
6zmvAt9b9obIgHVCyjtKzf1WOLiTl4brU9FtD3tCNhsXoJmFpWGb/boK1WOdFknEo54JUe1JaSH9
/E9r16oCm6oWihDyDbzp0ZXNkp1ZXqbOEAcU78ESox1THgQm+T9KMBO6x8g0So/NrpmQru/e8ChQ
kwUZ0PLoNbM52ivqq7gTNodTXF6NEidZzbk3BlM+nRGoBp5F9IakPaef/YLcwyuXFA3aDldG94pw
SdhIr7R0RbBJ0kR33GFjUX6rfesxRNfN9epRtKEGtYGqjFP4sXYBl+Lfk+oe7k0fu8upoJazka28
PqDvrP3yrVikWZRjB9v0Q5/Kh+tu6NShWHXWQmkM6f+vhPxAkSfNZECdno+O6g87NRlCXnI8ojKP
ap2ZKGXyu4dKVv1uhujBa1Y9D4LHJxxF06jXJDrhtp/ohz3Xt6sVzEstQkPVTa66U+g/S4IheEbB
nBXDv7TAtO0XEo0PN3cXgGIokxXMOqUj6i5Wn5vZ9XUSWwNOR8K0wVJiZBHidBUsbQidXDjE5Cnp
Aqxo9av88DICJy3Si8hNVfv5h80GsAtOpqEjobFr33LucE9zjPdw3Wtw0a29AiESGvx6cq1T5z48
w/2hsh4Kqvi5FjDeyhq9bcVrdYH1UgaY/tYCs7S7IxOljuuGW/9FBGOCg+z/c7t0C7dKDzS9ywdE
d2H+BcYiNRdAfN6YHXiGoavEm7od2La75S7WovytfJN1qZOg/DRfsJ7AXAFeUGtlti9Ij3GooEBD
Ubhyejyf91Jz9LyKBKMv69j3Hqed2LOCnWTFIKLToUPtZ2LcW94xJX/dmyyD2NNAcTh38tyvaAmD
iQmPXd97YPs6DTyo48h9WHYyB2SHQWN1jqODb6z4H9nYV2SltDfM/G13cre1dbRSdIJDQir4tB3O
2DznHB4xcrhMpgC1f/KYc/g+dQjuf6MTVy5ZcJXbpwm+3yPAAkBH2Zu/AC1vPpr1yxGvJPALbUg0
bchUPtvIhRspQHiSEGU8LlCEyLGyNNH1La53KmSNp2ZN5AUBzXCZRnzk+etshK41LSMrPhWA8tj4
cEtjKr0ASG1DYYtY9f63PlDqxeP/B0vOwieWFTRY+17C8tgdbioZ82v9NKNij6NZx0eu+dIAzUhj
fIGzaPsRnxOFgD+lipkG0LmrGaK2TXwAeQ0tOrbRIEQtHCoKvXHbSqcHZY9ljjOuyx2aDbtxXtfx
PQ8C+ESxeewuxAL30hdKsNsuRnDTdBTImXedbwWqAXG1umWr8gleb5P7yRGxmTaWbwm4qn1wZLlT
pG+if4KD2Q4ufk/5oaUb6z70NOOXdndaalw8VlDYDRMLMBjapM3D1mjkUH5BfnDwLBuDMApeEoGM
bF41sPlwGQ2GSdxSc4fCVpVswss1y5LKWqmirMfJy8gleBU/2Gj89l8+hNHxMJADPZ7Yi80IWlR/
1zzO9bHe+r9RLFYQvPqwduQVd/goy/SRcQAGWKKDcXyjYCNMBEa9W4iOWao7E2Tnso2j+YxToQEr
4hrucXAvI36+2elHjN3KWr1B5D9gVURYrW3+1ywZ2ujs9LoWMi0mWlN8BwrXzsc9FhUtWh61rbhB
97RgnG2O2V2mQyBJvfC9V7kr6hPbr4BRSa5ph/OYCtwZjmTrDSOI/+sSBNL/9t7v2jMnLguHhxVp
MKZJGFbW0qzP6ZhpPQYfzCrvKtXe0Hz7IebyCoXL6TkgHh529ni5o/r9AJHE4oSrOrJO0ZIgkbpy
CYJ+3KU0M6hvf3GmnGNKZ4ooOE3mh/t/rRABoKd5v9BvPATzn0ai9d0GEPemErEUU6+setagbMLE
IT6X3xlt9E2LAm9428aV6URsuXPLtVwzKkX0AY5P9Pm/7TjGNLBNK6rpYdP8xZPZp3QRHAHEknta
EMCcdeH1a2YpyXhHE2lhxEXHhQ7Rd/5iEkRBI7iBAYlwToTV0SM5m8rRrdxacP/NAyWzADfKfQg1
8In8ZHkzaIvTCP10VpOu/HHldhzeB4VbfmjQViWZnCDaF9X65rMTxPaC27uS+LTpbt3yX2HYXr2M
zXHTh4B8Nwume3i64CQU8OpJH6/XGK2WiJXZssRwCa+FA88W0018iUXlvxR8G/9T0Yec5Yysr2Uo
e8EXoP7zmnEksyGoXcONypYXldwMtiHUg1IkHZOnohA+pQiOewryJ/egE/MrM2a0pMDcZwh9+Gba
6UH9wHHRqvbyCWoGWcfUFNALY5QRPNW65nocakDpTVVNqTJPhl+KtILIN+sqbGzsxnTnYF4fNWpS
6iD02Y0faw6t10oy42fI+uaG247nUIQLnf5GuLWg+pK+iqX8M7HRt4v+phQnkrDp07N7g4PHsLwl
BnHedpI5j96CU9/mCe+tZXHSigBNPfYrqpQgS3sp24OUX1U1y5i4sPXgblh5gzG+46QF1CNXObO7
Xexu6hQICsA8sgUTeDiEX1vFjMSGmVYiG1EhcXXzJ4yhF0W6YrsawSSZhroDoGuIw1ACl6Q5elNY
rgc7ulatjav/u0Y2rL5F6TkrhiISJMRcRi0fsLjpBus8QoSDv9zatzeGJc2FVug7OMZ+AWFIUgwX
YG07rPuGNOYWLqRKIJELoUE/havdBH54ev61PhFIW09vqvzwBRWu+4Sh40qkDmMHK2Zli80algt8
wMYtPdcI7wwBtUajB2LuG23Ec52Di3lcGuh2ogzKrZMFi5VNvhKt0X2vnSDvegaCyt6ExtOSDUVs
09Ax31RZsumKSCdlOSWgbt7UuXrDhpW/vaA55II/xqfw0+OK2rJ9UajxC8SHasYmtWm7vkpF/4sh
Gi7JmZ8ii2s80/3hbgTXZbD7kYIJxEzvIf582Y1WLZXtB4brgl34MeX+6wHn3G/t/tvEGq8BnzfZ
+KKT3Vq9LnmFbpoYTHOYuW4PZfEZdjG+1w9todi+n7VIz34WuXYeymuM9KGhYYmoL9rUKs8mCyiF
Zet37jNWdTHIghJBGSWpytafNOPUpVbqJKnGrJ3wk5zyMpNLYvJm/n59WSRJC8+jYISm1WGPH7lH
3oY4MZQCuZP70Jygf2MrN4ilVhO2lME5hLwfNZmNF3AOV7gDyYdG76+urDrxqoQo8sTPB6uZ2r9w
9j8iSXg2aQPCkNzJkuEAVCyplBRQgl/RT+6LgHBbE+65hlg9ZGiKHevOerUXfWHSPpJc+xRniohG
uer4kMfGZ0dKYo7pKVoJemVvIowHXjcuRG98LytKgHD3BIgPUhOYe9080DWnsYuWQXHHuomC9iiR
XAyqVJs3w5TYVrGhlFZvgJI/iqXXWJpGMkmmLga+ALh13coZJIaM46fQRtxvb1cwHKao6i6N3IJ+
10DQhD1q8gn8Oux0RUS/ievo2Fx5bk/e/2HZQyzZFk6jGaBHV4sf2C//S7y09aZDiZIr0ZCxnZ+p
3Hp/AGtiv/9qPEbqKTiTkedZBFDkxhODrOqqQ4rdwz4rZQdzsctr+bKNkpTCF1oPh1ihhVC7UbvU
v3rcnevGDoGJlff2vRWNiuGXZoE+qDJLApfnSbceTlzXgHe876Eg9G9vIpOJNxAqeRqKbRs/3YlP
9Adl0ZuNbsPd2Unam6gmPrGql6sYFxAd5vAovdq0nOJ0XRer0wwlGJJErZKyMEFeu9SdID2Zm/KU
oQg36KuYOZMMkHPJIuKJy90OLlbtWTGKhXvaNfzr+EsUtnrhiGvV0i+7mMIc59HrgEbpTt1oTiz1
j7+SHKyJXPOnFJviQrep2J1wrirgEW0JTA4of41QPuEjSyeChMMau88x2Sg9i9V50yETwKm2wMGp
XMcCv+secSC7faNQYKtOJKIhGCmguMf0nEp6n/HFU16VSGoZaeRmiaD33K7V6K54WwPvQcyb/2d9
mbBkNgFGol1A6QoHI5cGLy2dzmuqeFValQeT0gOe7Agh1U4qjpklZe4LaUzjaxwn0gKNY7XCp56m
uIvsXuBdBQ5Xt/tM6m77x8sn/pvfB6BMpjinJ5AgkIWJ4oNrE77gGYNlGmEfy8M6wcfYXk/qiDC0
17N3Yfoz9VlCnMYJbuuWMi+N3fiv+5sj7m0LoU/SaGuceH08VL/caxJaqVjTqmFyoGlBXLTewGJ5
JEKvwkHWi9h21/clxA43RJRP4sD0bEbL6uN+EmQ2n47lKHmkv0VQENUA9UEDAFINOGG4/Ff0reRq
JXhmJmqZF8gSZmBvMx/Re0si/gLfbzd3BJVX61/1uMbNlOB8yoyIai+RYTSIewQOSeipG3HO7G6b
MCIhAFPGp21J7oJcHXXsZhb0MPuGqmaJjCJ/PPdLaB+W8NAJQqLjynL3BIC3kcay48PpVvfA8wAk
RIQobfainB10MxlFjN72BmsPNLH4gExPBZbuB/W1VOABp2LGUpq7f1v5c56+5PLvsX3KOzDcSV4f
OrJf91TZ5k5jPxqmnsaGuRZ3ssf+ZTgxkG7YLZiyOQagD3dRrqPqN9huhNC0pYcRF2MGHERiCv4t
FnBpjyeo8yNEiVLc4X351waYXZRzAp2Pd+gUQne28DzNSAQABjNFIr1VKEl4qO/x5Y1ALRd6hHIP
oHgS2SBCX54cM+Yoz+WSq/gUGrJMFQ0sE64YM7noZSgBlm9cAkI7LJDYgd1TB3JHhz+iLSA4v6uP
nXqV4VfgOkoXx1hKZPowzCJb1tI/cNiXKyRQe86eVCzmZpAYmPMFRPZadLzyNfjmvVwyqq75GjYy
tZ7YIbDlwQ7NXVpk1ifLmtiQmwrmtdmeJx6Kipjot3Tsq0ZL3J0UB07PEz8aXx86SDj5gY4w+SyR
gB4aafgsxgP9Epnj1Lw9G//ZRxVzRRCdyi/TiO5isfsdynB6EDh4EFYcJ5xFBPEILzNPk/U7RZkC
x6b5d4Us2y36uThGVHQRmPCfOwQGSwXn1+BDoike3aIMH6vFABmo7t+xTq4C8l5XC0CmvCO1Nsqo
VXnxENdlbDm8d9FX+iUKxC2PfQSA+VcquPwLwgtOliv1u7Nlm02tIgsW2X/n9tYVJooJtztvXA8z
sigfGhY5pddQ39CV3MmDuGqY/CcLzIcv0rKU6Y3BF65fsn3s7g6pvna0vqGDZuQNnbAKHMWPJobx
lGrMq/xsrXOHAX+5sVYb9NSwhDtyDBmqj4FS0uAgptzddHyh+b+QLzesIhEwUXLXF/7EiMfgXFbF
q6W7gU6y6MdCIj8uuZTBhhvdcNA9nX8ZcE1CxOVuSuPpcdjr3VrYsaro7dDYDZ9etAhDeOb/+2/y
7N7lAC6QO2gi347jPW47hAqFqf+CiwAz70o3dgQ69oOrpuuzT32+WOnvvTkDqmNhzTQREnuyFegU
eEn/X72z7sGO3JaRno7ZMkpRNhn6gvBxz/AN+6MJtNjIEkh06sA/cV24knn9j475WEAvY2H57iKI
N5Im1UhKpWr/ebcfqCPhmuQQDwvYyti+0Eb9ZZZaChfKpZdznoKoQLiY1a4sy5hrXZbvlY8WzA6y
kmrUObTkKi3cp02TB2bqH96d3L+CBD8z9KMN5Sz3AlJx4V4RGwkfZNz5MZTN+HkuPhvmchToFaET
bYrBtTcwXsxBysyIsnjGiJQVbZN9Ezlg/TUDVuegRb33S8W2MUGMN8dqClLQX84yUcyC/3b24zMc
GM5TrMyhNzOYxDQ8Px+ajhlq2fIzq6OdZZZsKu/HCZufQVcWShrp0CmbWo/2TkkPoRtpFdbx4Ryl
ASbqmbbg2KpuUgy98YGec5lz178eDmoYLnhXw4u2C0ovXNgJrXGnvSUa0F3ws9KTPdJeUaCloxsw
42+3wJmjlTpOV5ZBXPpyappJXpa2DD/4DvYL/50WwSVO27O35rslNZTvri2+X5XmSfrbxBvwcqmn
g5M3azsOibLVaJO/+b0Fl6ruqFWUAPGXAX2JClAFc25UzpDTkmXKzb0qs6Ri+rchn1hRy/b+am0w
gv0J1SuprAaoGOBEA3zMUEr+EFacyFtBVMVDbuzxpQPN0klYf3DJkETp3/Lws9egITn0nXaCEjuM
TFxw+BT7JyTl/0Y3wn3zVGDHgrXe0CLnc2rRSmHqZE/c5h9fjWnovEfOBik/7Ons45pZbkqewkX8
HApEJGo4uMKs3I6wWYJNNEppSj+8hT6NhGV6Xysx9E8ul+HpWozYE/A9rvzgkhqY8E9xRvK8zjFx
Gp0mJKMroOC7AWj/iYeKvVm0dcgLrEtH5Ks7p2ZSRiMZo5kTrxyXL4fU20YLg/3eWIHRUNNFV0W2
NcDs08KLg/9zy7vgLs64Y9U9GbwPDB/+XSMpMXHjAagsRoP61WZmJY1ejI6LMcn+GbOgIGfRTFoP
2ycQQatQSRdRy9oGNT2p0aajHm81G6qMiQlomUdc7Ee8dBp0nRK7TZaR4Sc170roP1YsNGjGs8tc
lj+uJirrx91HjI4l/rq5eXUe3Q6XzvstOicrTKd/3+hD486au2Z7f7ppykpqBNYe3eUvrmT3YOm6
GN9DoQ0+S0TMyS7rRVEgTcFmj5oQ/sTPino0Yt7Kbe92S2HtVONyx3UhhMuwpt0uGUFkY0jUtJ7+
M1ApymsBEp0swPPsdM3b8Gm3UKmdslaD4azp7pZzrYbW5N7e7PRgoGqYNtEPZlY2ay6ff+wEHTYn
Py+bnUZR9Dh6s15/oFFNxKOw79cXvujlUvH08XXaaeBjKheikiaxG/k3aiwidZNz1m2LiyOKwbZA
iLvI/82OnxhR6WNPHt3+zErKUZsSvATw0t410qOvNmcbMQwvDWaAibNwwN3YYfkQHONCAl46pTCU
z0wX63JIWj4AMbWZHH+YEGLQLHTMR17Y6nLve2mLlzn2b0oxnnfNTn2qr4DpHM7qXvQuDH9zqMCQ
Fmfl1GgljSGEYUNe1wnGTH8iYe40Y/ytnA5Rt4uR/ZtEgTGMe/DQ7bVclNPTHRgG97YFU6QBpprb
bjRADoUDoEuloxlkav5hRsk2+5MO6RByrQLPVi7AjLyM1L+nDfACNA9SrFf0fIdmTGoyUeD0i82W
5VcTe+NEBk7ItKIwf3SDlAu83NT/qCN9G8dwoAKGs5m8JfmWpwdNA4juOzCwwjZmzzi/cNpDA5r6
HaB2ladKcU6RepbrRUajxd/lIL9uz1ei2jzHNQGjoEnYwhX0Vqg12xhALrF/QzMo4L5UMKHNzGqM
lludGwp8dop5p1W8sESO4K8eUZ8iIuDpzZrXm2D+nsPXV9FFith9ETjhqWVJoq8CzA+DBZlA/gUe
3i1+gw2F8G6gSbu6JrDRZr/iH302Py3JLrvgVvhxNnw2CbFw4br2pjkLe8kcSktVPpuKap162dsy
Hr9E1+pNSbRqrdWj+xW5YTYpv9gjYg/yUzlWW0KQ9fSz66t2l+NmFTUiOza7r8Nh5WZdsRyWg9aP
GYGx3fpuIxixszEykycBLZvU49Do3lhsaCpelDdLm6MftVMwBLxyO+NjUHKGl5TaRmUupoU0CsEx
REaLmQYZI5J8kVav7ynPH+IhoeQ7Cxma3PmGPJIx7gSW/4cT0FQeGfWl/LGdPFp+TUMFNU6gvJas
9meqa3GAK1J897SXY9qDdt8x1gd9DlkhJjvRu0kyuCg6oexqXcNbhHmUruoRBoPebFASb/liJP2O
LuRpQ/Ab3/QZFAhZYoeLHnNAE7VRyUEgVOjhnMaJHkKmmENPkBC3j+ZcrVKVQngWJ4Sva2p7onnl
1hCM2qkR/vkIsqRVaUuzjoeIHHt6FPBXCJVZeDBFUC8wbVrsNbIq3Ss1+STqTVBTvy+qGxql7lDH
4Yj7XjQeQSRAKrXwsTOL4WqtVoUSOqIrwY5lwGroxm4Y2lZS2FrMSA07tW1YGkM57LpYjg/pGE0K
hboQrq8Xk/cJ3RjAhet0p/gthTsennY5xP7idE+WdHeGGAdNGXtkSPimL4Nevw1oczxHeH4zq2jX
biEcj0Pl/JzOgGRuN3zg2tLqXgm6cI1ReW2RS0imuip8FQe+mwRL2NOPssHQVxDYzY3Z3BLAqBiW
GjMCgjMCR0a1q1s+29LYnzzpdjN6KxDw2HAFbTjYai2V9aI8Wa8Xenxbp/LDDclGVt81pFzU0eoN
NJmlHxH9zjc7wkSCNttDr5II1ammm8llj9CNRua2x3zGMxE+TXksHEpXENl81AOZU1+K4VL7MRfg
D0xW+yx9i4u72M1qhym5QiVbK+fSDMwSt8Hx2SX2QYqJTgWJWIHtT7yHvxFvgKAeNgVO3oCnDaBl
FcJXx9lSx2nsji0f9vAHlM9JT7H92vvloYtsZB+QMnfMshwGKK8FRPvYSM3FgjoNIr2DWBVOiX0v
ltqsFfpvUxZJBBxhFdPQjRbUMEFOip8bmpgqrRcetBQhLzi+0GpZRQ6U2gRoH7HppeKdBj1wC6PV
GVXB+uOYIMH0KPhWpYCUHJY0uLS/9pyMl2k+/ZVo4oqga8QzzwVXp18cE8CSyma9oxm2BBOau2kS
IE6HPLlLdQtqY2qo4slIWaCspL1j7Aa/mPfjWmVofHE493ZKB87vCMQRFVIDTHGgsLrWbq+x4reH
sisa1fUUSd3FbwEItPQXx2Mq2dbRDXwI/BtlUDJ9SoL3sEWx16Hj3eJnTpcvYrT8BHZwalbMKXel
HULyXbl8EO71I2O4dP35lrr6Wxv2en5DyR59v9korpg3K5jFTLPACSu1RFh+56YLJAF/lIwFLy3x
7XLo1vqH+T3nxssjQ9bLRd+LBj+1Rqht7v1tG/zj12YRrlcPZhZPrO9/27oWl0j+MdUpa8G8lus5
fIJQ4Zd2FAWq6ECzsIzJfymvtUDkl9uyqJRxYMdIbL1IcCZhQZtySnjnXFccQb5kTxwwiZUibmvD
YLnjlVYpnQ72/TYcAYeE7R+xAgxlyZUT4suArKaXJoalNOKILEhmmsy0fPY/wS+VOAjMwiTKw0Qk
C07SFkCs2O0DA477jVU6YXzQoGkEmcBpy+m+fBszIPiGKrgRl/hEbBwld4r0ZhNGmA8ppb0L6VhW
rtqY2gK6TpAe/xn/nlKwa4tbrPPPqbO5Q/v13U7A2KGMVuFbfHeCiCvSXWNJp197vCrAuzlB0ei5
uuUHplay1CpMUTaASEBb0CPFKg72YOBwmonKqDg3Je+oW0W22MM+RoZRkEVxWRdsmoyWFuxnvVDJ
2YAiK2/XLu3Gr2VTRIHtQul+KenNObco9wg8No+TRLqJlGXyvEXxUNtnGEPBhLziuEk65pTQuHjr
GYN2RX4be6A4dLFxERSS9S75TkV7g9dxTh9+j0ibfbJZ3gFtvzMcQN35QZtmfGoUT4+vh4/a1hEI
cJsCSvrj/AbO+VzS5Qe8Uqutmx+x9ad0p5q7uU9ZHHfH/ka5DoWstBK46N8OGjZzk4D6dvqB7zKl
r50za3Ie+1QBoSrG79xFnvOhDuIsWDeR+t1sFXVzwsCt7XtDTLkAhEwegtitNCrKST9c7iRuY08G
JPkJl8+BnlkrtwMxFfTsBWFy23CIHVtPO7MUfdyFUKgLlDII6MmScs13XVL8B4JS2Y/GsUp//ZZv
6FfW3ABmvBXH7D1mM2PgPmTRAze2zRzigaCJOaEeyyFT89Muu/ogIEYXWwM+59qtRiMLuwS6gx8o
8g+AMaYKEOQXj2msDSvffRKFCDOgoR4sBGPOdGly4UhcRhc6gf1f/oxX6UoWWfLF/96mVFsU9gDR
YZxyc6JblcChSOQkvy9wK+q9c1rnjssmXQ4VdbqYtshQNeToDGksVP0Z91PB4ajHnsMeGuAv4mP8
kuFN7eF+AE2pcz1w9ynlY4h5X7cldHRRPGQZsSdx2g9BEGulD2mu3Feofj0CQyuMmYh6acdcw2DN
L6kP6aRU1QBxQ5ISG2VAhQt3Sqwij1w1Vexff+ueFduLljXqOyhgYeMCDGPMp2HpEOsOwCyfzODq
9aisB3qbYgX8Keu97nRsGYY3zohGjos9ipb5/SJWYWBpZ3dGoO3IlDgDf0o8eHPIWbD6PbA45J0u
6IaTff0dA7Fuq+4YkD11LwLxVO8qr229uHcogoya9+WbXuGRyY//fkEzM8L3yFTgUNIkotb4BZQG
YcSYEaY4NtrAvznnXxCZsTV1ZwyRYgr1fH8ow+CxEfOso2dIvJoBnjjT9aTCkbmd/4/iAS3jZPk+
w4x2R6AiYDxqIy/mJjxMHGqnjffYfJ1f3CO8AJ3BHcCRwzcfeRvRAuZDh5KUTRI2mrhLxZNUGvYD
7allZmJ3YeaEAIfghfV+HPrNu9ooAGdViP87ETwSy6f2dTwMq0kKwJ0UG/YGkj5XqtycjNX3UU23
qC5s40vBzSVosPT1nBek7bEoWDeOh0JbGT+08W1aOrNURwDBFvqxKS8ZBq1BqKzKpWs0sqxPpn6Y
vCEAgXg6dN9OaXdLBgeVhR2FgBsLOtNN0/AxW5PaajYOaFecohoF3VUZg5Fgjye7EXiervGAHtOA
JIsWEV5Gx0J6T5vNBHpwyxvHXerzZQyyUNYOQVie/+iiv+Wtwnz++VlSk4fQjflKAGLBlVaXrXxg
W1lvsNUfot/J9/+a+AOBReviwaCX6jXaAfVIZ3MrS8F9d/yuj2QDzJQnFI1DFnAPO7Qte4n7enev
Vp46SDFipFvfmKjenfUHB+rDV4L9ZQH2tCeMAiqMOFtp2igFINWM7o290ZVFnaLmDyrSWNjuL5MH
63A9jY/2CZFkkgYNPW+tfHPFSXDGgsQDgqhsww1WL5gKt6GriXOSV4ZdvYJaecCP1LTrVD39tiJu
Jug0VPGaYJe0ZMoNivVcEidU6SBZB6k+M9NQdzA06YIAQRadfzFcp2KhQ7TgNolg4Qv319TWDet8
lTMxpsfOlYbPhwPsSO7GVQd5dIdYtUFt7gzvrB8rvvW0u3qeyOf9SQ5XnmSqxXKEUGHWRZOryIJY
z8YEQVrPOTpc3zOKwLRvOVGr2UNA+2F4d9q4LNxmSxeknGqMuGhXG2ucYadfsZ2D1UmA4Wj6uTC3
T84s6CcRdXte7Y6MQvCN/WIlsmXZjrfvyHKFEolcdr/GtNrFNx3fsrZ3tiUCfbKIlE+WMarp8J6x
czHA+t6rijxFfvbku1NEAFVeP8xQ8tJsuOSCJ5OuXCf6PAoxVrkQF47K7PxZSbzAjMNjxux5gVj1
3DsULtrSdg3MO9rHejgjpeLn0EhaQQBR19IIe/OjjFsSMxkB5h4HfepVx/eXs2ijT2ELOuOZC6rr
5IVzxgQAC3LZvnACao/T7B7out6Q0Zw/ko0zExrxaLeeYv0m21nO5SkeHkt/SxdQ8FXwGL8H6SAE
ZSuIZuIFmvzaqKG3M/pjbc+w/vC+Z19Wpa+m2DHoYC2yymq36zelGDuy7DLmxbja/xf7kUY3KR7A
BL+nZAJAOxVs5DAmW9jMlGI2xreEJmnM/aLInxBTvAeFM0cgO7Uq2W9EADMvlLWOuRhq57/6t3r2
FqLavmDMa1g6PeiC8CPnOu5vDfH02fAg2AKHyU4U9sHe+Vyv+gC0/aV2numlV0BcKEEzDIkgg1AE
HelbzwnIkvtkuYUDC1Xdm5z05KYTqWQksPefZGEVBLIjaNK/TbKxbfIHItQhaR+uQzhyd4vlo8RN
aWXAIDLtDsBB2fijgx4v7TUhIMCMtRlPgGaUZWT80Xf8Qx26NY0x7n+M8BsxQEDbazSio57bP3gE
cYaOC1rvjnXAZUDl7pBIh5Swf27Bg+OHiNtMqsdqHIDePOPTFUWoGENWtBXHwHjFmoQMWmfCXlhi
U4K5n6S9G1OaqXQXfaQMLuOlOmurrlnsK4oJYCkhSxc+GTb6ytz/2kbILyS5GDmgGUYDJEacUCp0
XQ4evu/BXry3JZRz/x4ouQC9eI3Bq2hpLpPtg4GvC9k2uLRyLYwr7xDTw96Po2M58stF3TbtWWgJ
bbOZEJj1T0jKlt+8Eh80I9M0Vd+GSx1yVg8QQh2l9Up2BTJ34ENZfAPx5Wf4uQQDU0R6aIKcGft8
aYTEtkxUYr9+VDLYssjXSY6j/2cxlV3eKOMfkdWwCkwBFg1FiY+ckVMLyxDFVBdxX+aNpYZgsnPq
TYH/0f/UQjg9jubt8WRv7eMeKKvn9RblbJIZ7tVhrQqnQ2N1jbFHks5qUWR9e76fcaJMcWcfmLdx
hE7MESeY9xANf0X3j9ww9xGzf2FfsiAtm4QvzAc8iGGC9srMFCJrOw4OPdENt6p+3ehXFc6vBB6x
arc3ASCUGxwTIVv+yCRBpBQyx0WN9IiFGoyGn3Lhd3xo+u0RuDjP7fEYqF2IzfODSALdfbvkHiO6
5o4/XGT3bw7+kbwi0w0O1+5dKpelLf4AkhdjchHlendIjK2oaZIklN3UD+jUaFpXB4Dgz/xnS9v2
badkOcDMI+kQ1DzslxZVd3QyGGWjMgcmXYV/imGsZM0vkWukXwx87sq95OeDBhWRtYY+vlAA/bgb
uEIy497F3QG+8741cJ4OvPn+llaqzLqG1CLy/yWrfqFm+NqjRck2AGH1bEElQxbJC9/WXrfsmvL2
zqIQ824ZTuEg0gt9984xJZNXTH8rMIh10s3ayLBDbtCe91SafRGZ5sG6OOU0Vm2IJjHI0wL7Ng8/
Xy98Wb0skwf0yXIGiIzD+7vpiIzMo2mQy9xPW7O0/VR8xQfYM3LCtMRLBWqXYJpQxYK0BjnBRrn/
iZIPasT+oRpAWNQPCsHkq8rMgo3xb6g7Tz+SvHyEp2hNbaseU1ooBszBiAC2JbH8rvbylco3QoKe
Aeh0opCQjhHTyRKQBTEQSnmiks0MJuprEYFDHBa8hD3qbQByOpjZiM8Y1p9+36D20lK6uADsfzKl
GGlfoPLXHcGD9msH+fouvMd3hpkjQlf0j4OMO4U0MCkLAySydX0oe3dA0e2XaM2n4gwibDPg22OD
PUPHUecsNKYsG+lLqNTS6/HZQmPtjXKbVobFbrIYA4VjFFTgHF8nNDaXADFYkKyInnegvWVuyD++
cgGQJ9qMEgD96nhsap8jNYZJF39bSe1seIviS3f3g5cv+CY9Tw4X4pGGPGbbh8bKi4GMYBVjm1WI
dO61LxFzNX9mUSikv8FSP1diAaBZ0cTRjkDWybH8XZPB1VprvoUJM3bzrFGQYDBM3OYL3BUC78vw
XB9wQvsyDBM9+bCdzWw4c3Vk1YIYvMr9ynMQU2Iw54gJFuL/l0Kmm1lTncj2CLnQrumYFKtmFOwp
QC0CdzQHEkkHGsYMeQnvTka61+Mk9DUUCpfl+ZW27PMyDeJ5M4iTmY3mWlbNPXJZQqAOFYrZnsPP
tjWhTTRcGDQrcdRnrtcCaybiNIIGPN1p1YTtpj0KaynERx7ZaySCCHaVzcEIl+OtYcUMM+77DSGl
rT3ERH2ZHaE8lSLy/AesSsOGkFr4cvnj2AozjVbF8xjYLsL1iToHBpalhNH7lLofIVFf3WPGmuc2
0gKFm4OBYaSWK6oZLZGBN4Z9NWZJn0VIvPi33R9IRLRcmt1VtYcTHSiOck478G/eln6a8FoQRt0Y
YfPRCsnLyosH11yB89C296UsmnAAO5skB/6euwXEt/4S8HzGPFEra8/4S21Y706bzl9NCcEZcW/T
kHOqH7gDwIo04p06fD+aS5B6ZhAcryMiUQoCHuGcNZzjFg7e5DsRjoVs9gpnxOZGooRh0/IEVktW
4ZoaAFGbMMDzlNPYBD75zQUJszTA0I1sFh2EED55OO5uQDUOk2vUuWdzJfVnL/1FdANJ28hOUzFT
1E8sn5vIEjZ3kt5xv9sMxWclsvdh178Wi+ZQoHXthO7VFftSWB8nkS1F+lsM/jqF6PJCvArlRh6k
+NbEtncW+tgLKaZEtL2QHOdVfrCVW5jICe/KU2CsI6yXp70K1dwtpn60dbHXRr8Wo1IJePqtJ1BO
vTp65BvXhIEuHxV3ykkwHOYSeACHp6Al0PY6vlXqbr1axX4Whif4F0BKW83fvkX3+ngeYMF+bGH7
Iphkt/YNNzplPpLram5s+QOTRO+6OX9wHpztoC5mK2zVDeURJlnE4qICGmBW1/KGWX6fcxa/gBWC
Zr7I/jdSk59+VJekM+G8CLDb+hua1y6xkBQIhFoSPR0LlIfSk3kuFoOwBkGS6XSS040flkqHsMzd
wjrf5gmBlkiEl4jl0LSqBiLDOFQ/VComoPtIKD3LyIu8f0jdvU+9wj/o5DtY0cSh2oUQYw/84Q5z
DQWhw0HFFIJ1KUfYCzcydSgEGcheVmZcmJkMjykr22BWNZvr9QXRuCR0q1FWXV4qN9LsQDFSoPE5
PdIKWGTLMbbjr1dchEkXo9p7C8T499aBMmqf4ZAzhsPNyCZLB8A5Y5bD5slqHRv8NnQjR4WSzkqD
LVxZB0wlHauyR7MtcWIpgwe5hJcW8tFmHR4LkL+sXEtpV3/77r3XT+ezNPW+v1pJ26/P+Xt8lv2L
+qUhHy1ZNfJXSBzI01bZKQIEdC0zSpJzhBfamdtfRqyUrQbxue4O6l0r0ZiDc4x5XM3dox+DxUFJ
ICUo+41Yoz61Hn6AQhGSuwPHN6ZFFNE7sDjkxTr5aZG/WZRm9+I387muTLRR51GYI8XIq756DXv+
cmyyDnCB7blTGvkEW0Fd+9Q0kq34JYCQUW7EnivfeG0n0AWj8kK7yg26NCT3rJdwvrVGtK5RtgYm
oAo1fIc/eFFf57QKVgGy0QksamxrpW92K8TxX0P08c4t7MS9F0ApHkTzqk1L9pwuvUbGuMtDZSdd
MCamBG+ewu2SMn2VYeNCnZpQ/JpNqGj2+iJkVHzK/h/PtObtUzZBV0jF6IKx/wTiwzkpDyah5cuJ
TRdMnAL4y17RfdPoeC2eEgMSuGfnkXt9FbLlTtTGIs7utPut2f6L+4KwJkQkVC4hOGzs7OfyxTiV
WuEiDc9NFs4L9HK0/3Pz0wpPI/qTXKrWLgjtgonmwGyL/N3mp96+UHXbWcOzDR7TCyFTC5rr3jcZ
/+3hTPe11ssjsRrayiE02fpdsfpvJTa6KrHF9U5t6L2U9xbAbljjRDJCtJZGmybXXlXi76ZB5nwX
XYzomdU8gvFBxBun3tT7uoSgTkR1CHOuM1Y558tHQeBbMOtX4swkp6FD3/De99z+iIVINsyRbDXl
HvQl6cttTGhtD5Xn4/+BceN3+9ikPSTUSF3XpYo2zZfbwSSbzshLDM8PgPLr0/wkq/k7SlhCKxPU
IF/vm7nDJjLJaw4C2nEZwdknl7ElvzvYVcooS1bCu2DxJ7LjglAYl2WlOHfTv05ZwrmEkLhgzNlQ
rg8jCVs2zXtJjVyMNIMSH1dTAVUYEPGKsLnmNyf2IgGCEVchs7bOg347Feiqg7l48m89bD1qGOoH
vNM99X2oMAjgt7tULPfYXT6RnYhjf0lQpE1SDc2FTnG/ya2OcNsmEzwjvfKDWDAHSf1bNBTfJtnj
jLNYt6IdiTppehDMwAWDuyYOs/jJMCDvJIVX/3QUocBKUa8s+/2aoDQmnHmRy1cRuk2MXFa21TP+
AYwB2hAuqrRerjYY3QReX7HiQsZ370gN0XIYuRA7jnjteeWywWZteQq/0oJeu+c9sG+5XEIO18a1
VMAo9Iv6hT/3PMR23tmLZLkwfUAaXmjzgyUYj+TJL1d5Yrm/Ny1y2YUakzAxG9gEo/tKW1jPTtmX
wpCowSe6e5DeUDuarqFlpsz06QqzkxMN0YdEjJjMpBS4y+JlDYlVHoTZEbsRmirwF60LKKGvCLfT
yiAdvjGSprYvWtKuOmvi0PzydjmecsV7lh0OGeLOYaWPUBSZH5GllhtWmW+3qczPaRFBgfaKcS0X
HukTlkwDG8p6vnaw5A1kyolczcn/NYWHOQcbgZDArDLV9ZZyvBjqIGJEv390J7MHBNiLbP+EPXj1
san7iDDuAlboKPdBiYFTBE1Of/deKx+qROhsbBfN1Gh2R1kmk2NERFAXyyOO6Q9FqhWv9Y2oRdc2
a29RgrAlErgiqSo5T2fSvkyt6nDAWWZyuSlC4DdqcOriVT7Fk5dGnGb3sHtdcmqQuk2zNe8YUolc
hWigRlGRGYF5CR9uDmiHqTOGg9M8/6xshglA1Yb0r1cYf5BBQqNVscecS3OdHFMm3eYzm7GgicWt
YCPZ/uOkmF2WKc+JmNRUG45a9z+DTknrkiJ3OeJ5MBzoXJVk1Q7WQM36fT6vFYN++gU5lcgvbetR
zosQnWKhrZUzA/VkfPGQEKBFwlMFurbSIAEoRR6Qkl5dwxT9mJiZTRJqoHCJ5bEq4kW2CrHV92F+
iLSVv+PK1RL8tAOwF6ThpecvMPy+HZDpfqkaYqBnA6eQKi0OXPCiD/CccnzfZ5xUVIab3l3GjMGK
tY28R8I6I38PR/GiQrIcnIt2k7iLLT44Vw/6/8b3wH4aeKdkDlvaNGKEwFHN/Px0vODiuqMieBqZ
XYB2UBVBduRbYL2by8oP+qaa1dNP8bgVeeyyoqWQX7uqEessYjh+wAzLqbDVKYeJeF8sAmHCAziw
1NFMVBFP0uuQzNovDTw2ndUk3RFYO81oytv1RG8Rv0Xlwjeq1Axel3ccNYtEr8m3CmWDOZ2Uu+8d
MREZVU/GefPjJMwndwQZiIfmMAqKE+VZF05FtTzA6Zk68PUSIeZVsB7mQnd5G8u18S8+C1Rqdigb
MaEjoxnGh7U2nKBSbXEsgz8b9neWeEyMVghchEfqDHWT+RT/5exDPdNc3+QlHAE9NYMf8NlxEgLs
rvo34hnR2+CHcT4MwSFolM1iUMdc+n0ujDutWIAD45ubpQWAfJ2IQUOmcqF4lsURhcHa2QuRXca0
5N4ow7pqVHM+2bIFRQ04ISVwp4PyfH/UKB9F2RCovHLazYBZK+qvIB1QVEV0ozb1kZjRpnXebd5o
eEwuu3gp9VDc0RDm+UKhoM1/ghkqbPo/3hZ7IWsyWfBVD9X1+ObYmks+E0CjbJioOydLcma90Zf6
FW1m8RhQ2Me1EyvefTTViARS8+9F+F83O4LOKdlY9h4C/+9K2WcyrCmCLYVtWMQ6XV7u6/yPOUy/
N155sV8B0uSAvaTMZQBBvnCarfcK+XjtZyiv07ZprPWHjej9QVnibbfw7iLGYZGiNwWcKuV09IhR
7Y5mVwwerkI4F26VvDmDDXNcD8vVTfwjAHeW0NqD5OBLf94IrSoOxbWvihS5sZyeRILurSLLXRmH
6rSM0tPnpa+1JOyZFcalm45j+Oxkq5Yed8iHT5sLvhBuvQMH1oRF109LUu9VBfy7z6wjsgcQe+jv
EBRjuNyx+p4OcX8YPI787rbSHmfyF1er+a78Nj9OeByabE9mMXHvyGpCtpQPyOIrtm75233DnKpF
kPQo3Oh7wJXwcEtRawc9QvdCHJyj+NPly9U/B+EIIJNt7l4HU1CKHk8KcPqX/2uPG3V4Rjl1IdMW
SJmToeEMvniYzf2FVb/JY4ujzoIIyVGUnRq9SPaK0BOHqT4VhkVzLFiuaxZlSVJ22oT380viBPfW
fnLDekE1877pbqXufwjoXuC4lLpYdiFxG5Bv/Lhm9IFNeJXjDZ7ULpTj/Qa8shSDwjwT4VsNqXPp
hQuN07bLd6bobYMxG10vcAMzSEQXlCc2jyX2klT2yt6gKh5DKU/ppssPe0/FQJsPkoKa3kbPA2pT
cji0V3wznKIDQPLlDTTixfVCk52lW/0KkjZBtAxaz+3mU7ryzF9z2aZM60cgYDSzZNfHcEXs/OG7
QNqBbUG/lseAjKLsFLShpwMLzy0o0B00atGsBi2ywwn18f0+urDj+/WfXE7iuC8ZP+2ZJcNhX5Vt
F6SajR8idpV8o7ytaw/oNVdeOBVS/EHSfXzC2mA1nfix8CB0MefPsSWQVToF0MEvhl2ABgrGU3Pm
+nc1lzgt+oWmoDEuE2l0SgNcLYSWcSfI5CQvTp56KEhJo87ZgeRSLQ/Gc/305Ajk+S9V3moT2i01
KRYqFsszGk3akwXbzKGUr9k8f5xLEXCqnQL8mQJ40saWbN9ZCW0UoMgavuQOC4gwOmmpCSgCOSZ6
D9E6xjpYzqbYR/SJgfVxqAFsvTyko4QsIPIg8QfQ8IKVquXZby2k5a5C6bY4OBg7cxDoSnnJQVJ5
aquXTm2rPyek/m+1ueGixFRiPyCpIfAaxKSZt1DoEwJs//jfAfFuB3lTDDTkTNr5GlZZdyccD7Rz
BwMelcZyOoQUWvYVTDj9c/jjkOz7wJyOR8cnAKrHQQx+CIdFAbeaFeicV2p450sUa2Zs4cwxmBTw
K/VBPUFe3KBRF/wGMD8pRa9uk/7vcPTvrCA08kut1zd8gKwTjoCIPKfqxjRsDyCBqe+VbQ9zKFCr
I/ufFf3rpwuuUxKXnjLJ8qeYl8ENTkeP5eS13BQO+QQ2Xgb3Ekt2NpnfzQQG9MHfxL3tnUUPbhNl
fnUDoLT6KUXHRfKmjLdBdpoErzz9fplUJn9PG+ddX6qMWsbi6qHdcOzxfoUd5jrqQl4ebSx0Qs6b
v0MASG3CHThbhUqGr6OBRvwbFU5yKiR5qNC9g/MfIBaroK6Wril27DikUNNiavihc4EPeTvwTUq2
1RxtWqCDf8gWEzcYIYWjGZRBaewO0irdefaKFdOJwpwtRGY5bMR7iMZLZ2ArY2cnveYlZIW7W5PU
o/TalLIOj8RLuwanU4CXMcXDuSEzcrz3dLWJKBr7XczuX8voKw9/yZJPAVJPPITePP/Z9A4Nwhgx
+xycMxdeiSzItG1pDEY753HD+/HCW7hnrXrbyHV74pHEgTTBSInkbVi+dy8srGleaLS4URv5Dnh6
ZUP8xWHiNvYf9P1o+kCRwfp+IXw5iCWej4nmHphPh0By1Fw5hsDqtRoHCFdavxBGm5c715tHcZYb
JbxJfTfiCK43i3SgG3HewUsHoBkk+VEuf4lDyOse7/a4fErJqFB2YY5tBmm4fUrv/e7++n7c9nXy
EFYWFxPKfxuN8BWz+1s7coNOPe3VF6FNO9AVrSQDo7wOnvNIurAG40S9C1YATQJIh+oOfwrmcuQ1
SljrxqzbnCBR4hlRGg/mJVehdj0Gfr/ykX4bTpTby526AgUQHCvQiP53YJ6buZv/tRfmoerOaz3K
gTZiZfO+OhGRA50EBkJV8QHRjvC4LqL7rISt47a6i5tG8AZVraPiPjqcsenwNuv+dDlt3fEbOmIc
3QyLuv408a7TPWwgE0haQyGcyIobZlHSuHEnVD459X26ipdAcYAawZCC9bhR50aRFDQMxJ+ZN+pt
+Nvh+nAjBSIi6B3gI/NBgk9PX1gP1pLJQA9jXZ6vM1dikoSpNXPSvtqOlRKQAnnCAZkeWMR7ZMpq
b0YBt03D+hAjkl3W/a19zL812YNv2UbaYRvGhP/8AX0DELHr2WccIzoEhQ1fXGCBRmlIa4S9sbTB
StwBbHHXlm0iVT1HwDuooTIDX9nstNAYc8DeNpOisqzkS7Ty0crtMfhWj2Ce5a2e3947mIWxnLLB
EDzR5pXLvzYkTVQ9V+O8DiyLrPM3XxIseNF/+qlvqmHE5rtfiNb2EhB10kTmzOwhYledGUYHl8ku
pngdRcVVxrKOMps+4uPoGzqHmVOAZweM6XgHwj7zsa8O1Jlh72eLHl0eaXKN6GzIid9aiWd+Za2Z
jKd2BgfeWOaMT2u4go+8+enjxhCBv7QvUVbZXzEdNHfL3aBd7EwBfQROFn9cyZ4zn1oK1HwVUe/m
Iph9AtfH9roeYEvnmIEKaY+l2gSWigzX2A2L2WlYUe0OIdT5TuOEUhB0yoYmUSrL2WSDXcTu5hqs
NUnfKjTlt1bWrUgvlcICP+L52f+bX1zcPSY/J/IZ5Tu6ErFvpoR85P14kom7JXxXGb1Xlt2+cVOX
0VqIj1Q2/R71UNlncexBFNSE1X7RWh0msOHIgTi/944Js+Bij3FXu981oeU7VvjETp52v3MowEVd
UVV83ikTnAj+3zSG60jp5ZZ29ZIh7OLYh/h8JGWN+qUwJDUklMuAWJ88OwnfyZEyJqiwNHgCLu6S
vwbjrfmWXg980fCziyfkKCVqNbtLGoIsL+1zLVEp5sPkDp3/VL52QYmfKlHum+ajLLjCq9pmqXWh
GOcA8EnAzJHnRqzV1w/i8HSGpeKZ8DsqwYFGYIqf3Fah44HwbTNiFCxfQMKHpwRjIZQZXhKmkOpC
nJN7mOroSWUaqeqS2kk2EbkBiSzgA3GzAS+kisfHphKWY3krKxHgyzUNKOmIi736opS0Tp5BNTYb
c6hovUwNK5L0cUxDvKjBDTknMQ1o86qgfer2gQJ8iU5odFRR6UTmBPIzXP6qE7A3JRvtQ1sGwNBx
U1wzjvzhJKoLDGW1eHLpkHswdFGtICQaGnYMbNMV0a6b9CTvy44sbGaItMAzS63kzCk25j7hfdeJ
+OPUqR6yUmHb6wDsIfJhc9cIdvlHHbU+5JiXOBOx9UyFfrsG6dxUbMgZbOO8+hHscXD1+qcqmnKj
wjKq4ijzyYvMGZI7qWq3oO25PPWbJFxYmZH4sDl7Uq/DKmOsOMEoIRseYGSDyOREWjf77wUzx9r9
lTq0odQhgVbI6a6LqP9golPXyXfPYicBFy+lD87osZMU11YJTgAI3lltKUuCv2wSDib3Wl+6bO0U
yLL1womc5MjPMnt7KfNPu0F6FxP3/nI0covUklr5bc5LqTzWCQiMTWoOl5LRjVpSZgtCNoryGU1E
YvSG+IgwgwfTkRK5EuAnjMxC71U3SsYrqRjw6HAB9UYn9KcXeG6eZZM6g5j8Uo9RxN+t0axGxqcg
4RLoKZ4htacSnsBYA2tVbMSF1HwXPNZ+wu37g0WgF+BeJe7Bv+rbMBrIrZxHohobGYyAE0qju+mt
LHGuu33SC4gOCnYl6Dl4k1mxP9qHji9AQebSTHji+rKGo/ZKQGBBO+w0PgK6aPYcg+xHiBONHWNN
QeQeod8in0vIRtd4SMlN6MN2f9S8AY6kHmqPu05qgRvtJc3Ic2HunfjWun4RpqlMRXt0xljNlpiD
AP5KZBvXmfgMj0yKbFMIfoCrQVroYZnmJSioW/pQ3wqCMrgLWt8JVWeegr+29sB0Nf946RcouKpD
KhiCL3p3z6tYX4R8S8vI74WdvAO4YmZwk4Zn+2qYdmCvhAgNjpzZbMPztkeEtxZA2KkcxeUfjRAJ
6oc05WIZbIbAvtxrM3o78uUC/9+hhJJIHvOGdWD6DetJNiE+R1uMLBeQi+LzwwTPVoUF+BGFEf9n
/0K1jTU3UNLxmF/cGPiOaXZDSqwNQSsZY6BLqLruDc6yVAZ9FF5mXXJ/RMgom80rYw1YASdyxL7X
v9NC6XYCx+1yVmlCXcdVjOB3C/o+M6ke87qEBOl61Jw5a6nf2PUTTLgMdV1hBWl6+SJKWGjQtyIj
7IDuMbj05rE95PO7ZbU/EShqYWdhU/EknVadH+Y6+B0XAvov9gqdIYYWKagtmXo/6M7WdhYiXwV9
/Tv/l9cLxroSWnXynyzF4j2NwW+d6lpY/xuTXLKZPHUXACT6q/2RLQmQU7o96MZ722sY97s+aNPz
KTi4mpHoDDUlVEPOgpPRHfDs7Dr+5cEis5MsPovHog+cojwg4257GnbdW4Z4eC/dGLbE9asgIK2n
qwLU0PT/B5yaqKztBh7ByAXu3oJ7ttmrOUp/AP4c0+JTfVxJA4O2NbstVN5aYKYJznfvFNjuKkWL
1OaMTbCW7x2wDsNjJ/hYZv8E1nehuZC2pr+HMMR+tlXGnzVWm2go5FO2o5S7mJNLdZEhhHdc295i
/EMqDRzKzT4sCuxCjtlG6dWNUvdQzNvdpT2UbQgBat2EeTSiDB3pdfrKzrF1nIVHUZfzkeUmFVD8
97PCGWz4ak3+7e/d2ZfjpygszJoNYeoBjTiRfQCM8mE77e7WaaKFI8+zh3/kuxnIV2zV1RUiVgbl
CsSAsMuuhsKjIV/elR9BiVfSUEjNxTsYDB0scyeVA52tgoWu2kpk5WbA3RgjCbNHnGobJ4bwDkX7
7zYr541sXQz1Bnc/CddTjMfkgWeaVG57DDgBwotCyIhlrRkm8hpNuBL6hkYYTCCqbZn+j2q4KGWp
qDh6b1uMjAtb7KJrUEM/fwBrzREVjiMVEID2aKGSbrw7n4ZXW3ANXnR9EQwFGBuNvAoiDOWh4FjM
H8YyCHFxf/KjDzlTdj3TaEXG3p0WyCExOyGwCG9UHnrsgzd9D3m8BJxmeVrAV0c1pffNJB0wrWGp
Lx1EMctSdmFBpU95BuooiNHc+fbzAwMV4+osHH2L5gA6pJ+AdTBOXR8HC/qxSNnJN1pBgZzmuJwV
hI8rjE/vtHFn529vp17Odu5R3nDoDuD2FtfWzUe3M+AOiL2P0hSCyC2Mbu0WnlVLGxkx7fRCu2wb
ceQ+Gyt/OcGusurpixG/GinGjrD6Q3KIN/mKbluuugnf0Y93VEnuDepEnK1B5MCxA5e76PXUkRLZ
ab4aDpUNKvz3MDzWCkzimVU/byLVIlTcHf2hcLyTImmzTlLPcoE7bEphAT96kZcoSPT/aOWWcYIP
Ij1jUkY85TaSx0z7Qq1j8vAwCeGiEjqHdajfb3BeXmty+vq05PO9DoM5k5Qd4Ir3nVxDDr2ubnYi
7JMv8rTNP2Pnbq+PTq/zv4Q1aHchRlQePy6LcvbqTr5dKxzt54e/E0RPqqDXEMeLt8DhbtcEnk0m
QFmTT3E8gWi6OZi8NBCw0vbW4lxB82/5/56SM56104gjmc/qIsGJpOt69BohyfzyynOzNlFcFzKB
A8Nayu/wuoABdfKTTdPpVuY4n+ANNchk/ENroaujqYKKsmJLYL+YP8vYPlFAeq7kiKnDkGEvy8cE
QOMk0esI94/5CApb8hp1Jd7et/stPvHy/ldNec7PWFzI3hMCDmu1Fw8kkcbOVIlMHDHegyKr4YLs
a7D8A+2Pgt24wqlqVajmwVsWtYGm5lyjn7dldfog2RGQmK+uc0wrzEpEnfB/t6jQBUsPRFH7tFPa
fS4nca1+wjZcxaf376lFjeZOmjt/CBCPVMydtmbIS/BfC1wy19jmgWZ+Jvjc2GjbJXjEz0+eV6+v
swCixwzHFnmWrbLj5FQBg/GuDcGYZcDw7bfj7mCxwNKqXGnPBIAwluRcVASkVO73NiQJBcdTKpwv
/+5TGEGjVRpVMZABZZf/8bqzhG0+p8Tuk7JIwrhpsPZIkwcrXeuVq9mA6DewhUdPwpmZ0fm5+Dxw
BvuovSKQGxZ/VXqSMk0hZjd2Cl8XXofYgrtb8uP2eWp8mJ4HhYmt4CxSz9gZhyBX6Wcf9edWCv5s
7rXdG2WvAb6oTJ+myf+6Ik86HSL2obgqy7tSePruXrQRz/x/bCn1Lv4ddOV7aBhIhkOqrqVDX7Ok
mWznuvF5zOfDrwzD/IfpKXwLYuKb7PsYdYqPwJRBMqhUq0do4Rc/7l6UUOXjRaUEr1UXcSLVlnd+
M5ciR+V3OVkW7RTegBsvp+TX5OHCy9SYhYP+gbn132OzxUtZMqV9LVDAZm6cnjIMPztWIXbRuzRQ
5TPQdhV5Dt8nh2R5tBh6iLGe3rAr5sr980Ps0cUi8rqHwl/V6fl9fMZJPvJo9G0Fl9DnKBXBJfC7
+riEqH/EpMKmo3hbOmnhxUY3bBMB1Uqzwe6tVIn88iWAGORaaonbFOV4oG3L1yLtbIKVSd+Qydwh
+H1xc1k6huPzLumuVQ5VeCZbY1wSa4J422QbhWZuln6p0lrrdHJdC0kaFGrDwhUW3uj7cqhuEV6/
IDJDD2n6bzAkW2soTrrPaGnmRwwalmcLX03+yvoEENJD/igJCOFIPdMnnCiPDqCa7Fqcp1dW+Iog
pIwpiPkWhIxZ6HKYiakZ3Tx/PbjV/4ZtAcQUh4x/1lCrwcCDOGgBkS1yd+vwzfMBsdkUIaYH7jpf
6i56AduWXYtvt26HmJ770CJwcVpDM31APIBz4+2y6vxwJe83w1Uc6j4D58ZHE5NWCQT/39Yt8/s/
rhHq6rTsUIQnFHjpR539+PhdNzYErR8eaVx2RDYP8LFAY+HqoVQmOqnACSN0jxLrTYJSt9eIz6d/
9BwZ3Jf1Bayq2mPGpKdNM+y8heAxA8gbvdI6VDn5Qh6N1FSed54JyDr/F3+C93VIk+H01ZPX4BED
d0UtSQxdD3flpLmWbZcXHGdMoxymAlwZ7UtEjsnCpN0yEpErQrOCBMa4E7q/HhPxkpHu5H/ABzEK
6tM7teMWO6v5bxxd+QUQp2UmOD8+CU9cYTg8FaKbzl6Nkyv+Ug6moEQ/7kNnQ8XRkiYHwAAMVW+E
MrOfPX6/yMEQLODzQCkJfo1hBxjiCx8qM8j1QI2JKxyn89YCk6BOfJIxEGqfiMFoyqjzZwwqkP3g
FYVQ/4jxHvwVw7V7hZgSLarRxDpZExTGSNCt7eAFdCksuFofIj3y0rGllsSXAQThOGRYkaurtt0z
xw9uMQ4Hlqb0fb4qQuQMZtSXdmNb68BA/tufGft+2VkrgfT3/CnxtIYl9WgftY3vhA80EB3NMOhd
LXtrCI8B/Kp+E8ez6cIBYBEk19E1PgXUPlBdYqcYPpDd9yG8X6azFfw5xEKqbboO7KjG1f3KXd0i
wkJyOOYbRXL9dBTUh8f7dYJGKC+DNZj6f41njhLtMdgB573pi5kQ+RAsP5uINIKfc8t9Eu4sRCxG
OvN8+n1krIZCplOb1vm/kf6ib7PiElnzjb6tQaxRvxKjrt4caU8ZHh/rtPpb2oruvL5Zs9LTCEYO
aJ7lrgTDPBD/q0TYflqDjKO6Q2QXQnlQEva+ShgsCpcjOzhnk0zWayd+099n3TvkO5WIqAAlS+22
a1GlEIuGtMvIQKN+eDMxaGMVosnxKR/IyYW4X/b/xb6fEKdQg54384pPOgHgTDVYsOZAr80Zaa27
EI7BxVuqQ623aMxrdUImSaKw57oWZ6qz36fbgykKjCsCteBKng+jKSltoKOsFGZ3y3KpSxbSNKPf
ybMVVvZFtBQJdFuc7hvUOvSo4Pjd9fMIvZO5ZrRZHeLwrTM5b1HxqbuBevUsBGE5Z7tbCddZeY2v
mjinoJyGpKb19F01idVayl+24cJEFJM5lmNo3RPe+N7niqFghkmWQde6BPVJcCOzx5mKjDXATI+G
zu18rbuleVvUr5URFX+bLg76xTkDI+FzFNexnyxFQJMPMAiJt5BUNA6dWGdZ9N2xrFoAIXCXFoiQ
x6AoxdCIsB4j0QPJcWVEkgUdnWG0ciY9MbNULRj1iIu9JMQj3t07ANFHb1FdLnS8GSDf/SDUVINA
sqNNv/hGuKREPHU223RRcPcMjKQDf5bBQ9j2jfm9Qw/aa4Vp8wRMSiWFj3VnTUpaVtkYB77Oib3U
2796IlDZJl9/yrS8mCsbs9875PhH4wRi8cP3DfsEisNDHYMc4ywa7PI7aREo3rzRApI9/59iBXy/
HNELxk5YwNd1kpAnbRrVBVGRwViIFGIbcGyxFtuoXNegeLTYGr0Y5mRcabDBalJpyRxMWD1wgcdr
7seXTo49UTAu3LHKrCyToj6HkvSY2MqsTLEgBO/qN36sCTxxI36ewZ5lt5zXt3Iiv9fY+9PcV6W3
e18WwFish1vdS9rAr52jp/Su/ZZmkovCWpi4trjJtRONFjVz4ByV1lNiLUJLp0g6oWrE3D6JfUlo
wewjk3apDr94f3lRnsvxyFe56OwqI3pY5YZ+aeZbaXTfze9ir24+x78p4zVOXO6Dn5tytaFfoSpg
R5rIxcCWCZpDtwg6Dv2sC1EUNbuAq4XaGeutrpO1QfCxA/UkkT2z+5nE3RyQCeAHSEFMoxAom9jt
OTr3fgAKpyR+GiiKy0ihHU8t1H/+cZq96bjgI9XFQQJuhBwffJqc3IODUYu5gSAlB/S19c5jIlxE
uxKX90wyDEAONTR66PNuG9+U551DyA7G6o06GVIZq0obzv7LTNJtNna7xBCad1RRzJ4uIsgF5d4h
Pxn+I7gmQ0MR1EBH1nMN+hsoaOJY7LVhr1d8BRhRQvu3z5TB+5uVXr6GawLlXWJKdtXxTPhlwVNf
evFKdOZVA7GZR9SGVQKyw0jpQuPCeoB0HlF9czbnKny+DH9+kgcwqD+0pTjKoOypv6kJrAQMzEas
Qxmp/ptPE7icBR9JnUGgGHKciOthSlyOqVDYe/sl95e6XkHX/hGg+2clAYTsTtCtEVuMUTsM7UAW
aMjXYay4Y6aNvaqVTJR9+Yagjt4usYn8AapvV4BjnySTbRudaeGJOspIlKoOyv8pySzEX9aEgKqI
wy4lra75TFwpCfHI0/HMPtGGKud+NI8P5gDYMZcIWsVQN6KmN6sIjtLryX66K2XG+a6D14G7Wi+b
Rz4ZSj6BH82+vapDQGdm5F8hFTXclNUSg3ss4ZTQg6dOzeRrrP3D+IRDZzZ3gT0+R+3Aiuxf8GkZ
Ss2tnfrIXtUgutyG7HRIAhLOtFYFMfCWu8xz7eKiDgSgno2COogdGnmgv//JHLAZ94Ld4KC4djf6
YJ5NueZXK8jMBJPwzx8W4wGt+/xhObf3y74Se4Zn9xiMH1yoyeiNG+dS8v4aTo4slVqOmE1npIiM
rcx/FVGqXIfa4nX87y1eDfFKD/HmHow2KmkPppTGyQCB+y7tQA7SKGYkcrww/PujoafI5/Ht9HFV
pw1k45kB7XjSb4rZIG3Mvuawlc3ZvXYiwgfdKMmPjB1dIBl+6UDy+f2ZFIXBqG+uCzdA8cPOH4Cj
BDN4CEgUakf1fFL7+0dq+rXwCwWNCFGSfS1U7VpXOgZ7J27HQnkN/vVmMg3uMxIlybB8x4cSFyI6
Wofe17NzG1ee6blJje8OaiJ0lnTQqDfIwYpskHVBE83hhixw341OB/DJr5G4SubQIOILp5z+jUY7
x9OKZHyaBAgyRa1w/F972e9SQirIYr8lKO26l+10eeKiyRcZjGWEUbDAgCF1xFCPqLJ2gRcvGenL
mXG/vHNS2XbI4xAZe5BMGsY6uvJHIzhi8Z+VYCuFfFPghp0rSjSCMSbLOacGNFiCDD2QiwDswugP
ODK7I1rHD6rawKPNsLzjd+Ow5/ccb7KLfKEnDjRHVlgHvAfZxeL2bYFlwxPKEo98PWZSWv5CINUN
uU6/dPdI418ncodFyIt+lQ+20a8sQOXqbzUQkIFN9epsMb4QkUPsxWwpLfcrYLLW7Ocd0Jg+ooTN
Le1U+ZCczYgKiZckvTGluISe5IdIra+uEB6u2RGrrK5vH0cQTP6DR8E+NbqX4ZT/l/fux+BoyeYc
8WUsb28J56eAFhbS2qGHoV/OLMOAGqm/R9N5qqxIQDpNWWiwP26cpj74YlxkRqnwFd2fVm55MjwV
JweLBfmuDY0vxpuxhpms9pjboiw68aQZyaV4JK6rlNO+/hd/SH1U2vpE2l/zYarb2oIRFos4CtDm
Pd6kmQsVRTA6L1tJn/6BViw0/IxAGw9ZJfm5GsjJrTlDrtxPopGPoLvoBe5n9h6yD5MKf7r8VEgd
//rzWv9OKTvDx9PokboCRsZcY8J5ZiHsqbvn1vUAJpuNY4P/paXfPylSGnGPcnlKRLrifElth1vD
ajVDRwpWncCdt+T6L3EnROSHv8s8Z+QkG6yURalk1RnnVQ6Kc0TkL2yv3CZHQ1nlPxivSGjbgCht
5Fx8W14ESdA6Ks3CsBpiqJCurhvLiEdHp8raccgOGtw+v/sVihr0lHYPfXKtZAY7Too6QDEgE3cR
WHN82e8Y0pBy5c9lIuLAcKkhRP3/5IQSFfUrWYwCpbcxbJnhvMjayucGqyRWcEUUYioIQuU8SI4G
Td+B1u17s9GDur1It4uPJICuLXkNpFbvTD0gmnxiTARBLXJkeX61A4p2o+dikyEJYYw6ap1k1R+l
d41v+4lmeGXiNOgPDGSu/jv/DB6b6Yh+G0qk0B3ik9UfyDtBeLWLboffgUDbf7bzCWcKNqHUsJPc
MHSXX5ccBIxEqA31vg7kFreiPMbGuawhq4b7X40wksnhUKvW9AgaU/Ao45/66erIgOVn8qMGi971
eFxy+istMMEFGoN1R3sQKMfGNLFhpRRJf483ddVrYF+G0aclhEaH3obKfds/lON9b//1zpmkVlcz
g+Ww5ee2D226JyMBjNbRHWb/U+X0ZtAEKUaaps4M2EfZrOO9Tw4nth5E8Cs/TPuXY/EIT+df8F4S
80qiHvKyeucJlS1FNT1KLZrT4C9yftl5LgRCrPBn4glvd4zyjYYfrz7RNTu+mg1bjHbTf0nXXDjS
zf4v+vUIuMx7NChXUs7j/x6mmDecQYz0Mhxme56IcsBAtPVPLdzlUxKfYJo2SkWXIPu26gCvPyIf
PJnjqK7YGO7EEt5W1vkx/ch+97nU/5pWoc6TZ4qG3C1LeAjExoTLE3rL0RzKUHSHsJbP57D8cyxH
b1Up4E4/4xTXbQCIL9TgT6oGKDKHFdlvdpKzD5A8IhVjBg7MW3f9j5Byb5VQGowcIcEXt3zG0kLR
eXtDwTYDRrSYMYi414xSwjBbWbOZ+f4ymYYyrsKx1hxPYcyT8Ei9CoBwivl+pEE5hZ9bwgB/MfpU
IBr8iMux+wuJIwZQ9iMd6il3lJ00FyZV2ZGWcTsGaDXq/VnGx6GZc/sHHuUMAxHgevhMv34+e3X2
IeCHuNI9VbxXlNcRqDNc4ro7CyY/CUcGhXrBX+YaR7IIfYZ8yLREvrMXDc2Bo/SHpD2xF3KOe0n9
xbzYpo1xeVhYdFdrhlBV8xGzXh8FTBO+IN/6RSKldECEWzWLHgHtsGpyCnyrBFy3gpRsbQNRj1tV
11FoUH9OvR2v3f4naZ1Vf07Bm0DLOscdITiBU/SX4z/a5FEwn+LKy7XMOrx6ex5EjYgp/Q4onx6b
ShBbWWBkZYLu7vYxiOfs+e7oWvLsDTe9jq+LyMgz9F/jUHaywn50UZmx+BrAJE8Bp5AcrhX9nYrC
A0ey/HRqduUdbQdnXFoqUP4df9pQUnjP+bqXQtPElnj/IpkVA57OiAW7A/s24ZvYRyFgSOvdN2WR
3l2apZ4PfLps/+zspxxw+1+C11tPjfKocVfNnUVYfi6KjOsMxFsL+R+XDbkfY/WVOg6oUQtaLu6o
h+wmL8jc763H+i7bhpkFqd2JXMMOOdmccA24MpbPqiLFWaIFC8DIHm5n1gsGz5fVwVBO1yygVUVn
hKHw6lh871H6HMkEVE2M6olm0abRPEjqzaso6I5bxrDN2ahJv+hiF5IZKDKHUcfNmsrXJ/nWzjQN
xG4nDYIULS8SOyh59N/e1jAclV9b/UflnvhCUQad8fzuY+H/xU+CiQTZ7cDQxLoF/07RVnUl711T
CjzXgH9BU7H9uKYAfcXLnVzWjIPcyIcOPchOAT5yqkElOOgUXXBZ+CZpKejaSRnS/2lBUlQ15RZN
5i12qzaI+XPD+NRoNc3iqKlZUhkDPhUfx11ZifIy2ZwrFoSC8KhMEHxZIPfqPDeufeUcQ60GkwAL
GZD0s0XOW1cPGw/rM2Kiot+8rYokTh5kyji/kku3QV19pQNOCfuKtm+HcDhVHfPdqTe4DnZq18+i
o21g/6vyhppaCLm+28cQk/TZX1xrx2waN8t5t+7V3gU5Ja1onqlbm4YC+b7wrBnuDGPOoY4tQHyl
aJx/li9L4L2MAj5bZfKW6TLxDUhdTH2C6etHfkGrDx96Ahe3TNxnkZKavvqDgpJU63dPjnwpI0I2
t1u9QdVEX1wSNriskafuPUxjNZjNwuSZSVfYmfZ4cwL7uNu2kkvrDn3P8lpvI3UUVJ9PWNuiLMiE
X+K6/02tAOX3wdMegTlV0jmYyHNLopDT3XBMymAqVqYYIFKjXbUaH9aO62tlQ/mkxMaYaiUmEzRg
ArHG2QjH+9u/fg5HZbbUVruCk2UN+9Ppms6n3Y9W6FtXM0OTzm3izBW8opPBrjQflngV7fz8788u
t9AB1QWqHHb8bgooiJ6OCj6xh2PR880AThAV09W0UTCZNY+SBhXYVNkTKoy0EO5rvLqSdzdXMtR8
oTCOEsaxZSbFcYDSNxjL1JpzhgdnEQwm90gHltqf+NrPiVpY8WRu7c6kiSIul21w32SqB0sTa/E6
2s71QkixDRLDZOhPrUNU0FHXVAlJmlsToLpNt16ZsiTUH6DfA+KgwgFiT1sMvgEPIw0gKBleOANn
HTFu+qIL8FUaRKCl2Gx2/gsOgZr3SyPkjnQUKg0R6CHIRGwbl+r/ES2WJ4El/v9S477sjHmZao0Q
ithVCJSVZI3KDV56a/8ezCbOCuoqWVkQ9k/nbuuBr5VEf2JS+xkPjNdo0R7YUp36Y7mrz1gSyd9A
Du55RyUaR1BnpjgKLGrxb5Pl+qiISRMB1UsCtNKhNpCvMMoJ0BZYK5UslztfFX+wckZ2BUwG0w/i
lXd0E8ucG9dply/Lct73hc+83S1JGPIkU3+myvHfHsdqcJPK3yIWgHC4s+BOPpsBWQXti4AslWvl
1olhBodJm6AaIQd4bUJcOW/yXTeQQqr7SVYda2ryshr6M7LVPPJFc1mcm6dKWL/wsKf01s4q2xc+
zdpp3T4Kv9b47tKmdOsGjc03DKMK0UsPTunPh0bvFrsgDt/5vyuZy9Gwn3zYQLHU8hFr8x+5/kRM
Cy1DR9QRBZrPhpSZmKGGPkPcd67NipjcBCnNYGr2upJlKWx4ARyG5yg5NF+v/eJK0xLfD5gYbfDT
1RzwkRf6iYd7snhlWrkIl+Edb1IwtScj3vBrxmE4JGmcOfvmPGADSHqsHMEUtyrDA8Uc7OV7L9W8
vjKFPd6XeVSCh50KR/334wOOCbiDfKK/ZVx+WDy2U91GuhnNgaYGVKQkQ9kjRaZSelmUTnS+FC81
zL9+VmPsRY0PmJb7tOviWIUP9QgaAoJafaAL9lklc3qAR2SLJUd5sKnozR7Uu/gcF7iZJUmp+3Iw
d4ORtO1Vd4HnJ3NLqSITH/xsoZxZ38dA3up2CpFdxNVVqF+NiWi1zRZvUz1VJGEJFwr2tErJZSvD
k/wSF77WWIP8gNezUNjxnGPfM96h2vqgTMLMbTPdiGDN0jI5urntT5pW2eyI2yECUlz8azZhP2nN
DDT5Dpujz3aRC7gOQlBDK0lGv9jekEmSk0blPO12/sPCl8x9PccSaF9ysj0KfxQH15dPCWOtoajC
7X4w0on14tx15TOsRXz+bO/SrcX7/8UiZBxeuRlqAz/f2FYLRBO7Rq3aabjK0g+6UqCEYGBkJSgX
9nlCuWcXgoqFlobnyVpcSvtmX0fS8l7oc5iHhzHhnmIK2eW/1yc3OgUhsIZoK8gII+x5uWZJOiWf
7D0JTs8jRDINnVj30LlSDTLLysSTCo0JVWnLGNF0QfQecs71yqZdyuW6eU7MW6PJaawNIUjsxdon
kjNVReYAPdGPgzd4KGyKhSYa5sKQLA2Y4axgGT3UWl0qw0+k5LBZo16AIm6DDqLDSsfaQP1Fh20o
kk9wsbxd80IN++nenPhR2K03LEeMtbrD0bKLsICfAkypJv/TlBRxrm0crM/tqf54Qcg+bHHjIXJt
/guB/E+bEATCSn7zF0gasz3nnCYfIEhs0NocLYl+xTpYqRILTv6vklvfvIk3O+VQxh2usC2ToEaD
BCrT/ntqjKZabgdblhKbNqvSo4JOYMD9AjTS59RuX/GS0OnVsP2+JHzQRtLTJ2eHcdNkSoQj9UJr
Ka38U+x3LNAbYM+P10j4QlvneSADcs9PBnWJtyaZdeN47xMfb7X829p6+mbaMLH0POcVbIihmqmG
4PTPbYM9O3hl0/JlGsbWeBMeBqWqh2Y3ShleVS3yDsOf2yidAVNhS0srALRTSM5XJ8C8xHatIu7T
Uyb1zrQCMsug50rRnmVzbABYLzROmH7UvZS8yK9ssBcZfOd6wXWLVEGHO0wUk47seTl1FhvOv1S7
yYooaq44WNNiG4Aohs2DxzaxWH7D2i5L3YiEvXsbpaa+CUToZBfgxpy+xk/RtIYZlQR+T+/21Ne3
nuzrOzPnatVA1rgEp9521GovvvFQulM0pwwL5eKvYSGOmSW1ZaZgAKFVhYGs4LKdfQJPThnbpxeW
4MJ3MposkETsUzEmEKQRDLUmLnmGTUx6Tm3PTC3mwbwRALyKnh5N/ORnsKL3GjIcUx+vyqWtFx+V
SQ7SRwKbnD2gxCzYBwl9nss9BpSSGP5BMV1zx4xhzDlPRCEn0gSeYVq7gvoQmKHAJSyx/Bi5HZgf
XMI4y3FrouYUzb0JoK5s40q/kMsvBvefJZwEKmyT8pPAw2RFffarHbEjsRmuL9nLuIJJrvdpAVTB
0CVGwDEfxYapToSQQvzWroor9EoYz7o3TdVzhP/Jx7Lr11y5AmawoavP548FALP24g19NsfkMJ5+
cPkAP930nJl9I2kYFTRDWFxwfPhXmpK6PUJM33UFVhE76jSpCoc8mX/iPR3QDOIXJ5P4UWZjqiCX
tUDF2u/nbpBllmMxZKdfmpuNAFkpULHgjbjIlFmi9EYTFiN6qk3Xb0q0C5+zmPc2XaR2zA9hUGtk
bxOi38LUU93A9MhrE9hW5T5ejHHDGgduNjzer5+u6KgXmf1TChLP9aBugg/IoBEgMqOa0M34aMjK
EKUlEVZ0lwqZkYGqpVKns9Zm+Sb48y1x/wLnyfWogNzVbIvkzl+R1RKv52N3JG7dFRgcZ9qG3OL8
NYDmEnuqrai6sQnO/HXyou5sIfqbTTektjp6cyn/NZ/oggFTW0GaKIgvlyqKIcbKjcAwhGCXVw4F
GxFGzIsZaZANE6Uj37Buy/AK7xDjVOS6xA0nZf+Z8CcAW7BmB/4Dm5wsV5z+CHbwJx5h7sMFVsNi
4wOXZf7t5o8zOLwvG9VdiISwoT4yAOZesfCG2tgUEvx1A3ZmW/87tfADWwWnKolRAvlAdcwCPIgA
FVKDCqkuxtQVxRhkye8EHwtLTdBihwuTrC/XTvbKyi+p9wnZztbMyYuexP9dYRF0ziCqVR/Tzagh
ZITwGIPX+cwaFmOGFutZkJmfDbpYpJN+LagfjTwU3Pw49eCB4PyhXfXlTcUBTWF49brY5ytIuzVv
S7GAadlOa1Q9xNl0CVp+p+kwHydmYW7Cvh2fZu3VcCrKnjdf89dwn3YWB9PM2QQYVB45bLKp/nzl
dtLkvsGSU2YOo/CTjmotqSzNX53AKIKATsw14WlwJyL1/HUk/YVWqDEIsuv3epjwcT84XT3jN87u
c3a1S89BthHtJ83wY8PF+wkTsKBv3guuxPrn9f8NJHTGFEP0gM3HPprCf+P6/SdY6vgjjVUaTBS8
C3uV4u1RlnzaKh4HsPmUekA6VhcGy92gcgpZQ97sWBsH8orIoBAJXgQyXEggDmbgL2nIHJe1C3uv
1PwHkhonDOmX2rOSNAOv62LM5IghzB1qKfzFrIkMp1uu4eY82xosoNh4gQ48PrJo3h7JHPD4uiYJ
Mb1QzPIB9X4momxaKV8Ojivu14cInMWRdc/qPty7QF2wUpXWweB/vxE4ufmIUuOFXoKAvgrCU8X1
cAcuqTmm5gJ/GgUjvdEo31qfyjn6pM9daQirGgx0IqRsYKdUO+NhevbmWmuHVS85cMloEGJcyBWd
aKaKvRmolfCuSnHW0FbaZ6NYC6z0EXynlXwECO0FkI0bfSA/Teumh4nnJJk9tgcgBjlK33OfjfOT
ZgQlOcrQcbN5CSi0B2021iSm2ZeHgYBK9LXRZWvKvTKkBHQ72DcFJl5Od4IyR06HlVm1JpWtgNlS
FyJr0FdoRotVfEs5jHhNTcMtC0dQVdyz3ARcPa6mkeqEax/PmRsYr9+g2T5zokbtmXF74Ux3lC9p
HmvfuyDHqRKQ6Rx+DXyrxCRRTdHrT9sh6Ka+lrpFpZTTOo6puRoVJjs0IJLVxg4bRdrJ8eIe9Dqo
UgzkoasKCmuRiU/yH96Sh229ZOfNTcy/HR+bTh7TOE4mz/Rlt/7xKBIBAjSe7jK0dPAMltazrIXo
92cTelNLmpTdRu0lZMJYRNP/XqirVD0kx6Ii8Wj54dTS4RNLMjL6EBBCOSV5/UhIsaxCW6hwVjll
tj1z7IcA5YxDIGmAbX0ZtN6vC0HNZn9m5AOlBSfMrOTVz5UM7V9fQsaOxNrBDlGyaWFTzCCyv0xK
2DLHuzxXYyknJ3R3lOm49l5NmyxXOPMwrcICVAKmvna1qHMqrpyaMASvLDEOxbQNkIKGBJA3kYEd
UJFv25QBUppi+Zt5sTMSNnErnoTreDvvHKsLM0rYIk/WFOhi7yIf0Wzkw+Ssh2aFcGuHnN6NNw5V
+yS1DiKU25DbsWQyplW9nh4a3DAXwnheGByHw6wXDU78n05flBbvEfrIZAIcSpKXtiNXw1WXDgl5
NIHXRoDvUu9+f0Q6JFcNZXNom5+T2Lj818Et2ggoA5TwYJ+7dDjIPw+OKMDP4PlprCQ+0/HUWEO4
OeVj03Yw6+8NU8cF/9Be0Iwt2X+3CPbEf9mB0dlz70sAEVQZ7kpd500GjCPCyE3eL89Yan/wCRGR
JrmBE45rRgw5mA+yA1h/NXtigPKVG8C1y05WtaeI/UENMlPONw/Ol/gpcPnyeZqsB2i0DqiiLYBR
D4GpXTm2nmwKesiN2bKys8ilNRuKeVCQKx/46tW6n1HqpDGhD9Q8ug10z0om2SVmys5rwIqW19nk
YpGVWWfYJG4BLMWk60R3AgEcAKCFpRGSKNTFVEVborjYgX15FfZoObnje2r/ns0Brg7pv+hVDsZQ
O2ETp9a+PAvAHBNTR/bbaclEWos28hLFdlmiHPFKa6A+jMXe17RGNVtqH/E1WEeJvT7Nb8YjDtyd
9gCrWjdBWukUb7UNxGqUX3QG9PSCunlksJJbz5NoE94fvvtO9QR80CX8HEBQeTA+pAlInvOjhjAv
GNvlwGAhmZG4sNVf4rywSyamHQ6bRcrRq2Q9+sRqsDqz89XetEfOcg3hJXZ+/h68Z9xipYhamBjh
lPRMmvmofJaxDrv9CGEXFjYzh/5oIfsILrN4fCq8biU86jLOjoyOacmoMQHXP47RgFon43IWf25r
etId95N/+OlVv76E87Td5khbUkySWWd7jxiRBkBqxglDI67JANC1N4CSBz5YzrL5PXieerwcUBUu
/5u6z0wnxtbokJ5+nPz8l2i2pW8lQFsJyFOG9Wx6x+FZaWxjxh8XpqlGJE1DCfKFSAyfCTMXVGBO
wKiUsFvmcZdobPXrMzFhiF1SUDytmxWAvfiYvjJ3NimPjWuaA5nqAFGgEhgmPq1Cagz0HTqMQQkU
70b9T51ODMa5I81xQAGs8ANzK5juXyzbPSXWFFH3qOTVUJWrGcdnjr8sxijnwl544UxVXr0+197E
REclCW7OqPTX5dQXz6fuV+k7HYvETNCs94qUdetdUIujQqXuoNvP6A4B9Ui+orBiDLivfPa9d/Bm
w1mYScaTODJsJuoMEki4N5NN0MGXFCYh8qfn8IFnfdGSxaXYPu0TqJspbh+BF9GO5y00syjJHNCe
WEdxMo2NEzL1vLvm0jzrHMAViS6N6YOcuWGd4DU8MMFOXwwIjA/seZjNAeX329QIrIKtTWTwGbJV
Krl8hmgsLL7MWmRMBu3riynyNDMpmwDXwxDLutmGwt9f9gLNtE/9V1ZpE8u7USfUGEYxZHyszMM6
HCMeLGvX/ozJEmAhkvqufmuAE9f67GAQ7N+AuGLpEHBds2DvW874cyekEGTPLBbcWBBF9bSD95GT
1CKIYWDTxtCL6ULwv0jY0sEBNYPuUa1mi5soDjqr1f9thARI+mlHkv3Son8q1+1jvOn/GKMR7q5J
oUN3im26L5JG2DFXfk3gf+dUv0GEERj0zpfgph4zgCmH6W3thLPamrijmBGb1ckqQ627BcFiTo6Q
TJzowhfkZC1PvJuITxPlcjONdlxzJQ2Go9y1B4C72YMqjU2217+2/xsidbvmORdsz4xrLnqyzPy1
ptUDBWhJWf3UPE7i10eIQHS6WNCgEUqdMxytFqWBagBeNCW8qEhgWzH5AFgXWBduZnmzFIN512Rw
eO5WH3wHvfI3vqDZcxOK5JvSIna8W5GjsuGPAFtxdE100CiQesIQ9BRrOAXapOWiw/6z8AKXcO7F
0JO14Kr2jJBv+5yfWbuQeshwT0SFav6CIbCe2SCUmudIaTQ2FOWN9tb6HtCWAxPMUNrgPUmTJJnm
5Z34FH3GEZzVG7TDzHJLo45SX2rab8KAKPrBsAT4rm7WiMtF6/S/ltwCYQDEi3OTY4ItekB3Akz/
pCPdAvJqO8YLctiomryVGoGXz2gy6yjFz6zI+Vqe0zpJgTuWKq+K0yv35s8iKJGUtwwZ5VG0TDq8
trw4yqivBWQ/v9wHKJoDAYjEKGmxwrBcVzfxu4TapjNIQ//bJO9LItnHbPzykYGO4KT0ug/FnEbk
MFLpLrznSzwKH5mSV6VtBXQrFB4e4h0ylChV93mRvbv05Lu0dDErjojSoVENm4EDJgHjcnppIfhT
VQfqkEpwRB2uOy5JOPJWnXoEdXRD+/SNmu1Fmj+ler9XvFZz5qBpyIUQoaUdehkBGytVT6b41+oo
4VAmer0MN8ThNr5de/BwoeFBCLuBChnce6uoNDkeyHCBBvo0NYuFa9bHWVm8QoGyw90rLvzrdZYe
11J+x2yUcZ+bc2tTqJW9bpSI6ahfnz0hDtea7YHZTNbodeUhIxMXk9ISKnW+GWh6OofokOYxKc/m
V5ZFNdw9rTL2qmsJODHKpziKS5pPr74ivyvWGHvEDq1e3eLFc17LEozmoA4nCwwKPqczbr/RECD+
WPzB8p3a6TfLw3imKulemgMKM3+wCUuxVvYXgAUaWXrbx3E4XQ6hE9PtoK+olWq/FEqVbfgyb0Q7
R5CWvYShguIoEP0ILLf4jv7vTG3yuiDeXH5Wm/Z2RG6fY3zMEBYYzxDGoKFQRPmPkCr8yw4flfMg
vNsFiUQ5rI3USoXMXBSbc61BZlqUy9uYauxrkGBpvucpV1Gy1xY149LyC4Wkfjm594V9d2lLHnYH
hBH43rgipBobvUIDcxEz/Uu4Q/00Mb3siyyKitu5jKjFcB+Emyo9Lsfu6xzwop3TqFcMm0WSMsCT
14qHYvmbUJd1hGefiMiHhLIG5FceTJe4jMiT7bzVyFzjpMPJxhtLfO5dVNS2borNH5Zbup5Gxg1T
gP6qSYK6IIFAVQTv3dO3yVuNDELrSIxjJelP3fhEnLa46h0LZf1EtXsamHRUkWB4k5a6yAkP29Py
qE9zGeCSZ6Kfy1e+QpoQIfbJzxjE/WO2eb6u9aJtqlEPJl9r4yuzZ4WpED7nVWI2J6W97rVJsHN5
hIkAiyt+LGvo5r0SJ9QmKEKaMfFsuktf6+Yllhphr4jAZdxxtDxthaIz6H/YcTzGYyLI1y9XBOQt
Y3IBj0LnsQ01XqidXqPpHiFmeBGpi/yUQjO3F1J+woKFG3gsRpZNqBUzDypJwo1Lz5wU/VE6KLg/
G6qlz94O6QHV0Mh6+Cf3N9BpBCjA3SUDmP8eKQ2HPATFM+senEsUmGciYSsElDEIdUBF36iRLzr2
CTR8jy9xAws0ggThUu4rAi5auUKWsfdHlaQRwfKahhHA8eclI0rxZY1TtnMdH8oe0FQXm8djm/l6
16iUXDhdjGZKiBbQxua7aUTJ/H+fS0Wu2W0JMd1vaTGkarsLMg+mD8BrtvWiAywfZ0RG0e1xYb1P
swaC4V6KqBzOujpyubi7f6OggCtnXli0xBmkujKcepOiUGznksGii1A9qlyR0hg2HzSI33xwksaj
qvDH1SwAJHgSNZ8tsVysq6SK0KxN4CDbXuWqdsPXyfRODcGcl9ZtCPe7PcJW+xALBRsUFrU2tit9
O7bQr5y1tXtz0wlpgIQq+2V4IgYMkjOP1BRDrIUv6Br58Vosg20iFxc4ajmV/Eli/2bGTVC6p74A
iaruraA8jNMGArWO7v8f+y15F9EdzIVx8Czhh5SkUBEV
`protect end_protected
