-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ev3PqqNzK5sjWuivHAUP2+OmkefofQclinLTdbFFfkb76pVvXQ8LjeyxIgPVHexw/1jghhzmBEj4
fzezsWrpybEO9mLUiDxrzwaWjBtHZsUyV6d5f6D/bArcubao0Ou7XjyfGDRHQiroXs7yYVXyWufL
QwISeMF/9COil3n2xqbdzhqa+nyeC+MxmKTcngUpwIgOJjsJavRytjXKkV1/1q0wtTOixJPidniC
WCpbYrCERT1CN4NHt+FyLnwAQAEE62WlRQNHKRwwgHTtCaz13ZQMDkOnNW7VgxwMWReoJhuJpG4I
NrEDGb0lgAMN4AT8CM7ypWUa/CtoyCCvMeq9Fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
rurTnwndIEzx5HGeN2kvjCEDbos3FEgV4qeYGWE1Pnl8br05VOk2aAa+u6QMXini2+fYcwJ40tJO
/0QmAs3+iOnxJy9EFLwtUAhyVgJIxUKiHbWlTsOWrhFHmehyVCA2R5SIuJLjmfWaYe1ZTR9Sz1gu
TFBt6bOhx8P5TLWTohq8o48Sy7cSBRlZaERySRmemBLXgRrugtQ+MYMhb8N4wD159cURL778ydQu
jgYRw+6x/a5YmMSlHgxAZYINLdfRMpxbTGv7kKcKzGZP4NMVz3Eq4kGKczcjv+QXudNVhzX7unb0
G1ztFctmjb0r1kRL6RI+Pc6OP2CrObHWa3jPRLip41ZiqJ5l64ZbgdD8mXC0TXkpjfNSGvJ/+oHT
rCkKTOfDTugo96STYFZDZBeq4lTtEFiaiyVMWxDSE42TCsYKcPED2qG5erDqGLsAUD3/VuNfYOEr
tMiR1/c3CiFTg504FZ3/sjk15eTJxLc7wcfZ6e6qImn0mDqe/a541Haw/Use8W/lc298Tdi167dI
Wk2nQgbexh88bZEQ28tfHyhWVunr1PQAYFv9oMVrALw5fVTZ2u142ypXkfIN/1AiVjjN2tDBLqbN
FxR25vQ4z4oNinD6CBQGfNjP9sJj9KKR6+6LwWXuI46K/jopEp+t2+g5jkKXHvE2796bdR9NGvuJ
q9rcYON4kPIJHmftsxBmj3FgK0isCScG0JQLzd1tD2ZRRkxVyEc00IEanH9lTIrx1H1pAIe9pJNf
nHI0+sw9gP1mh/PkgzXFZvZreB/H/mziikHKNJi1/FiB6YqGYIf+MfkLc01LGgizPF9rYqwocgOk
t71XZLh2BIe6ypH3ZNNZtlmqc5EBvtFokl0WxfDdcC3i3AZi1xuBlgTlJVP6U9Xv+hufw6d48QSR
kriOUPJTb0zwAlZvEhObvuJFWHFuBLhlw+Im/XzOYMqUrjSFVWTxhuv7+IbqWzA9zO52Q5cZFpf5
1AOG6CiCqVOwN+tDoXye1C90ZSUhzWvf8gu2yq6IptBH4/PkmwpVRGoPZhfaYGSQOtLVPBek4zEj
cgoUxvO+Oy8XZAQSeTzBBpRB3evHzrNynJz9MzFf5Wo79MB/THJ7z0ZEPijcFUdBV8BcInZZu4XD
2zsUVBTS4HPRHw2U0B9MLqMRkCtosVzEbWwni9O7SJEizytOk+onuxYbPweZ+Po3oqu4zkL9Z75P
5a/xEbFdFUbCJBbuNHoEjfDtGiTJakWaEW26cUk5gZBIF6MvzRx4R9D0PqH71FIgPDhcio3FPsDG
hzPeJmoh2OLbEzlVWNmfYuJGe3MMf8uWAIgkXS54jB65wWdKvHZJouGX6NmQjdAzkZ6pR9Px0C2u
WCOemAYmxtrplXk/mjEB0aZ3X3hAvLbrON8AoveMxusIkrbRUn1CbAiOpfg7fFmF9vqOYV6UxeFx
5mja83jL/XQy+5JcjWGnfWzTMHWX+69anVbp5IsuYoHQMgSQdumtXcNM3jQH3LNhsbzZcI/xyDYs
/5OZo/uqk2bKVDhbKfmb3U8F1iNwBLamD8idfpshoNQLy9sNSELRoRThwKFUlgTjbnHV4Qa9BrCu
KJMFzFagLPia1R0TGrdir7SLGfHOPwFEIqQpqEXyRVkI8MDlFUT97Y0dCaPePLx+qIrKmqXyVZnW
5aNMKC8RNcr6xPJOet+Qf4nH70LAVrRNdMCbDkdLZaPZIHca5/ksqYUWsg0cNOUw3BEwptJSRIkN
naxKQ6Ra50bUDw6IJF9TjZlhISD32Twj3Hswm6/XgD0AUO5HEDlp8EP3P1og4fq6/L9dQyZxWKEc
+vC5E6UmxMsKK2qU7ge/MJDzeuOn5nwMG8uT8Vw/aM88c0wYCkHY8RfcMaELqutR5ysaVOY+ldGO
iq2iRyoAxSoBQGT9FmoL71RgexWsdorCf5agx+uN+WVgPdCPX3oLoTt2qAFJnIJxvTG6pK/bwFvh
m0flIqiQ6dXPhOCoCHoBlJJQSJFRP/oY9wSOxpbMnj3NcxckB/7UfGBVkMOmst+T75Smg2mcW0Hx
pjAYrCJcMKdTgqf+aoy9pkwy0GWcTBZpzDUYjrAOy2mxVxGluawVDcFEdIaUsQAy+Cgs8ruYoYBT
MDDnR8Ly+GuCpOKb4Z2xppR2WrBzFXvNc3hI6UWMNEPCh2+ProAs/lX0DJ695qAq5RABkBuKK4Tp
dAvktj9mgdt2RgydRsDQuiiCiMs8ZgyIlzOLw7ru8qX1kr/WmbY5iL1llg9RUcfLj6rHyZKIl94S
FFeGZ0zK3txj8B+p0+sQc+JASJiL/Q7DpoHJSUGC2ZAmuHeoCLv6aktFVVFMDEF39T2vPjaMZP9k
+fp1aYFBsT4CNgV+7hWRgiEqDDr6YA+jQM9GNDk7+Wr51GK8hmPh2BxRlj6tRVHShmmzTS9CrQ+i
iznUgjiq9VAhs7s+BqJ63PYc4RmyE5I/rqFFF5+FCu1I7Zl15Yg6FOygygL8Vo7A+nX9uralBt1W
5JqrUWdet9sXo+++Vkerjd2zrpZI4c3wVW/5uyDgbdAD6KcX2sV/uc3qCeopHkQS82g4aHLxbPPy
eX3jqUbmbGJeNqRAkmpsO3WLTKePYvcShLGtcwfmVQ+fr1wPomQ6yBLa2N4voHL/Xf13VbukPT5t
bCyPC+RG8vfxQQryndXUPgebCXS5Jq66I4AdlegPzHtiijkyDoqn9sj5LgY1RdubwtoSyjLCw8l8
e+iUziFoum6+GxacEhCSx5gRQGROGmmzYINo9BTgahx568sZ+S/xQ9GSV5V9pfwjLBYx7OI+GYf9
p3Woxn0duhL048y0a/KhCrbtuUn0nYSEtghu5qxC6Exu2VoP+SkErQ0O55tqJ4qAbLTtidi0rH75
OxCabqAoN7/i1FFxKWxoO7mCrpQQDTKQhhbDnXOBAm/uwPFpwbjuKhj0WwWjYqCXE5DRw/6yOcLo
iPUcgJ3EFQKC4CseQLH8Y0uBX5ngkAVsPgbiAsvvC8M62PnwIQoR/2fP4tJ51QYqVwHokJRnVC+d
jN0KbxlBeWYA2ODaZK8Y5reeyAsRjO/UnMlb05lcyOmsDDbXzHvXJs0e7Zo5Chmg0KunfgE+bAYa
zCoiNKwLq2cjjjglT+ilJrAVb/AypC7qU5de/f2NXGZZkgyW0x5syed4HhSfFDn/p7xHY8T2AkXQ
1gMERhzwS67v2WF3fWKvpQCixPHJuOLCNgpYzlZPVXPcTM+HF/Y6zmPVxiLIRXW/04iCsmwGvXy3
zEHLoqV4bEL4Jl24mOmOLEoK7FyVi1iQpk4BzjPZxaBJ1o4NNwe6cECZ4Gav4bOSr6Y83W9RFD8U
rotK8F6jacdMaho98kWlWr2wKMIeg7RTSwfSWByFumtite6en0KtmxygS8P+JLI99DAhqSGwZ6w+
2PULxVTaJQ+/KT70yHQ4RijCZBi5Se1h6kCIPb4HyfARCITsoNLv+QJk90ZQ8PIzdSU7b2EjneM1
MyN7/AmRnDe7aAGjvglvtDHkA0nMfpnq6Cuh3VeG/cSJOlzJ5UiZrPku8FTb3OJgUrOvMW+VNUL9
sH/x59g8fRIh3ywkZlWZ0zNjt2vb34wD00RKr4TGuCd+txyL5pGTjzLuDxKrwGUVGYhN6njY+yod
x742O1eASM0VrZUd4gw73XUtr6vOwcPbL6THZy0d0BbZwREb57zGR5FJzrEGCkm0JcOpzjOFmPO5
7qTkjNwI60lv/zU/G2pC/REuNrBEkiTjLWb2jqqUWE2Lq2tRpllXJymFN0clvljoYc0VIBw/XDBT
xAbS+hqCL/KXDL5N1+vxRocRy7hg1/1IxGKFKQt5t/7tHRXtmYPlmlZfU4AEQ+JCODNS6xgHt/qj
SoZqqwUBTucJN8siPTQyiR34iiocko4+7ncA4e774Yg8YIv1IuT6hkRhd3ZgTNxYyMheSNkWKNAL
q9YzDYlgVRu2QS7BNW1XYkZlH8EDfDBI2drpbPcqS3uT0jSJt0uJ8Nq9FyOtw3eYyAiwOiux6UWp
Uy3qNOf+862YvFBT7DKlZ7Rmf+uI241lQN7W+IWVU/3o/Pt5YvM/7nOXSrCaj81eWM0p0NhOxIg4
YtIWmf8QjboR3kwsivlfFan/2jAwA5EGwCQyAfjb7PS7l76pGAtqUxkSjH4/cMn8GC6NXV6120br
rZTDn35t2+buwVs9qvGmdx6e23okDnzRVT57ERn9+3DWoA7Qh5whzcsZKfkVzrDM9rWiNaRHexez
JM8Z3U3Z8brqv0uSU4ypiaQJjCYM4onvVvsI5/2R1PlMD9Kg+qUEa0idWMELC9thzxMPawalRXXY
TRG2rhroOEM4NixFDGHP8068rK6ob18rFTq2pjZAONZ68KFI+XPFmiqOpQGAywkw94Bz61y3PbbU
QdwjVW4pQx+VhiOz8LpqNwa8E4WPRGYheRBIIjHYQV0ZQExa+b19tb50kItq+8kHSsb0W+4OzJk8
5QqWmBLBFsWq78+/SbLjEkO/+HEPXm5EaxTJDrJwKM6DVs4Eo4iu5wipAZnKYiAy8bGsQWH0DyZX
Z0bs4+CiabV8BcsyEG7/oQMrJNDvPbi46GlU1QQkMJyy2h7zUP9o4zMV1Hk8t/ucuzScVQVSo+Qp
8EAcFE3UJng4pGyjLOWCqgXlMZC9dJGlYq4ToWAH5+CXIehg2C5fxS11hl63Fdypi4cTemG/+Nar
BkGm5pRlRtoWbJOb677TyaMRaYbGiib1lJdHf02NqquJ0j4bdRLanpapL49v8986dKozlH+LE9zI
FRH7lBzb9kJrLa8b7CEV0j80Tamud/NQtEK1l9J6VRvpsbr6xx4+3YWJLhg12S2c5fyoudksSL01
NlUszCx/XA+jd70UdtuDqxq3wFFGJP+NJ6zHS0kAPUGWSozSuzofJDD5daiLhnvsGD4EnATrdM9d
ON07UFav+NenoinXFcgTyAWQEpMwMK4wXOWP1gJTUkG0idO63WvNofSrkCzRIuVYUdxGo4ePnNn/
UNVTbAickvxvEmA0tGGiJUFPjmqlHZ8bz1y9EAtjIVaMaiSGPDEDUBIqt6jCDh+u3ESsTgioYn0O
ebul3cTqpYfzzgxBOALZ8g1d5CHeAsomp0WXDpcvPjj03Zr4auB0zOy1A1vr0l19cHK/cSnCdMRF
8WjP4KREJQFDaxG/MNro8MhVfw6alV+6MQp30/j9vCnpFLBZvTKuulN+e1UQwNpWFObgxiOSARcV
4uHSbJ3wiLVSevU2n0ayWmHWo6M8xAj7saSuzaFUNIpm49ZQ+rxqtxV89q9fyLrnm+g/Jyvo6aot
RALUlQEhPPLF4FaLvsqN13Fi2ffgiff267KVxCIw1YrRV/feL/S+Z0IJRmPwHtlFf0M7L5qotHG/
kFGScg9+zFaFAUUtNozM6ikUHojR1zB5iZB5P5Dd7px55OPOLbm4I5K/Pir6+Gf7tKon2QowcC1I
nJTA7AH6SB0hdnGPM5TT3FbAN2Ou6+dgl7LjEErsXeEDnktbjmor8mm7KBAWu46PCnbnG+4icpk+
YLz1l1psUthgbkaX+GC6OWhrPpnv4xieZHEt4AS31YDcBQ4zbwp/ivfbv0hVmvNPGT8GYnwLdLmq
xQcQj1+Kq578JfBsR3XnEVqCCSPDO2OrV/eMVxQn5gaJ/yioSS+bFskZbicx+lyjmYAu6MvVbWYb
HneCMurD6iDdBwQX8SHowVqvqfJqNvbPHUTA9Bv0UhLCwzmeNL53P5ShJAt0T4L/9x3rlsXdnqy4
4mNEb2HQWt2gDK3RWRF5BZnzGfa/0yuCQiOnefbu6f6aUx7Dg+96x6Rwd4SSL3NFQsOdlB9WnTcs
IrT1jc63pjCoG/BBmWI03xSuKaSLgjfG85L/vax1AZZVlg5r17794WNTRhEpGeOy0qynKdyRUR2P
Wg/ElIe3me4mTcQklScGkvxifXVbOAGgF5zaPHD09OkzCAtcGbPyOXWnn1Jvfpcl8OHBCljzurc6
AKKgz2lX9ahDUui/U2N/G8JDkcOEAcKHhLdMaMZV+m8fYlEEQycTKe4Lxr+7/xgR4ETbGcogR/Uw
Pdg0XjdUwdGbWs/KssI8llICnhXYDMV9VS77wEdpMlVEE2BSBvllmAIudqjryQSSc89zwHUr08/l
IhKNV08XUyG0ree2Iza9cmlxmdcAvIFQwyMTZPA20DnvWiwswSBxzUzyo2tqlLxQBm28nb/TNHq5
JW8+HpTZDp5Zlq0k7hHt6VcNir+4thFma5qnTSI4FdZHFMOxlXMob7E2KEFpnqXiQMmKJVYRLfP8
LW13mPPBChkWXjECoOGW+c+F8/Vhe0UOi+jXyu6Syv2FtLSJqE6/0+hZ9BwCQZHNZ0ESHC7rLw/h
Wgt3zZjwDxyctDI875K82eNPCI1GGixx2a1POm1jZ8pgRVgmHYgG05ijLdBBG9z/eZBK4o+pIKyc
RfXfkPhqdwp0O3B6PMqYiDNI0bk0gJnFxFKyGbzdxjnlpnPwwte7TEzSeG/1qk9OoUxXgXtlvKrG
NuaaOUuXz3xtXcIbrTbkduzaaMQ2o/YvJ3C9UYG05Qjg+ASFatSNggX9M7JJ86mVbPstqw6tzJHe
b8jiZqFXahNYBG2pVdJ2UopBcU2ew+D4TL7zk87cB2IBxl4N7VmMIXOMts1Ziup9hhH/f4e+y1jK
DtDXMh/RzhewkhxDcQeTSvm+xS4MoCwZGC0Yj5k2TIjos56auQH2HBdWWiqCPeujNQ4MXhPehUaD
HFfo8vdJmNrDkaBrDAwXPVesUuhHOB6U3j7+oi423vSMhFs3J3Rd7zgZAmQBmkOk3acajB5SgXk3
bptR271OMvQnvnAeJAhJ5uZAJaV9EHB8ZPVGZbK/6P1psLD2Yh0x3SeKd6q54M+PLfDIw5OL/gOH
HkzjAr6sgnHevtRoCNk9mgRUrCzxe75GoCLcH4+SavjoZpFPTXMWXSEpbqSGMlewirWzewBKWgjX
9vN74myGV8gFxrQQZddpIFmvhc3CmSqFcGXEm1wwg/MohyDsW6aF4pUIKtOKfcehMWibWiBlrWiw
0Pi8CLqmpZKsqVY+wkTfe6/OiHuqn9hMVZ3wja25F9Msf9EnMyn92iWmMucwjt9PRPvwIZNLUYvN
av2eFsfmZyTzze2IaSikbPusXY+j2BepFkwGowV657tZu4Hfm6iOsqT4KA87PCjoOAXmo+sKLv7r
p8QqPw7swVQUioOrE1ggZf+epnGpf6z5PpxHhphRWpt9IoCddz2GtvFMBwDY5qUiP+Zf3It192sA
OYgy3KxswjwAyhZ1YETexvRTYElqrWw5GKnlt1NSRs8zhCrGO5aHa7xbHIQuZ2jMAQ45VBm8cuwO
X9fGks3Rkxs6dljCC8gJwvDVrn/Y8brVeXRywj2FPSBxZxbSAiHL5gQv0nwVqPRptD15gOBwNIhz
LiC2QMdOiJzPKZw6EelPhrR+cStGBeAhumJ+NikgnqSusAcA8IwmpSLwm2uznL0tSJxXrSILXYBS
QVi5ApPJ1eNsoD3hq5ozf2zLlK6ibHLJzutPsAPO1cZd8lrn1jf8uD4EXUamptIjkABQwsiYq3Pr
1bDoBQW6ZY2ipQhKBXQfkqNoQdzJeyqDgVajG1wgk5GadwHWZh+FSH/AFWOPvf8dq9sLWNnuOQcx
rXiCuLmkMN2iw0sWyC60/u4lV6gBzy0WrhHmAiTOW5GtXepYoECZHZNwE8WtaLPuk7XGT5swE1z8
anzDmNktjETXVc6UqjmNQV1UNuUE9n62mUWO8Mev727xLpjtn+a+SuIVDIJVaDpDocs4e5Ijr4G9
5BLmTb0Lzy5dDs+o0kRR0BKd4DLvjJxoQP0R0nH13Vos0IyjRyyk04EHwT8OAgaYzyLbFmENdTia
aHYXTy0JAmIJHuXt9AlfEGBLtej92s71ciP2czdJL4Kc1QJopndbvHoCZ6ZTM57GqrukLzmrztc9
ial12suCyk6s8aABUc5OYysJSMzeHQYp0HiNZlrG/wC9W/QOl9Yl5IeII8+oIsDhosvbCkcnSAQu
Nwmn+TFGwG6HLpoXDDOCWujIJoDp0srvD0eDBrv5mr3+6bah156Y6u3AskDGExMSeU46mBQga5VP
+HuxzEsdNbuXnfBDi8/EvC+4Ncxgqzr6uN+5BiLXZfk/d+enn9eudkgofjWQ/wPjsQJUAT+o0L0m
kL4e+ybZN7XZqS7llbR92ArLOilrfLb3P2oA8Gk1Lp7kS7XvPboT9SNSxugmN9yzGqhRDp8G6Gxf
oVOmAZH/Zrmo8GHPL1Z6YyIPze5LTrZrHlieMuz5XmHBrLN7eYAXLvxzRLy+mXMaf1UjbCz6JuKy
zxOjDEuo1ZiRAOnk/eecD+bqyYPsk5VOJlgJNfRQS+Jvw7QwGUw9Uif84q7q0jPOaeu6MgeW4STe
v8yCfL40lUUAfMVveqiQotI6kZbBpPRIvFxyH3GcMo27PpOZstPrHtDiU/n5BzbuhMQNnwyym5Z9
4w14+R+ST8xxhtxLNwNL36eMAwh73JosL4n5d0OeJkqPQdhLTBjX9mHSL3Upwof2KYNWtrhT9mKg
lU2RpVpr6r/3jLNk5gxzg+/jKnr1s4CzdX2+dUcSuDG0RtKEwX1jgxF7wFY2zlRx/DhJZbx4fquh
DRU0b+BKsDKLShhkAPGhHSyY7NlRWkj2ibBrY9MQjQmKPx4J3VyVzobZX1FmJP+6doLUAoN+/pjl
yTr2ASNci+Ea15uukbgg2OOCSARK2S3rosfg5jguW340Rfzjlb9fxX2IvRqq/Kfz502Q8IsZCrHJ
Eit51OCmAPPAC4OipiS+yl+/KODGLTMFLqkBG3VioG+KJT6Avddff2ogUfCpNQfTUmLVeB8a5uZp
5JW0l3jla3HddqFPaKKH4niESxQxvHGh2D+9sYDr8I92gGJjeSMHAIS095WM7I1G6JMRtfKSbbPA
Zb1tRoWPoPpy4Ze0SzlL+8cTeL9aSNBIZZWuxejwllM2vEjf2qaj9zvdRSjHyNcy28TpLX11nVea
NTJLbpZ/+Xy4KlwFnGvkBqbZFEn+kAnqzDc3Dlr7fDZtDE5Qub7MOSWmvZvuSdlAjO8Hj2MDfMIO
Npk+yeZzmCbrOUtrn5BW76XRMiC4I6GA5kpU6bFDrgauTDT6mdfOI6PbpF7UoAFdIJMS/JuIy7B+
ZCbrTmeAc6yd3xag4qFZOEYQxSOaZmQ4DDmSNfCAFc+m0TpwTb8GJjycWKYDOpyivnhMkkceGUl7
xbvV5aydSTvl7/UBqrH/WWNzM3rl8oKDCboCjAfN1+p305QVo0h2NbhFTyrNM+1Bcchk5aI+ewBZ
wtmaM3MgrResqgmD+pKWmXlztXCJOt/QfonSMMaiXD9jmopyhHUW14PrxSgEkzx1XitxVe3HEE3e
/OWUhSTYD3s7l0yqpskMAUNUghN76wzpjtwJMMV+BbsAvAfuBq2eF214YAoFZUUAw6G5y9oCceTt
ykEIwQBuntpiJ/S7TezZTLYyd/q6WUlFVwxmEZ/pDUaKT2ab05x5NRrqnXJwfhUXQdsO3phVbSkY
ZRsjAGkVBwwRDONMfGOOXCylVv164nS1Dr/5uAXSSc4VvEQ2y9vG8k5sAeKPECCYfYR0gNhK55cs
lKoHcZqleer4tH7oDrMbAJnlM2H1oWn8lmZq1GMLZsiWeJLoNiBXFt7s52sE2GlLDUQ/eJYvVOYH
TZy6qYdPxMIndS9OY9CPf8POvXYXWKu+Ut4cRsB713kyw90742RtOt+h5Tz5ZiYsheFe7uoi1yD0
Mj1c5cfwc4DOobL+6HZQ+61MAM6e+qc8l6dn1/E79IQdaZn2I22oyo9VGS41LHW4KkgDa37TX6JE
fYTuLh5aonXGxPPD2KXw9EU3VFn2/ns8ivaYO8nJlcvuzu4sXA/7SoObLz61/dfiAE0PaTBkQJIm
BCraaWlrtDvr+6wYYPmB08k3evlwzcjiYhsCyYKxSVtMyhbZSWvmACGec6BqmjXVNQdtTnqtupHS
77RjHA1X8eTVVITLIlJpIQG2yQXZi3M9mNtpmH8ApdWEUB91prwXf/JRLDjPbkCjV+8vfXPGoVRx
9D2+kEdh227AKN/INZIhGBS94AcVKeuU3PWYyjDMy8lbbTnrzLTMlpVRwEvgaE97RSJJ/KUZFfw7
NnnK4ToqkjtMAb8cVsqbT+K0UsSji5IP29HQ0sfDYKsgeGKLoSJXCwOaJl0PJiZpl+XIrto2D2iz
TCbEvP9Le0Dnb5Wb7Ieh5bx1gAGs1nA3gOkQqyV0dIlqNM9q+lDWToJUJjIHs1jKWW1lfEqEOux3
UAPM7QLCsj0HfqdHz4e9Apx+DBz2aA2wJv0PVjlCSKglYfysWNdS7SXoSqFuav1nJMQInAZDP9s4
eW2Rl9ZmwRVFhT2jcG0RLmduABSci8Nl40WyYHc88PxalUQT5d1C7FejNLJ9fbVnTILNt7ouBq1H
8k19WHY18mHXj3rczEi60E/kSJx8de5DOOsVl4CsnYO77bXmJPeYookOySzRB4b7TXoGuoj9CXtU
E14wjvqS/V5UxMcEycavlvFmDyXcqizAqX5BKajWLdQYQrLrPOAGigk8YT/g+1ALVhmrw18lPsAe
ZtjMFyMPNJ6mvdnv6usBhZwlOCWBR5GPNojy4BX5k2VehRbwPr5i+lKWcf+mnBQbTx0BJcmYjfMs
MhWOH6gr6qczziuA5+j6xFjDp9gTvAtGo4t5qtFgefFNuP4LhVFa1jPoZKTkKDnWLjX5XHXtHHoO
aVv0L7nnehrFne2M4rBpwPNHs49o6C+ArfdQVVJJ2M7KbaY5KmSaaTw8DdAduyydjiSP2XhMD26h
K8oq4gROcqLBGAHXkRoDqlKXDtR8IeJ4Qj/ZNfO+T4Bt0O0DjZ4N3fGKvwmUzhNqhfEqD0xq85Vf
kK9fNmBgKVN8YhuYt/bgi2qE4s3PzSkrkIAgfxbGD+k2Sa9Cql+Pg/sV+Ux2gO0bAIwBc1Y1cns0
ixas4lHy8fyaZA7hnJyOH1mLcpru8oihitZPzcaqdmE5I/v/y+/H+EI611Ha2n9BzOap9JJO2SX+
T4F/gBRB7ll/RE6YRFmOtUU6lUCkoajzbPwBUAY1YBPXpoFzzU+pNm9rAC1C/il951rsfzUuZ+BB
ihOPq1Y3n+tjTLqdjlD1MVTyAu26d6oxf/qNVcU58zDNCY9xXTViwu3kevl7Oab6oR76ez67oLHK
4d77Cvf8EKJOru/NYq98Kus/oLrSTFRC8c4dpGTof4eGLLWN6z/OCZGDOuVCsx0DIXGV9LjDGs59
itmzy4cu8/gjuIU6UmIoSWdqa4IwXojJRttqUFJ3PgLFJFjw5Hs8DI0chw6Pl6pKyVUHCm7eYR6Q
Nj8soplJ/+DQRxVDEvB8oi2Iq81+Ll0TV7EeOfTHwCWDkuoYF+3991uXABimdeyWNZAoL4LrpvGu
VZG1WRRguh8pVdwkOkXnjr+/gW26siMC5QNEbPT+HpWudQNK0ESSM+dVB8IcWvhzS34G4hdheqTz
z2x7QFGyehD0gIC+6SNzlmYAWhRi3AOVSAUwcCNdgN+xRHZKhllS+XUnF4np5bIAJGSE/wV7TeiG
4Cp0Hkn7OFt7DMJCMh2JnPdccrm5/Vzy/VM7lu7deO3SeXLzIIaTRn0hsRyRLB8OhiR8Qj7n8d3s
9ZeSzJff1FJ6KaZglZtGnuxRyjWWDY9JF8NsT/yMgNXR6RqC3ojlWglXLxf0OUvqSR04BhDoGy5v
D5TsNqiw+pxORt4siY+JB1zNDW0yOXeGed9tS6vHUpueSdUW7Fbn6UCbhAW6EEWLrcW//sXAnu5I
Lj1i/Sl9jSbS59/jI1yES23Xx9l7upwpXeGByB86yrbwNgbQ9ckg4p+Eb24L+mR6I+WtP8h9NLmE
K1XTVpYyqV/IBsiV/jfJAdJZq6GYSajqEqc9C/tSWa3oDbFJBc58O02cb0Fdpxo6UR4LVFoQkAJz
rMLEh1k8YKkZZylPXViHA2v1B+AI6tP7Qnke6BiOHAbnUiaBIQrWFsvlIPRZT9RayormtGIVNsTq
NoOmbt6rMSl9wRcMffVNMbmQFqBeYdZLZiiCdT+ZUJjzhQXempqB+8RoOebD1ZonFZxRRxeDEEyn
360PyDHpE+WCPPxrx466ZJ7dWLOI7fis6NW5kkkeZ+v+GIYfir+pdSFeqfNgX75QWrxbcExflJJz
lX0APr/l3XsB8w+3mw/HW+mASYhfkm05XJcUJtyESBreKBN49DJLpKrzR6x7WZXavsB2dFW+tsl0
M7ZobBjw6HtgcVnmOFYPgD62xv0Pa7wwhmri84EJZ1Hkc5nZkz3688bqdO8VVWsjxxDzcT/VDDmW
7QyLs9yOoOkI92HStszcua3P4tYXckgZiI3sTOyh1QVJG3IHSzcngYuD3wHYBP3ZE87At31oS+80
ADFj6aHO5acaucochtbFEGiuKadAkNK01RhEFbw6M1wZD0Wv1DHDBMT02Inuxq2NDCMCt7wjXGKe
xhesGbqAdVqSm+q/ONOi2F+YPNUPBDihKIIrspVbmEG7U3Y6H5jsZmsN1g4Z/iqp3xKVouaqJCF9
C74nwVBE0tbjpNwIq++68q3NZ+THB1b8n9vVY8A5Sv34t6stXBIKkknImF9/EX6h58zyeXdp9bDB
gN0E5Ij0YOgC7CLbE4f8oTELFn6tzqQTKFZw/vUpCwybxCgDVQX/aKHFrLgGtlT3FjUQ+DuFneuE
yzyORa3iolIG+tB5bth+UoMfBC8VbnMoH+BdlT98Kv9iGiQvTr7FxXiR6VW9Kk5xcRrayUXu2Q9T
2C6Y4TzddspJWc91YOmj7gJf1tPYA1J4gaKoyHIjboEJC8umx1bC4pKzU0GR/y2VP/PUJ5e27H19
fD7aXnCnzz/l9mJ+tt05fxpk4kOKuBUDlSWhy4T+ZmGBzfD5+FxODekpj4DLCSbQkzAnorWBpboL
rZ4NAKZlX468RdoMZ4NAOS9sDwN9rq2qn/3Mpx6cC90PHZlaHgjWkPZcgyOpWimJHelVji31YZDk
46Q+x5e0aK18ew3/u1u+Q7pBuMVSqFJg2KQQjGq3wIKw3P1oWJlbhLm+//C3bQ5KRXPcuDNj+NcJ
A6R/I9i1Thwf31gOt6WBJVFDqo7P7sH+HsNwY6hqU5LowBZxEDt/32bpWDkVD1+hfQnbGG84otC5
Llw/ptC3BChPLkl3uEvDHhfdsxts1kMvyE89CVgq/M13HTpbHBMyr4c7Xohgm6kIYsji37oVqGbX
1z5rvVeUBOMwY1e/VMHEmBsCqZhSSfR6bzSDK6edhKKyag7xVU+C0sHLKzjaXDwx+Bmpx1T5zUq4
Lps23V11duCG+NC3tdSFp8xQVNN/4MYCjbVdnx9+yuqJbTSEb1JcXHT9n25JCsztTIaBLLTYFGt6
1IWXvkoUi/eekFgwLOcj2KSEafm9OGN0aK0h4O5ND6k3hy1g1QgUXcZJtChvLlV89tzFtYiNzSx6
ARrszfihV2IqM1wHW66+U9rjttyWemCQa3jRrHny9WYBMhJY9nUm9vhlJ/HWR9Sfl7Wxl9baIhYe
N5ls5nmeR/2Y3xO6Je0rqH5ce9BgRMrOlMyHMEEGdfThVf5hL5c83fIjMSoWcj7ypjVPMgj1Psaa
E6Zx1hMDKW2t8GPE2nwjJykI7wxd/Ts1a6nE/8dlLrsEfWFC+ivWzXfP5S4Dc/4CRJDyR4aG8ZIT
+RI+yETyYS3lePtLRfUQVAbBT9BASP5DVzEE50ExpR+Q/kocrPKoY2fCKTPbUEJEpZFAHlVS15E/
jPS/Vacg1B17j9CeVOu4HPfx5iCk8+soOXky4bDOmfe+SBZq1G68DX4XfMAi4RmRPOViy9xHSG4M
NB9YIN9gSUD0V26uAWBymNPUxOjbIyVTb6u72TUIhfjc8rzCEEsH//6hsiIPqotErQkZ7uDCWfMx
MT4cbBiUgMtZZfS32IjkRjo907rGceaj35MwJWtabnPhi5YMMrLsR0IAKC6V/ahwk9xfto8FRrSN
RqrD+9JFMwHLbdXdk+Z4IW1LOp3bTl6+58nFGda4VHICIM1U+PAI60qktnkPHVVHOdqpQU+8WOHa
etl48r9G/LOxot2MH8iEFRvTX8Wm6yfxXFt9HYxT+/E7136tMiIr+ndrhlV1I4qovyimoGwcO34C
3Qk9Dmd5w3e31mEicSFdt/ex2Flrl8bAk5gkcgtOPFAKc33jd5FZzcsBBokZ/eH3cqZptt4vTO73
3dqy/wyFT4c70d8cxplFt/bIlWP5uHOxLpUuZl5l6qFnjvMet4q3Ognz7H498TzinyptGkZw62Q6
+W4vdlbeWOvqRHFctPwH1XNVKfSaghUhd9bXr+x6utG4hTH9FiQM6aDq7A59dwkn1QSROHfawyvW
0ldgDhmltK9BMmOq2QBMuka195aJNHYSeCj70aqwZsaYmxDsaKw6ZKc4BOF5XhBhlcSmC56tXivh
lNP7kGoswDaOvUzwxCtqvFmXj5BCVN0YDMsdoJz1waGhdAv82YJs/0b9OqGOSy+SqJ/SZBBbgOM/
PqFHnplvpgICASpLQcGnqVMROpNXAfuqbm5hg7icwjAgknTHctiXbaAgn4kA3q9WIvl6f6pEkMr9
nKSsb09/916M6m+Z81Itpq980U0PBAmV7LmCL2q57u7TMCEc/N7iPTWR3595MWCadrWyyeqBlOSW
4zF+3RzUtAN5UL+l301ADJ8JZazwndNiMUsox0/MjBRDzbt5x0BPHRZD8ovQzlheJhOGCwuAUz/M
F4HlEqV8riMUyiJ8A4SHp/2AX2seug65MYKDZVBrhGkoPsWsxm2XraET87aiDruWBLqn6eca5Eyk
NwLS/ekcybS+PgTo7Mh1xaX65ngo+FguGxv1buICTnSdNcwegi8A8G5X63wfAOLCAGArpfIbh/mt
bFoQQ/1M9aNQ9Rchq7cZVOV1QE7MM4W+DYpd/PQW9jf1a2YA0ViomDZ8bc308pJe0MqxAKTtGSOJ
KzF5FCQx7rqw+yrEX7m8Mvt1E854Au2vxm93JWly21egSzk2yhA4vrkdkyJkU3vlsTM02/LA4OCr
aG7X9Pm6ntM81nrvlJ3qLSmtXFHlB4BdY/cth+k2V+lQGHSOWQJ0klMHj7d6pNDemexE/Vlynded
CpQ3U17O5Ui5mENeNDmuCfZU3uYd1jfaBPqf80r6mXk0DlC5WDUsvRJatodV/ch0kpkQV9CWgM6j
8x0A9UqoQzLvOy8ZMlFtAXUEqebhYKd+OSEZaD+00w09UVMtg8P6qi/N4U8Dg20C9UaEzybnZv+I
IYLIlg6LjgCVIMmSkWuzRT+7xsgJninrJSwqtzaRuw1q1uE10b0sJdrBXJOjrv5oSAm3U1inHCQA
AW5xKO6m5pGzTBU8l0upjsLsHd4i7a3ZmvEwueun4ycsDxX1ZUgkOceZHLnzCjBGficgr3nyjCNz
RDqF2RAxar2dpPV6tcMrS0F8LWfqqjFzFyrWiA3CGHp7UWwubBwgexztHAMchiW5gq0c/XsIk9vJ
wX7QITJLfCAO+KMUF4mtzKuCGSmqshwkBXk7EXfNmf6dmJIl877JF2ptgZUr9GMG9qyGNUavz3M6
ZZ28FBIriA5cznelRqJJqMN8nhHbDyX18Da404awbgKKoGgwLDM3eQCbbAXegNugxbmS2J1ajJ9r
NvQq/0huBh4OTPX6TG6W4Mio18Hn+kW/pxP+ExC9JbkB0X4EbXNoHpxBMLX2NRF28/T3cf0AcXpw
LJMFUgDKbNLopoGc1O6WX+BdG/fOy3oNmsM/u90srE7sTHkDeF+7b0OardHSXv8iIBnceM9/Gott
ljpMpAi8cJ1ct3b0MgF1CWY3xtSI4wlk8WdHrDNh8kiLbjDuAawpnTARpQNINewpgO6Z7568j/ja
1l6l6LZc/MNl8U40G6W2N+MNWTZaefzXrnAugFTXveVK3sy3IecTV+kthQAqmPnrNBytao4Pd0sf
JD1JeSc5j5jiyFBWy+H127nzRybaaLBL/9qjAlm6C4+v/Iwx45EzeM+4r8xBAU+8zbIKbAeP8+TA
98AHGTa/7Nrw/3PcGvwP+qxV5qzt0zcLEDGgrq/fqUjluVVd2XF1EMMld0dz7ScKN1kMm4E78miZ
OU8t1dqG1TVM7Wt2Jn2HlQxPSc377ujVde5mo4gQBEjJ6lC600q0xuExT91qJ29f17eHUQfZuLO1
Lm6eARC6AJLBdCnbW/l4zFNy2K8B3O/vGwCPNs8Aag4EEjpFjcUxKqYmj/lCvAXcrdxkfdpQlvoa
F49d/YGvFQaEjW+IJzD58Lz5is4I1C9dW9sd6E5581R3CYZDc8LrnO/0SkPe0UdM5viN0HsbnP54
nJyhqC69m2lEYoj3N6N648n5oqJhLKfLK9vzWnzWNhn+AzKKd+XJzYrInrOtuVhS3o7HDhhpSC9y
/lfDbyCXO7qGQLovkOBX
`protect end_protected
