-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lflvdr67nob28sSL0x0bWpNl7MuydevtFCBBUezd0mDKBnmsXJq8JLMt4HqqJIKDZ6Fvq/mz06e6
bvkRaSta8QdLfgTwRxDMNwEbzEkK/3GFt7nlu/vsrP3B7jWqUxGp3DXiI22pWAyNWJwKchOcw7a+
AzWQYBpUMkW+yi0nwnRyByS6UqvGnuaPc/T3TP2sRgf94P3v8Cj401KhjF6bS4N14oWFlZwwBRqy
Uy3tig05CGzefRozdw1Z5y4UmnXOtyDzVyN/K3lAsml1/b9kP16tljJqOCBVJ8AOrBgx6ZnqU7fN
wsZbs8ha7F82xHBnIIOOA8HZePk1c2VE7mRWOg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
4O89mgm+TUp1C9fet2SMwfZ5f5q6y6RB162f0exwtJ8H5xZ+5YaYdq27RtxBljVO5SB5dmDYjXZD
Amk69qSL+iQmT6mLFBb1JvOwqwqcgWMwgh0e/uZeta3sOQapnTwSVG5BKclssFvamlMNLQsyruUl
ejd+1o2r/1tZq/81d2cl6bDS0BV+QeN/U3ktp/wqm1FymDiN/sxwsMaL24Bo5bzpbbS9gJRW+1qG
86YfxQigNGsz4mruMvBHqrQQO2u3lMBzjJyBzsEjGPp0qEzgrzT0i1N9F2Zl22jDV9NQ27yRbMKB
wMBI8XmFZWX6wR6XFAV9MrjXKQ0vqTo6BTTzPfgOOS6ZsEkKmp1CZpHpewvI7uxeKej2LvycQNs7
VbOc7DZYFpUb21pmmCRnd8wGjicwQdVJoHsBqBPVChoXiaR1XjpFaZfeXczhpvUZPHiM37pE5Vze
swOSl9sEueSyqKk0hty+/zU8GqcrSfXZ/CTzaQFO0glVl/Xbww/gfHb5OhiB0ibEo35RPs5LfsfK
+0OJwCUHArAcr0/PRiljzeaL70G4fNzlyIOSR+7E/aL06lj5RUTNdtSKqzRbZGfBIxBZraFPP3Xp
KzRJ/JPu94HtcUrJ2TfWJ15/Tq+ysBI1tNHRLNZTSeTXQv9B9nLbd6w+VAStubwcBMNVwCfiA9co
gYikV8yJ5Cv5fQTmeHEvYmENbBGBHz9en/nEjSlvYZLtHx8oiAWe+ZmdlyPRGmfcL3CaTlfa3nT4
2eM0jia1qUhSoo8hEkk6a6P9aI9ZVjEXoyLWeu5PkGE3TothhmYUzWOu/xaj/7wn3LvP4DgoKIOd
8abQG+vGVOdcca8iuXoXoepU5B1P3mOjBvtUdLIvjqRhu1JRcYadpb9dupnaC2BTo0RSWpup2mO8
BhDu8GPHC2lMKhPZrbAtw2M3E0ZTBycwjVOuRo1E+ntra4i41Wyo878Rh5n2+iYaXuE9cOEOcbLA
W3qvzjUwj10GqUrJ0Zf87I0s1Ig39/X1w1zFIP+t/RWkPSbumnZMLaSTTKcetZwJKDr9ZTC0hVP2
UY0VAwUbRbvkRAL2gLRsi4fI0nm0eKtKQd2xNAv+lM/afozAUaMwZITPALgfZ/rVnwH/4o9jjV4B
QbNmV3or1Hg097quHzQWuyWbvfjS6u9ZEhL4nvc1yqdsXghVVZvUmimyV1ALjzPp3ADWlCjZwzEY
2B3ZZkJmRmO9ai5qdkrP1dtkcoxOvuFI5dGR3LvkDDFrGm1ms+DfzWxsEVyaFhX1HDeL6WR7FORr
yweL0ZYx7eecomI78EsPba9+zV2vbtRqdQOVntcgBD+gSMgZW445vnkZ4hK9eMX3KIPrHyCGVPtA
SE7h+ToNep1Fa0Hz5maIOpSNpldjFWwV1rVUOSkHmlS3CrbI4VHP2oijXwCMIyvZC9foHeY0HWQj
1zZ3+h7X26K+6qQ7gytvB0XsZbbNz1TftAQrDKcgHhMa7RZsoHnUPZQNOLPT9e90ifM9XLA9HWU4
4BP8MM3/jPd9xROLy9O+5nHbQZTcNr8n/U8FwOXirlNQcTjylB/ig89Es+GMRUv0glYQ+AIqUxl1
C8Q1wsXV4VRfsiuW1zjpVcQIBNGQQUS0G84IMb/3Xrd+tOxH4dao1rIC50HJzS1BI1nK7ffkhefK
BI06cRlyipeXZ3QDSDCt61gllBByLXkqkEjv5uynBibKY8KfAPmDWL7QEvPidqMKM744ncOh5+fJ
+wwKnu+GtUXN38GePLoEiUdyKC3Q5OFadjqAa1CcsqZeVHgP7XLKlRSVfRWAZUMfy+S9OAxeHt+U
P9KuS0C+Gh/53IOC8rk9+0sv+WOD70K3Dpxn4NW5U6W6xPgMMEtCeOX1d0n8WdUwB8f2rQjLeXTx
cGnJqfI5l6IUVFvYzi8j3K4LzgcTSLsXoeUXwf8X4oajmwW/6GkuwGXXR5WnDwy0Zvpyd+QivTKy
QcUUCNqW34tJt1ps9ry55Sa3mm0nWrPzhB+vc64i8qTjBJdgkmFcoIxUM5vJGSDiu7c6Q+DhAJsH
as5i5QnOrkOA5hk9sskqk/27N6H5Wmz7Q0AM90BCU2cninNCSaD8p3O+3iNBPRdcWvrI/cA1FMff
ffq7HWLsr1EFaHcZfVFlSyQUvvf+sVVFOLqwoyYNQQg31tomCLCwLXy2SnYxv963gLz8yrB+ZhNE
VDhg+kxBsF7B1hI+ccMYhj4BfsS4rbg1uZhZ/rVXas4xtq9I6UPemYjnTpuhoC/ATCRP8jEWvahf
AsSrd3U3J7/gWEkgXWDYy1XIuiuLacvuiQSJYQcqsnjdiIMkiLu/jrr0hgfPQi0nmEq5tn6lPFen
Hrc/444bSedtQCfQ/f12Erb88Onj+rUJhtzAjNQWpZxcUn4W8FZ01Fcu1lfmn2alv0nqnUo4FTgb
7aLI6fCyrxrR32ULtUhKsPBvD/N/84MT8AUmHEFAuFWLnSz4j7TSQayLgY7dxpTLl4Xn7JskvEOY
FeIUohyvz2jkkJCrvUozLOX0FlG6DeuNel23opd8LSR4j+7yOr+Xhja4XXRnlrIOlR22YzASLh9n
kspS2afnz3yovHK0fu1jdWxJ/TdHRwCvnL+8Ya6tOjvTr2rR5WZLkfcj/Mr4VOBvQz6KWqbuJiRU
5fPkFrqIrdPR9HQ7DJewaY/aongD0w+tRpRqtKv8HhrdOoxCcICBjrMONtTAqHx+1s3owTp1ZsHQ
shEUAk6QqhUpmT26bmvE37pZJGeHD1DU6Prl/eyHibm+kIlo8rUWzysYPdWz6d+BgJdbGQhF84Hu
E4hWTjRBveHhVFEZg9haWwDL7EfKxQvqcAnuBZF+w/yJVRpBG1szz0qb5AH4h0VVWmyxqiYZF3mJ
x28PylfQjjOQrzfXhwZpojtMvBhS+1S67oVi3fgBAFGWsLc3EUGxmyWzzO49NCuf15sHglbCJHCY
pto2he4pivAmc/wT9inFa1ZtuAkzGl9FSpUzZBPo0dOx4h+WPPg5iMpMUynlG6ly7oCy2tXVLv67
JXfDBN3zeg6lQsZnUv3C/RVFjSOFLYJ1FYa/a1Ac4ehDI/0/lKp+vTdn6lIxqI6l09kLpvIXX/fr
zrZ5f/rTS+5s4tVVhQHCrkG60OdXdF6pO4MLXO19OXKKtt6Xnxm/sFvGkS2aIX4Sd55CdRuwP2V7
cIRkQypeJhbGUR1mIX3fOTgk8jTnRWLU202r0OUH9YzXsASZamh8P4+oQ/sqoq3vLkpr4Fw4Hem0
BuusC1yb5pX9vcg7eZi0w1wgA9N6vr31jqgn5y6dc1n2dRkevA2O22nOxKDU8yIw7VfilN+eW72x
dKbgcBd7ILp6Q21CAPRq+jrAj/NrMUyKYC4QXGdRVNZsjHwW0XuLKWn+DrOB8EZieZNqRetuqRQ6
RuogJIEbtbc2HnPr8Run369gzBh6foA4KTfU4VdBj0Yeq1jsxL2eKGMu5QSdD8i5eI7QvoFEqX/x
AJfYFRiIg6xn2WwqvzpuFcwE2njTkQhAWvcFlHstxix/dMcN8jP6+VsIDfJtizihYZhzyyTXm3i/
YwUnllSw7kCC8ZP7z/xQA5g+06FBO06J0d/b6Lp6eJ1xtoj1zwBeERPmZdqgTQB1vxkz3P/dObj5
l/G60rfgGxdLRDtGgw5WXUwrS3Ksd5yQ6FMDAA0LL36hFR1cKm1SvaoJZ6xvvDWEA0hyPY8Q1K3K
2nwSd8G8VAbxdz/kGFHUeY0npknRoMCEWoGJT0hVlYYHWjozMGQVG7jJKvM6Vmxg5tkR2SZk5aLB
CqswfB3VORzdhysE+dX15Lpkyx3oBhJUgMCtqGzs2HnK5bed4n+ok8r7RyWIz7wyfNfoX3BwXpxL
1zazWyvZwyNVlsCBLViL4CfjCB2Pg6ei68DBVsp41G9L3+gBbSPcp5XFp0WrpQe9iQYnaMF6Kgrb
LE5hGkaEg6MNUO4jzmtA767IihVAnskvLHBrbSr/jkNJ+hAEMxntirBYEmhfW0kr+9ljIUjLwd5m
SxsTk+tW8fS/GL4NaGUTeF0hGSTBOLmCASwxfzfYAaUEVza2RCVNDp1ALAeTQIJDtIS7MwXIr382
shTW1o6pxbTgutZ4/hgRokq08uX5Nsk7S/D1D04wGk1PDkTwIn47Y2NSWtiG7jkmX9jt2Q45UlYv
tHpZeJiXwQc5jl62tdhcQPstQxuSmFlhEsPhtizclX6YVdTlFlpL0oiR5feu5Sd/lYKK4qkk1++8
SQCVkaFIX9mCgMouEWgHLnPC+D+CYF3AtEndZz2xum3XTInVKCjeuPpigplOX7Dkhkd34ff4aTCX
PprIQxqELg03QnqkvmguAht7i5Tkjok2Cyz/uVKEw7IAiAowYWTKLv8pCWwVhn4QsxVCmzgq4Uzx
09XglQS7lEWfANacWJpeUK/7dnwRFdbSUGRgEyb5O1Rdm3utOkeGPL6eJTbZQuw/uw3m7TdQi2SF
8lu69yzEr9FRkiMsrzznjh8KrBsOYn3ZEi1ex9sJLaoWDSQIshsIjWqlIUdDwLVTruZnN5/UIg+x
g8KkIjbK1W4LXmlRten1a/14TkEhRUZ1eDeuBZwqHkUalSjaf3I48yRPi4PZgBrq6EkslyRwiBBP
ZBqlZecQNOcR5WZLSVyTCqGt0UJEZemsbamkqZEMKvadznrm7QXveApjyHhHd7OYRfpwrgJRmo/X
1ywSLbAan6LOA6ERvORTAuHGF8il9nwNAsgMj+u4Ti23fdTDWxEwUyxYCnR+/0KOTyohm0To8opL
KuLN0oc1nbPMkWavqQ+lw5JINoPy9BIeVO4bv8xho+589xIlIm+puW/y9R/iKz2VAFgUYWaRsUzy
QjBv7l9lKgDJJipfcr4yGB+BSwxQOKvEBqiYe6MdnXjT8HuKaOYSDh17m1nIqRf664KjhF7/jrxN
nUGyS25Nm5R63FtFQPFgJlSrjb5TrdhUdyHcB7sY0W9TbogfBE6YorIhrvU5EW68rVZydrRqyqUk
RrPv9fPswu1osHX+H2M95j/5FAz+WnWL6HtdNB1j8UanenIosFNLxTsj8gW3Wb5wd9tFpfXcdJ8k
fbGpDv5t42da0WMu5vAdqAVsWlVvdDpfH/Lta0KMehJeq8rsFE1odqpotj3GEBduimYu5F5onfxb
brNXWjM3PKBQwKBLHMxbqzeHdnHFOvFPyfoafBwtRUG9g+2+a5k4qXczFzC+7n/xRFfA1DD1UbWX
LsYiQINLE7L+M3vCbRpG+rd+4ms18OfH3/FojbLbiI89IsO+hr2SWLS1VwoAuti/W5Pe8pVlg66R
lxLoS1nWL99KFfIDLzkLCjuv3bA739Ymh0kMYp0VGuvcNphmWAJ2s/SSCxejWAkX4RCFFJIOq/Kd
jPQ+qiuI7chdPGflRrtV+6w3cwnRw5BNf7vU+ZgChsSRC+3/xctMveX+UK8mg/6QyZZOJKO+9Znk
JAcZGGs+RsPzUuErYxNy8+beqhDj0pW1rKpp5VkLMbyglQX551m6VYDxF7RFzF6B6+djcLAvYtkG
QkSVLxtCJhfVeiBopiGYdw5s0jUJKVpA2eE5LkhYNfVRbwUEM/Ch80SxA7PRsJpaDxDw6Q7rCEjs
6HdC5U+e9ziNsUu8tRA7E1N/CQNN/36Ya2u/rqKpuYE0bMLBqlpi9iH8xqPMjzW7ddS7H43hHb4O
mqtenIUVHJA4haCCN0iBl399MTpdbITc7AhMI2EX+Jw7L3FCYdsFjWpGWdrdLGIC9/TWpRflUZvG
ESWAwTQPBFoCeDZi79wXWy39frRuesBCFIgYnopqIkP5qeY9LcPu3zKiX4DW5/YvRSuig4SL6df0
GyOq0D0TUH8Ra5gyYiMl0JTGv/P/fVl+2peUbYP5OrswbVOPece6b8ogZeERVQaKlZUvbTVAUwDa
ujcosN6UHOM0XhHEVHMvEpFj3bGHLlGQhof0L3kdT+NLDtJVJI8A3LDeLfKeiH2urMgzh/2pS1Ad
yrBFSnfh/jqRNY5e8x1aUtobytXlTngqi817Mq3nT1URXlXvQ8jrccLFsupFOFEpKbMkuEDUvTR/
aD/wdXI0CG4+VZcqo+7/tvbvpCScOHy+vIE6GHebzKeysGrXP5mzXddW+ZXeaij51P/8wgwqyygA
Ps+/zCexf8BRXZocPFjiF4UNfmZQeBR0JVPii3GcIxypxYUNxmDIR6zrB+gOqs0tTw/lh0FnAYla
F/TXyODSjM50Jh9r1rqGpDA7uX3cAzxS3p8m0S4vt5PhzdgXC0tGQLzODKeJkc8ShvCEGT5qSPN8
50hI0MAiusOeiycKCWuFbaK18kEBp/izZhsfGm6t926Zowi+Bd6tV9KjIcFDB/v9qnwdvBm2HKuF
jDQpC51AtocJ6U2FxVXkkQ27ZIHBbWB7Dr8DwGBAjteJLp1r13Gs8Cwu77g4r4qytT10Grh7lYym
90lnspBAosqz+7859VEm3vL+XDKJgBl28oLviCmsmW/FyN48OHm+OZZgaAvkdu/ni0ulUVaxFpM4
ImUP74HpKJ1SeSzoPm018r3fkb4ntRTM5vbew8D4miJfIkO/gdZSw6r7LtjRiF1J78GZi1PgK38X
byQg0Fbk97nsGQ19EC+D34Bm4Pvd2k8NOlMbIDNhBaearqYO5ZMhLHrWu85kHMormPcOuVhoR7aw
ZOttAQeXmRtHYBS2Eranw2/EOJylh+XqpTp/aaJIT0xCDglgpzhCm4mJFBb6kYWF6ASqpWmCav1J
0cKQ++Jvgq2AxLOva7t33WiBHxRmyxE/XWa9lgC5q4nNKbgm4XR87FFeISC6U9QlMl++Iikx8lSN
AtvJ4jIRVhY1YbfEhhW2RMVja0i/v1HfUsDC2gX2v3sFhbi2wANRzC/SiVGWT7RaCg9R0LTIoV7+
NiSEjxoQGyxEq+CSt9gm+z5ShdhfPo25N85TiVemL0ldHHVOqbC+tzs8Obk7kooEy2hZ0Cm7DpGJ
dvw7yEqeFFOMPHTOhtmWfttCGMnPrLdUYjw6eQMSnJQiu+TZ3B0q0+HXnKVl77GOX9GnlmZNJCX6
Sun2gTm3/ZuZnZR7gSmH8Hu3nKa0OIMFZHNVp5DC2KIBlRJzzVfQGxME8+dbSm/vBY1kiAZy37uG
6beh/BT8CXWknkJ1O4uI/i2gn58ZCT5v6FzQqimoowrWCd60GLLTTKdOEkXOnKNg15gY6iL+xmP5
q6JQN2jZuA3TUraGx1UMvS3pmx7TBxuhBPj6LFOkj5hUcNzw415jdBihE0gvWobEMw7Lam+4uBTg
2t7AfzbRq4Ul94o9m+ri/CMrpSy/lyzKAOMyQrtrFFmHvPVNBTZV9M9X4auXGsWhBBpcEgDJHick
WY4fnBaH6eUIh86cIYUhGPpf8CImAoyf40JRopeqyTgtP9Z6hjxbz2N6T3PIISbzcIpJ0dRBVkSu
j4rSPnzVc8OnF26Uxxgd8Jo/Vw0+c1+wl7umsc40jyG5CGvPJuGuqfB/PKdqxS3y6bGw8VHdCZUV
d8rlKWMnlx/d558rLPxehMm69xBeTbI/bz3lZfYLWJeRtTM8NC0wBMD4aKimTrrf/LM+4YNEljlN
V0qyp9YOES//dcy+B8wM6KpOYYOo7wbCxZV6bAJMAYwwFgkng6nMvlrRGoew37AFmLxzU1lxmn5z
aiJxGROjzvwxtb1ry0iuV4Q7pGYYFIN/Qh3Oqfz7s6U2nSmKQh5sCumtKur1PJM/Df2Ou0Z8suCr
JKu9cbt8BRZoE8BKFmdgpbf7PDvHQdJIiYrXWfniVoAaucCFzayj0hKQQzgl5ss0fLFo/Ud+hfKG
uwXGhV6XF9HySS5BXV3K2d0cNEYWvbZv2vSIksFaisEUcvPyOz2wOlH11QjKkLr8vRk0PknE3akn
LEGd3waX4ESN8Y9nqwPFSZqV4jS3cqap371dZb+mFQmbObtYDbooCUczR36pZG5YM6GX9iGchyuK
Pmj5yJn1Jk1yIpea77EYr8aGmEEB1tAmG7otRRFni+bPK3EtfIat/udo+RuSdssfQRzwLUIrzMqT
sTKkrgozN6yjF8Az0mytwbK9eNFDgHSdsgbH1dPb47nkIeIMk7kvpXfL0ydb7LaPsxjC6S7xgcu4
vdJgv3/OocAagZvaHZcHnsSGUIZ2gmZKozO44N7XrFHuLJtTD/VEwceQ3Ke/7r50KXaGtyJIrhSX
LZnSqxNN9GTf+8UvEk/bZuJy6YenvUHkNE16wyVV0F682DP6lGy6iHPN5IHAamvhgbOOvCSjcBQB
dOFaUjWGiUYTJ9vbySTsrxLku3MTd7AvB4FSFyaiQ5oxPQOrzTPsrs+NPJtl9OxIHqNg6cPTvPZw
3+sXImFxJuovTgnchCNchHKQ+JJUHRPSXfhfIML/iy1ttF1Wxl+2QETez/TUNpQyIqbSsg12803A
KT17rjzjths1AGoz9K03tC+HbqwuZMs/Axb8xRbL87PzXdRCY4zwCQ7SrqjwEqYaRuy60L3opx/6
J9htPCJDIBDqPtYw5z3i9u6MHR1KyAP6JY+C+/MU1oIVviKiiQ0nQxDbbC0ukmYolyiAx1FwHgOi
M17t8yaHQ4tshZy7vA7FA0Nv3hPu3Dpaozw2HldKGjIg4Xzv64I8M8RrayvqGuSOuuB0rQgBnxhw
1/OKF1c+c19xn6phITwb+kQVNB6fTnKLKAN7i1Vw9Awmbm0jzVjBhc8lWyD48UmtesEc8CR7HpXR
9QnoORz/DDS1+HFfTCgpbTw2V2iLHJrYFFKGTI93GWgZsa6qcxEvZwh6yYIvKfBDLQly9alXdXUF
sCa30N2HoPnY7b0b6hwRxYGjINFqV8+K1uLEfYHBTE9uvUxYSpGA5KQenyUM1rp9x5KMxGmK5Ln9
t/lLLJ192zAQRuLb19EwDPK20j8ccCqs1Xut/F6c7VTlK5IuGG1yEEWzz6RhfKFNZWHHTNwBiuIx
5RzibSa8pU3XLwKT+fQPjhp87UH1llSIyAy0w1F0PIZG+UDZheAzc+Z70OjuuXrhDQS4pjbovA7s
4rfv3r54t4RbCmzeknZmIFkjgHo8kyCcZZ7aKwAh3zAAzlNkm5FQut5Me+EKYtceavu3T9csyrAX
IWkvEOB9o2eD3v8tKtbNgIYOuAbwWboklNCJ/Mi54aAgGT1zEB/cxW49xw/cBB3BI1RBcvha1jwa
RHYeNjUMR6hXQP4Xm85I9qLYc19/ca8RgO2ksm+izG6TOx4fyOiNJ/GwBVLNPNN32RS3Ka8hgw1M
+yRAEWyQghkY3jjL5MEqAPfd/hOTtY0LNfgZwpKn7ZstMWBdYvk61PXCwGfPdDgGONb6L7boprTW
cqmEctFO5zIZUi7CrPi55GBnJnJvEPLuUy+3bhlyutLk4WXH7KUzsRVmLv4tX9b63A45Xo+8vfNH
53z6GtN2U522vU3rbO/P7e6RVilyjIEvYF64zOqS/XmIuNiyoAo2WFYhgcpYid7aK/k3iaBzk8rf
ulxWDyXTYaj1REzzMHCpCFSHzdFz3tgb8+D4NQRvKpUmXBA/BFkM5H3ZEa9DBzemsgo9bozbCY3D
cbkaxXCyLroc4vYm0Lzu/cLQyyhoJ5CmeE6NQqj/lDw9+50Q5SLRQgveIF3fzsQAEqqvBqhZJo+4
koWSt4WQIQmh0SkPZ3AAZWxT70PDhM2wBtwKrwFem7BSdUVLqhPZSU/IAm+5BYVfp8q+08aJJogN
05Cr5cRkBXCLdm2x66TuVzRgztAps2mOdSKW22XZWAyeaGRSj0q2ZggUCD/TUyk4VVR3Ry0BhMi/
QKlFldX4h8kGzS4JvdzaPxlYgKIDOfMJBJkfbIbUmWQR9AN7iNOBrC73USB2Id35gssavagq9l8G
hWNOhH56oaSo6qSnWMK+giwB812pgOar5kefswxUSfcFaxmxKTwPXbMPE5eetgjViMGRAtY4lhF3
WrN+ZFPqaZoFfNMkaqTJdXfpYKlrAWdDzfW3SEsN+N732ocXYsWtcZycoNqTnTqg6jKQ5fMIwMrB
sRAuE8w0lbans9HJcpwnh6Knji4I9hMmXiXaJ2RhFPufYdOd6LlqSl7Pixkpe6UYI8WkvRguH1mo
KemIsnG3zbhVDdr26+Pmj8IKOifuSHlTkUjuYdjV2k8fh4042hQ6aGG1PEORsgL/ec2QFlhPI8Ou
++ETPaO7NpxQpLBFCR2SfbyvBt+BW6U8uZc3nafY6LwaM+mdVeFRYC/1UU5+u2aSyMIqbaLTwwOj
WfKgTwvGND1R1m7qeWbyeePlBCQHgLmIu+GpYlv7sTRj5O3L3ouo1M8h2fD5n9YFldvayBbcJnh/
GM/eSQxw10k2L1L09BUyWQC0HOIAdmn/kRnpe/v7CRhPfuZ4OWlHbzEF2LpRdTjZvtUGdUaax5wa
DRso0Ds/u8TERwUfY2XK+O6Bly2EHCJxibXg6ZPJ1aQECnZ5ql5QpUIYI7bJKJSuIcZyZuQfsx/L
e2FFtmUdBOGylwOfg9wlx2iy7ndilzDf2k9yur+5DTTtn/99rnMyo4euq0SrqSI2Ngtp6bWYvJWx
xcFu1yf2OhqQUYY6DkgD/lsK0w/Im/CBJHn+l3FU4/p0cRiw5p92JVnwhz+yk3j94Bu/UzkrObt9
gwg+MJYUm3Ps6kGNDaqUY5BMwBlcUB99swLIydUTxbZmZjcLydELtwCK6E1eJ9erkeFBKzRv6rgT
k1nPffrki+eWDytjJdvE9KqA0v67hmtNYxq+8sjibu04WmbbbvVw6K+D78BJuCnzYAuiuTARZ/4x
Ddk9pwj6HO4PrSAEaA4N+47l8/3Ye4JXpeuHgVodkug8D33c0W+9bM8ujFL5lNjHA503sRxpX+Hw
mcq8XJxjiFwM+F8E5lokW0GrucK1lQTxKYPgDAIU/gzU8r+4Pr8UfUZksc6OJJ+E/j3YB6ohlne+
tRhJQIPv9Ymx2xjhzpMjfHrmepwh984XtCNkEn43hFHlUgOsrgUpZ/0iByrt+4q2iCNv7Y6RmKaz
t+X58oJC5oHHm54M+Kr6wY9m+5fNk9H7KymCPgAewHohlDUqaElvp4QJ4GED6VrSlajz9h30GiOX
fAI/+QpDRE1P0IgrAzVl+jEhGP177o0uE/BQoYSxKLVo7J0EItRPhhhr89KCUJCen012HUqZ3a3p
yn71bRFiRlxahahvtWoz2kMYl97Gj0/NeiuWy0uJRmU2f/5oGnQe+Ux/kVM5Cd0lPDlw3+Pm3wTo
u80VF9iGOFUGeJVLHvebHlnopGaBGWtS9RxI6PG9AOF7KhducM0xjW+Uz8TN3Xrr/fUchxvtrFNC
gNzulh0KDYeG4XtohBs9UDAAle70I8+u1REkRDjnfHBnoe7QdrlsyY2RRiGyv73iC5JmfG771UH/
qHusXjB4aSuHul1+iKbWwEDcNYeLS2xP6F43mr+vVb1Oc947ywKiQTywzJYpkhMiO1BEk159NUpq
FFz9z9k6zGPIczU3bQiULjId4pmss9/O1gL3kLABY/3Cf1oBF3Kwgdl2d7I3zEpZoarpVUIq2kpH
AQP9X1EAO1ijAg0TJ04kysV8wZilnt8r5p8QgnT4LbzB9QvFcGdqeMAkrisC3neMxJICmVhkKICw
wuv5uiajNqfVC4ylcO1syUZYZTvFmDcUQqM57uk9aT9Fmu4bfQmTsusJMCLdTBWSxg8IyQkfpvoG
pokRI78imDcIsfuesE2gazBrUMB8vSVeLfGrOJI/BMTgdJmWTQ+GkVr8GM96fzAFQsVIq4KzQjYL
+C/HM6tbp387EmEdpd3HxXIM4Sgtwa/dfPDOhdDqz1EUGIxg02E312or+/Ru6Lx+a/uUH0p6MdA2
0/t8Slfjg57jLC3vYwHCabkqpevmmhMmoQKKmbl4MoaUUWmm+6da4ZGdiUjwmYSXrowLd1LFIA3p
XMWBHQ/Lqih+PW5O6/N3cyAAtasgHvm4++Vqs7lcOjlbDIXuy+pe3Nv3hK33yNSjAZQ8eedP6dqd
NBSYqgmugbtaeUMuK5ZgRwdKs4YXK2F2lGeBfx9xr1nfmmQj1S574BSKrFU/BC+3RnRu0KV1srt3
3Uip7eOYxlOhcQ+e2RJfcn4KX8LP3NWITdvKR1Hz+FZ7OKBKKoviDhLx1/Xdu/iprvK75QsHnLET
rAjya54bnPaLQqc41pLZpwvdepvdrGZGG8OOnMYUM8k5k4FVm6JcWLuaIL0KvUGSN58ZgZDvJXEx
ttlcifBxDLfHUjFtltz1FhG4wcmjutMUOyH0TubDUqFUdPEKA4lhr3YQIlkUNPVy2gGQihNqFuFt
SdmO3uLmJeeb09RwdIOkDVVOaqKGWpt1bYkB6KUZ7lDlNPmAFnG2b02R+yYeX+fadd81gA5OuUX1
u/8wtbSOj54zxXclXD0ptF3hoND5px5MaU+46jOu2MPaVfosqSyX+7BWrjiP7xKzwSyJm1Czi+Cg
0EDNBJGDbeSdFrg7mQkdCQsfmsaWR2+1gwXCb//vC8368vrNk3n5qVk2PabzreqBLQV9sIRUYf9x
LSLc4KAL7xl0fl+ZWdHJOYWFP3WskZZnlsQAgd/5UBVcNJN333iihAPGHp/D2D3mAEyassI1cJx6
o6lj7+Wk1p3zebC2N8BlmOVCvc42pJtJ0RgxehscIayX/6G9tFiPcJl/L1q49Nbzp5tg4eD50XTn
M9FDJv4suY0GeB2+8eY4XtyIXVeeoWnZMjMX4HbiLqqvQtdfR1ms9xPkKjw3/aUIAVYRKX+ZveWz
NEWnjKPrXIYANeo01m1Gi3jIyuv/73XNSS1zz4cSzJHBe9xOjGn3ZunCbanPvDhbxTonMpolrYnx
bZ6781ZQ3R3ucokmEt135QFeG4+ZJdrqJbNwn3VsnE31Rym6/LBHUWSi8jVkkUxNjC5GOeqbxxG6
qCJgr/2WKET92kRyn5DIkPurA+df00WqGCWsheTHUdgB73jwkr9frtpA+R2XCiZSDPamVOrgLHqv
POdfZaaE1v3cAcK8nlL6aeLHXcRBOMg7QVxxGRFa3zV0us/pHHCEVMpSw4I43GkJ+sLQGcBV+O4W
zAIf0tAVozwNX+YfF/TzOC6PN+Svz7CrtWi0rpJn5aDGXJKZExJMm8uQEVexIOQozkNGzlzxOPOS
XlrsbYKfSu35y840opxPGfGfENCDYrus5beZd6GR0lrPIuo+3gzkPlNDWzaX2c3C8lNj3msJd+w8
poZGACD8J7jyxzenhkxdp2Va4Xg0pfcvFmmhuiRTc+J0SQEO++RIC7wRVM0XtQvtndFQ0IKb/wQx
Wylxt9cy8Hx/PXfH7iMJxHiSma+W0Ww8oPhfH/9UeVIJD97nZFsPAMDGoYlJiYryQ34HnM2HzTBw
JTRpXVqG4tESG+3UQsSywXQvlljLFNCHulle1Ln0qRE7Bap6KqRpLFM6/kxBmkIsQ+b3YOwyYANC
MVK1ltRQz1xymz154UxeIValMKroA0VlyCqp2tt6rF0uIbg9B+4masixJne3c1gGvtkJkJHUk0XF
m7gAXRNw3htbXKuh2Sn2ZUuyDjABxntsTzmFeCv2oB5HCEVYqGVUxJi38giPk/qgx+qVWt8+itaf
5t2SJ6rlSTV95HbNEbdKjly8NlzYhhS6hKlrg4hi1NM6U/8dSJ62XNapFr22eXlbXosis7c1xhC0
5rgGFWOlcoKd3WJ5EezGWEXqIA860WrLq4ttUC/sEpLq/ddo2OQUirowNxaxJvso9H6om4jDIG4N
LXqozOfqMk2wccudSDmyEj10HNuBrJ/811kVZPrgXS4ChTHobWjBFf8/VkBqpIihqVMfaSpjjZ7Q
Kkl34H3ynu35SBOf51NmgHva5Bgq+8r4+9JRNKpx3OA816ZmIvtJPb5kw+dZt128fw/ccG5FlvVJ
1SIrYS7A+mnod/Baq/klyXxcxMpuER/dbvP+eyJ/EoeifiDUj75GKsFIUZDlbDnJqVxKlGhOWZcy
RQO5TqmP1QEndDl60141SWUeKWxdYdxIMSEfSVkDF+/N/etNKA+Y2JRwrjPoKIAX6MBxgZYTfrLg
X3CvgJtiQGhvJ9RsRgbMMkQDCCB1gKtAb0acHV+y/cNFUh3dW/QJzCaAiUNyaFiw2yX6s0+MBtIy
sZNif7YlQxVF20v1UH06nw63dDTssSnpTMSWlvgjrO2GB9qHyAu0Qva6ZODWgvsThSiPq33LYApg
46MNj4K/qH82VWu8ZZOUyIN1jGXBwW83NWptK4YMIFIIGBwI4S+Gu+9UyU7cUZtq9o41lDmTnBX/
ZiPCh2tjJl92lDZcrRBzRaRcFXJtixXNmDsj4qkHmCV6f0FwMPug8SKwLwU4zSL4f+ENszp3e5Vs
6Rhn+19pwsBqj96Bm9/osN5mOVkmOB3xV67gd+CUP+z5AhqpFnkTMyl/SucuZbE72O4gfcbg9CZs
4vk25XWloRYw9TDU+A4hBuZ31DJLnOX/8zEkH1FCOgsbgP2ym8uWZK4YOzv2DN8D0UfmCFTY+8HU
QLO59MF/IFADTfZ+iP9lIBmdT/SlihFuBSSxfp6ciKBJXzrB+pGWM7raf7g9K/g0YVyhThK6QgGi
76aR1Y3fBTJ4GXhNAWmxtrInEexTj2we7x55/HIeyTWSQRCoDiz6eB58IYUlUi0luQ6QZDlHhEQU
6JYn6tNnmE8i+ehZZF0OEdA/wgFVHOkuUZMVWvV1tLxAWNzOLImxswfE9CejN3xRobIqWN4+/mHw
ErYJ8N9vRwEvoBbvMbmBr6HO6Zd1KMIY8jtP5FHezL4fohxLTgu4+GjUaVaIBGZRCABSEDxKYTua
7bziXB6W2R6GoeddUX+FoYhATra78fqXU7xe+8KemyGBIChsgr6zx5KQyp4RVMT2N3cjbXNcIzHx
pGuh1aDBgnsxKqG26ZMGAMyAN6fXZ8UXm/Rbgfk0HnXd65veIJs3gQ/MBBFtHBsXuvPhXvd7Azzg
zUQbqLnhrDsf8rXoRrVhRYkwwb7IO2yLIGOxO7+OgnsQSq0axukEb4AVhHpbPPpcakT5VoD7thkO
1ynUiRkf6uO1L3ZAG+cUgtc+mM0h/627waOhaC5BjBi5ibBWeRTkuKSDetiU3oF6Vff2Pk5z49co
Sg9Ijzi6R2sPpKmaWriRE5LeJTAo09Eaej9HcmGMqL+sNHs65W/aI2BhQyMB+2CoxGfAu0f1PYrp
5uvUZom2tOpXmkMQabw6JI0FwYNG4vcYBAWsOe2Z4+4TkFv5hJC9Yty1Zl2Wp126zR+OnUU7I3dK
iKK4DBweItgATMadS3fMPTBidVz+3u6b6UXzN9kh3YuMZTXTLFBntn+8PCqAege1h+3XRHMijE6d
gkfSCVvYMJ6ReaWzFGg0CvREdRf4fJ6wugpCmWgUHB9UEFMeeRGZU1eIf7Kke6pxOE6rSQHzPE7J
lqq6tlAPDvurIKGGgins5HzgmoqvFdD2RlZ6Qao4YBfUHrE+XM1fKKtdK++Q68Slc+g8LJQn10ls
yoW4CQIiy+8fMN7wUh+9FNzgLCmAHMrsEUAb254kDrmbuEjrO0PYi/YoX9bRwBxWuyx+L9QWe2S5
KMXxAtvUdaF8QbY0nHwHxLzJZTBGr07NB55SUOTBKfZAufsE+Xcl5+7KDHmaskwjjXnUjOQ7a8eK
gftYNShJDe4lDIyH7ARuKSWDT1G1DUoQ99Upm8Dqz/g5qpefYY3XE0nP3EFOrtpD00TuTQtCv+7c
CUTDrmbCrRl3Au5MPS41xKbu0PSucaOeeW1pkwAGWruVjBz2uSr2jwNwwope0W0dTsV6epGse1P2
DJ95zwUvaL5/VVHVr/ip0MqBQbF5dS0WczcA96v8LargJNPjzJHhMr9viAbHC4vQVgurXHEFQDKL
BiiD5K56lN73nxrTVXj3og3BQrXtXxAJOo2p863NBGo6trPM0ovy5d/ZOVjEe76rVNnWYnbNgQWM
1GOKR20VtpkYlCI4nwqk6fv2mM0+aJmvO3GmJV8ADiOoFqg48gTtlpU2R7WX1wPSAIOJO7Amcj7H
LsxRr97w41CnmnyBNoDdk+Q5bS7GDgTBB/qMQku6eXk60c0cCAmvf7NY0u2JYm9n4u7OXCpLeBNu
mA/Hthjx/8cGbURXXwTwleZYsjWorG4q8FRujeZRgXuR1G5OqpUclqtzRNGgSErWqNeT55FGsC+5
NBAo3554uEhtHQC3Bjb0KWExLIV9RG8A9DjaJCCzZ2uyrjKVDMldDz4/yyCbFNSzJ3fy0XqjW8fJ
SAopl/rpkeAP57GqUJnRscyvv+IIznx27WM9ZdSFlAMSqvS4Vhgwxh3Kr/8YK8tcHAutmsoplFDv
rTKy7hcUW5OwKL73+s79UzbX6FFzA+i6lQN4FzBdNYHQgcKDb3Oz0uEAy3lrPqSqmU5txye9kDOt
A5M/bF2UnPz2pAHJKdBpKvXIk48jyWVdg5+2Kf1Hs/cv+dIC7wnqfR7OQskn2S0huTtF36habSki
2+dE/DzOkmYUSMa2H9IHPIn//TXuKqv0GCAzaPApY0erIEYKsu2aSWomPWFfY+9BIdv0nFUW5Eiu
EqApwMLKYxkB1t1kHTnTYFuPd0Y8qnQ2eDv3PlWE39hG3WukSpYB8bJHqZ5Mk7WzGi5+zEzjDX6B
p0h5uwtQ+sCV8Z4pk5xC/1LsWqWXVq0FI5NAwIHVsZJO2DQbxVlqn4/ZGHM7tsEVRUfbPjR8c1pC
z5hpKnyu1c5CzvqdxtoSrngEsC7X8itEJxZhTgk7z4SXNs3796eN6eIkV4pZj+4EMxeeN/EX6rrz
+852rNqLaoa66OPfR75trn3gHnmb+5lY9ApoKGBCpf90q24oLXr1ib+5lvkMidcKUGC4hP6JVYH7
3WPC5Jaof24pjpQDseyzGJALfwbhqfmCbB3YvdVX9COCgxYd7UJRvCMFGPVmJFqjyMYavyHinWWY
k8LsnoUyDUzdIMADHPufugl+w5Nq1S9BfEBo1+h/5qqxDqP0h0GGrToh1I5YITeq48M7v6/PuLT2
8bEHdfYZ7Fhw8iaIGac+pzWmhAE2qmCUeHQxEooBcAEj+1emRVcFMSEj5UhB9ExAujF6gtnMXx1/
Z/U35YxdsDG9qcH4o4qBTRQf4r/kpX9AIK44Ue6HKfGj+hux2buKwnFNSfq3TXqnmCTBrqiBtCiW
g2L4NJp6bAPxdwqZq7biFo9iigi8zTUtYawNo03O3NEjVAGKd+NVEUpqx62GJ1HrkIfSF1CXvH7+
p3rSPA+yUc3zjOkgjCGhNxv6J9XNxnxNbqge0jksjV7MW8IQajAqApBjxLdwzsDatlsPJAUcwzsh
9h/ugaGWg4QuUn81lelnk1LbyyQga60ONQ7yjkVIGsQt5vOa5oDGzyUYwKCq/xEB789nL+EFCzvz
pWWsKuL1G1xlWzlJ89WZEVG59Xy1a+MYZXuH7FUYXUBF69TvAfxjK/sgyu5fCm8Yp12qc2R4Th3I
ZcB0UcrFsxUvXPGatnmh8iP1Vhs19IKz7ShB6isCjDMJoFTZW1dJrh9XjtlZGweG7jnwX/1fhBsZ
2HI5lm5q10LLxIDcCbKEr59fM/2re+oc3A5EMy70HDbupk73QsgdSIiGNmMNRKB2oqFsvS4DjcCY
7/ElzVhnQPbjUpqvAXaoeC7g69TjelgOZjT2OrtFPLtfGvnTF1WrAEktPpUihAOliY26jryWWsv5
FvJo3+kSlKNo9K4IWLeColR+RB94HYB7H6Ppr/8pBkMvHPunZw3D5xSOQkkU2KWzBhjnJmIOTbNz
yWBdignVOVd4T6bT0QrcW7YlVhg4JVAS3pXQrfjQ4xXPgk4U4LaiUiE++qxpoUzzVbQz/NSjBrmg
UtJHn0Yuo9KUTNTHZYXW0da3Kv7YMCGVEdsAa+PLA3uVHmLfXTFUScUhHbbuSMdSck0uOsEcVmi3
WOm2lMtJ8nP6KDFXGEV+ygVeqhQ0BOViP1Y+ffH9h+wOpo5qehWLvDzVgiDm7Vu2LHhTAhuFlxK8
AKo8jCZng/JtAQph3IL6RnzdPlwstv6vvB2bxiHtFYhJk2xcg0LRm/Zbz9OrLrd9ClaMAzFdEWf6
3/qygiFPc3Cz3ByM+430r0+JPnhe2dgCphxaHy6Z8n+KavfT3aABzcQgNlckOuzFsVJ1bkHNrtO7
CNtHKg7WMNFUHAfhjWReWLFk4j9oXYT4674oCVCPKSrlGsSR4RokpLTru557BejPSHOOwixVp/ni
i2mpveCvy+i/ZOR4wGzWFSJ3q8wI2NbduZdeYiA/hoW29ME/MOOCXgTTa+UnmUns7bM3jI5Qyfhr
7WrX1t+kRrQqoUTeEKGLV6pg9HO1txBcO8shPU5hMchMVn6k2pYg1wnIID8vcEKW1j21xtMBk/oD
xCkbFu0UjEBBCVlK5lWkEqKqMUDfY/s2f744X0Yy1TGgPRd1qiyt9PFmVabrx0OmdZvEeg4asH9R
HTQngMS5w6tArZwXo5p2D8Iu7OC8AHAWF0Uo2RZsZDLzLxKWX7ncDS0Yag14H0hzoywbqeAybWj1
AgAVEUFNMXDjEhfAd5hcjErQl4nzR0HLTT6KouhRj9mStIJKQtCwppYIO7uTw2MDcrJrm43UBVUV
4JEPO2gFX1s4GXXSCWQHnMJLblqPZAqJk8rIBmP3PxG35WR7l0wVHlcq2H9jWi1jvHaLlUDkTxCG
D6+XyZchk2u5FOQnMnru+G7x2D9EnYBWLipU23JOsehWnZW7ZI4HJekDymjLyCIRu0HrBhIcqxyT
9867N7FswfSuuvBcilsWkSa8N/Yy60Itm+aGVXonaVuW3Fpnu44+gn3SuH/5ucAR4KESf+SdMmM1
I1Q5tsUd6ShW/bdWud+MPqPEONGO2lLwl3DdpaedrKqnZqyYf4nZl5gUErMvGkX3ckFzb6RShYs5
LEogsddYjOW0ZE4guRTCTP09BzZrgsHP/g+7OKly+d2O5NMY0NVyowBH+yBDLGtYh7KNfWtcuLn5
6HNMD4mVMQ53BeWSQD3bMWLZiEjHAlnkjgkcwS/JYyqGPl2jf6mYP1mN0J2aFxm9qLEmSW8ALDTg
S0o+IEaUzCYX0oC6GhHBPaXYW1OfrqKnmX0A2pZNgbIjrgWq03D8ypGymYs9T1n9qnBIYix80S28
fK4ao5P6p2mP8VetTIL2sZRg9RJuUo1Hyz/XoHxJ15n0KG1ula5Au5q1dgoVJtmAvHrcxB5duF+V
BQMmTDNUuaEig0OkJuR2BeP1zbIPxl9YEKHFg8mME1AP0AgNN6Ug5jucCsifLEX4qruwB9Q25992
HzyR7Syo1yYZMNtgEhpttzXBY17FWz7mJhEZQhejtXzkXW4glQzEqz9/IRzbm7YQ2+sjPJmhmbGv
Coje4msYqNFVK4NQzoqEC0SZnsyewCgIwu0KS6T/2k/zinGvm7jllSh5cl6hJtDfbMVHVqvbungf
RRE9bQ/M5stbANMZsoVrGwROkAYD4TPATvAhV56Vo3kUJQy9vWaM5pabkdlqzsBNPxeFb+GFL5sX
TC6XekK0bN03FYxIbDGTI/8JOUWPkUn+s7sFmfGKKeBg8BhrTV9rtl+HMUkFyiv888rV1G16i1hx
C6bdpQdsoROTxZAGFCRXX1qCZjHMiNhbpdLI8wplvJFimTf7SWt8NdOd5QKRbMZHt/ZfOXk3HJaO
ysy1gSLYKToKV0OrpfdQmEZ5X2jBeV/oUFKw5o9S4UnFwED2+HaZqiMHIR5eqeBDW53ypKuLdXDm
NX6ObImfJi8+ZOp4FBUKnex06P6yG5JVdy2WsTVGBNX7M9TTwU7IyOM4vskC2G1RtyxowJ0gMmzU
tk0bNNybjvvdeQbv+ZTOx59mDAUOw64SZmVj7wDHfeKLm6SSE1RdenoX5iIuzt5nF4Gl7GaYFLey
XUCwM5U2k0vlOqd5Jdf07Nx0ArLxA/n0mBproV/x7RY99aCKf4uPAWjJgg2vjqvH9wh3oY79CQy6
OZL/DAURuHbeJ6bbKjYLjd4dz/QBizZ7S4JECdU/rm4KLa3xOPCVigcCL42VVaWULIu//P3Aafjp
CUzNG4/aIDOE04AFzqWWCJfvYHuUgk9AJUxt29HVNu2c+0fPeGaWM/QB+BMmcp5OtDYE6ywOi/mS
ZkBpdEoaIwBM0fzSBzDTZ5DU0Qp7PTyUH6KcGiNt5qLWAp9dd1gxr6cwriyrvX/PQgROHEaVLZOa
VYn+brN0aG4uTpov2hHqGkS+olQuXzVdHASSu5J67qjsNdRwAfLpV/ZMt3wuKYR+2AvoTIGqyLqz
4yO482PnxYwB3wq1LTuS3PJPabG1VoVzKYnqoSeIica0ttgHdx2q6QFTNtNd+zmKdcWTq5JepJlj
yNJpZ+pZC9ic8oZD1JCs74yjQ1EtheIiztpLCtaaiEz6SDqCy8WpAaEbmobK8I2jARkZVYR3NlZI
3hRGfTUfok9vmYi5tyW1+UKPlU/68SvneR7t3IPy3yimqX34KFYzeQjJIvH1PVqRgyfwBLQNRcBm
tvSezpozgkiH3m0lUDy1WcjnZ5t80RXuASdffcW7tyyN+I4n1Q9MidbJspRh7qM9kYgjTN8a6eVE
OEsXSaCYmB5KmGtK4BSw3leL2zZjYX3Jnh7hBVzL+BRg4KEfvskFbb/iozGzdyYU/rfWH2HxNgby
uLqHMANjReK2qu2C0ee5N4UZmEDdb9Nnsgnk96QDmAXx/xOZbX+ouju2zKLonRiUPJIJjiXt3QOU
CdfYdBYn0JkX/fRuMepAz5UpTFbibYt064e0w/FsEWXxa1/Ln1QOCOgbcNRJoultd8Wwohx7Z+Z8
Lc72nw2FZxe8RB8Rj2fGMNr5NcQxAlHm04E+wcKMJFFqKPULiMat0gHVYB55ITKbLFSI9sbGQL/j
QzYGG3bQL3jr/yz+KaeQpmVk5SeJwkPNDwK/g5UTtgnw1IAb1BjoKQZC1wg87ln8y2DsbbdH/Pmc
nWWHdrBiVeSBY8/FZ9h79N9xejPf/O4sey4dYCDIrfQp0dh6mUN87CqnvA7d6sDjlYeMLfU0abKS
pb7somK2FiEE1Ehnnybn0dGyE35beKRu4dgZCvXIgN8r6ZZMJsCJ/dSpjMh6HYjlEa1mgLVDkGNe
GPoxG9lOjV5CnM+WuucbPCeWTK5fXRFNuOjERwwNw3+JFqBUnUFxjIhxwbQyLzp2Bp05kD+XARe/
dM6DljCPnzgq/fcrsANLD97FnERsw8UdPoOz2PjHae2MQwmDzgzuTRHcSYFiV+xLuboSbuCjG7Aw
gZf41Wj1JtfC1SveuvOZuFtSbuxSeqJr/h1vkR/Ey3aPWVC1WmxhLRL59PJPaBrVFCRj9eC00kDK
jdN4QwwLMMKp8zj7bBiBJ9iYFHVh712VVGVqB6cvC2YSFdFXUtD2j7dOQOt71V4zoFrJG1WyOK5D
bKq2Qp2L+XkqmrKz7q9jlNkFUzbP2Qr6JKM7g2T+kaOd/kRhJdNR6y4lVDZSqiy3pbnfW2A0gB6M
+abXKIozWLJsKVZiGBtnSoHIdBZpFmz4ui83sVSsSEmTE7qGmuuAolVMQnLt4x2KMXYPD9/iDlAo
tP8ugHardEfJdAlVpaSV9SyY4fciGwjKILxdkhhHCLYquARdD1WrOOHRCHve7j6YaqQA+qVL8TfM
9c9tqBl6f/YNPlCyMWOhJp0laRefKKljjFbFAQka9KwfalcAd7MGGyQKaYJqKtcuRmnhuqHpSqcI
olFNPlNzmblZu4wF7Krv9S4NMQ2zN5Uc2uX0zcFBRmCuquOW3uv+Gg7S361KMCy26+yczT5uJLhx
+o0EDwnsGZ0h1Rp3TYZjiG1hrmCG4tjl29W9GJj0vCoevkxjV2NmWoHT1+CMr9MGLNrT72zMTRyf
BN4Rf5c+hiRb3mggpmW8RtCPkwQ9YFThwPkx+kTyQnCZHV/i5wSRusAlbV/mVenVRCEvfvK6yCCU
o5cSfTfT0djSCTNshFvG2rm5VC0CisJ9Tiva+JNIFZYToNAE01iqr5h7cldwtZA51GcLLL/AxiMN
spWSLCUM/56cQVGo9KGccCc4jc4eBmtbUiWrSwuJDCQTEdjWd8gn1y+UDxdDnvBBjaduqm7UdBzr
q+tKRqInJ/DxSK47OAC2I0/BHzK1rd2dzcJ+IWAiluJPTTC8s9mDApYpRsUDSzeCjdei5X+fDGly
xAOBayCQnUjGMhoCOT7lXD1VeX+9uRcmJUgz25DrcQENK1Jhj7SLeisfxibQNG2rjcZaBOzpNiie
Pzu+CCOUdijB99MHqCXPTmqjErsQKJTlawzt+UFzearYYq0SRcplin/hS4hBW/p258vg/m4McW5V
sTOUgLKBL4hHIKKMtbxlPGNOYnZtsij7/ktUeqCSIWENaELFT+4jNVXDw/0aBN/3hsRL6pLnP3KA
nJjscu0ZqFcRKReBvUNTZhaYBlKSv4oWVs17p73UiaVFFG0Pi7jjCS5+DDmEACzT11adhUplkBcT
SqNSlT7lXsKVGCQoDeErXaaZC8qTUw1kfYfwMxpzR2ER8j/p16qiaAJaNgYidDVoHc95to47SPbd
qvhCv5Kz1PsyvLE1WVouZxcpv4FyYbXNrxKQgJE2+h6HUp1gc7XDCvBkCfPB5Hsv3CnNR48cb1Fv
0bODPSPg628pnKKA3xfVTdzRl730Ai0hUlDs7xCF1I+n/0xO0THRCPFnNaWNz7/aHURYfmrSwkST
Pi+vP+EgxMxa0IMfmJq5uqpqLEEwkZwZvH2z0/R2nXuHSZFnBvpnUHoHWkEod5kJfoOnUT0bTtH3
/OD/LfuZpzqBxcvHfBAags7TZH4xqoYiS7uJ265B24RVcmZ6c+Qzy0vavQs9PyZI5G3MqCnUhfM6
zxWmGVDq1glRD2LXTNpxVDoiRmICINGdk0BGZoxBh2NovnKp6PL2jje73/HEijVx0/w5Yjpbmsxy
fK3uZqcVxQM1P6Ama/VKmrKFlJPF8vVWuqr1TLJGV7JYlHY6lUjOB2ltLL612hUQ1Aax81UNx3Mu
sAQF54Y68JY7V550/pgz216UssP+FgxQvoqScHk6MNQXXIstXaFurdI0EGXUsyNvS3DXCyMit6kX
j65HXGrQA5A0ZLyb8ZkCNqZYMZw+tmK1X5q0BAz0tQy7UheAexNywgCK0mBTBwcDNDEc7bSxHj++
63EBSU5+N+0wYxxAJzWaKaDnUpmOjsMfVWnfepGVGFv9Nw3VejoNmAuMd6NHjkEP8YdYxRLSTbWF
FgU0+tx5ekVyVLFiQCmAhc/pK+myrMOIz7wfg710d55xZ/P0brPZN6xhmcn9TbIj2fLj5Yy+6erH
R7/NmH8R5WrPitFDAXki1g9QbIcpDOJp9d4JbPPsst1KO6/eTC6Uj/bYdvX9k0tEMr6CnsIY+5vC
rMRVj/Hrcl6925mr2/rlzes0pi/KgW72tl4rwW63GWCBWrPDnW+7y0hXjEKd3/9qI37fXkT5D0wg
Fr1ajNmtKO4yBXRNlaPmsuLx5iY97qrvHMdLV3DRkU3PsDTsjHa/CWcp3vKzhzw+tTO1XlmtutNB
Rk89ebnByiOHaNw/ZEH+p7bsJm30g0gmYZ8rBAZGNOW/UC6d4adQN8RhM3gZw/xgoPr1fHzq5fIr
kxSKCZma5M1Np57452cyeePlJBYADnzVz8S7vnIdfqTI6fSsIeYzTkwKnAD6FIEUpZTJU1G5s+sM
pIbFp1QExQazgJBRw2nJysXrnBWBXtSW6JrPG7tQPlVX74J4ru2FXv2ejagSj2qT6mvxHmTHKROC
gEogT16BYNgNFJxAI/ZmzRielrbMm7diRhg+O92jB+JpYkBhtSAA9bD+emtQJPGiIi+9m3t13CqT
ig3XDnIMAxipL2B22gGy3YTPyffGZ6Kei0PfZDUV62b4ee9mSVY3OUQ/NHUsB3To/8+NpERnH6Wj
7WJJkh2feE2Dm7yBrsuPR2ogs4C2jfyX4bL5f/6sqi0Ebir5Pa5T4vy+swP9MX1kS+pOQCrMNiQL
QugW0TYznZyrgqbSuUrAihT94ykrr6eE9Ank0QgAJ6m628Z/gFNDEbt4u19YeR9/gdsAFXo3Wuo2
pbUNBFj0IhHWFcgsbIX2woXVx0ggyl3hrZIzkC3wGQ5XKpnBuyXkEeELUmWHWy+CKO23OisYOI52
rs+Ii3LITlFuq34aieUkcgoXrWrKJlkS1SJVoHF5X8HmRvt098re9go664cFRDhgPIK7OExj8ixp
AgcpHjW/kogZ7/UhY93GfzlsX1YabDWE/fbwHM7bz9hH1MGWhoNCmS6pByW0zVBSa/2NZ/YqXD8D
vGQoUo1QhW3pVI6Lwa7V3eghsiectc+A8UjYxU9Ni3vinqHZDUrZkWAb9Cje6OL4ztcxn9GwREEe
okw8PWuvopw/Uc5vcda9wxV+YAZap+WV7b7Q79nkx7pNke/G4RXWVYNT+6L9vVokufaa2cBqIKvi
N8RoFiRxZvJtJY3OpaDbfAAvcHcxKyRUpPdCaqKJ7EmbWL7QrJZo+cE0YKNK9KdKPcBGXkgXgbAx
hy9Q/qrKQ445wsa0BZJloxJWDCACzdQulZUeHYO6FOEcEYsA0n4ap8Bqv2UEKx5azEPUZwKO+KQK
djhn+9iew1E6/nxoZjWP0U/YTsiYcdnZbiwEGd8DYRG2SBZNaNGO7a+iRG3tQ873SlgOfeJSscJ/
e/ubrgEPThmYx7+Q+w30dFbLQntZzE8qB5Kln8fkFSK3ZcLkp91Hy19AU9rmP3WJC8Ch+A1VXbZ4
lJ2Y6XD8QTzV47cgCDp/VTLU+BVoRsFspwiChAplNFLYzt2waF0dDW5+Ei1xvynZEyaf2uIaQuig
FrX+wNqw+e99xjVJ2lue5Xu6n1/t2G4otxfAEf+qgiLtoFKhNSx2uMkNrNO3xB5Q/qVAJTCaKbeo
nIXbylPl2jaqaILtvbJ4hFt09cjzE8xvhHhUrggJNhc62UOAcQrt/193ooN5Z7NztC8hbqb/7BNH
/TaQStrpqbWYX7vt0ophiSC3+4uIcpKu9SH/ODQ3DuRtAEZBfZ4NAys+IRnkxX0tTv3sj5U5Ozf0
gBpEHM1KDX0RexLz5/yRtFSlCiyxG6yio5q/+/Rh+Hwh/APBUqfTqm5c+LvdsNIRMIHntlcIlYMW
udt0i2Xx0mzHGH2EXeQrR4GkoMKz97LhY70dMvhUjhQxI/pBAdjdeNz+WjmkrccueN6J8hx6W4/y
tbVCrEvyDOg7ZfMLRYieND9o8cOldCfrhjlWImhTk2MJScgPZuIJxfHpmpl6W8vU4FemuzNWcNC3
mO3m9OcKlvfKPj8S8FLuuVBhV82xDc6vYwE4c08JecsxTcE1OzccYSp7t7OdXQOknwoRPyndm5tI
U1Lgeu9sL6Z53GWMEw+EePaUZyxCVQbVfWpto5DnxWe8bKhTTzsHbzKkiz0+vev80IDGR+LdCEIZ
7DWDZwJtfpIc0j0APtYY58CVWVb/6cWwxTA+BQWPQFjM2XuUdDAFGXd4QrGXzPVOXq+fnIRgIOte
fIoobzm2RbRz2ptdSh5QD66l/aFUrlEgMRiiOaVkkRzNjlrOsOwyFI0ZHzvwMyprGDR1tOhutDLh
NXzkMxYSTrsJvzrbApBRMgE/+hEIYYkk7EO0k/YF59sJxFb5N6Lo0phyQLwFOb06FFavtEJZ2/yL
7PdyQEgn/jtYZfXb+gmfzK155EHHHNi0bm33pmPqhU11SzZpc/W5FXWiNOl1vRmGHDnBx31PP2D/
QAVI8N1t3P2boyEmfPqCpnMGZgDMHShQne+f3Ptr7OYs1WMMIZKaWp6dN+OuQLCoU8Whdqhg8M0h
qXVeXkdPuPf3oSnyzF0fVI1izdwO3QL0oRMrrxOqvUYmS9eHTTXHApSXWhuJ4hsNvj44PGz7F6YU
am864CF3sq6nOFb61S+Xo5RpidM0/glnZJg7KbT/rKy727z7OdNShM0qURGwXE3zF/w7pc1Uhdb6
iQpbleZFlXkMObalbJGe2uydKc4KL4qLQeKkhnbLFj3fZ18EMPfR6qlDP40GOIwrBw/KCi/dpBdc
/WOMC2bXs8ybbn/Zr8DCWgzsJxoB13N19Ep3SxYrGiTeUCVqn4UdTRo6QtcRahweR8ReUGviKUNT
QwaCtVluUP9NL7DcgZKmWzhA6a6Vz2q7jNydSogBj9F7Ii/J/PbBWxokcaPtBIte3BF3FxeOBLuL
UwXvJmiWAbKFYgVJWMon/iPSt+RqCRlF+icnd4xWyhZN3czKCmiiSf0ztRKpBWHqMUXz4aDxRIaW
6V54ngd0h+IYcpzBHazTDf3egPexAMxvS6Iwyksc8Lf/FZ3IxA1ZbNAZK6QDIYqp7adm8qDJi98h
rMT8IJo9ALwLV8j1E/E3AWnxFmOITC5tJzFDwiO3HlWLGHlXrZT7fi7TT1gmVx65ja4fxwWGM90b
3uBscKmh2mLa/74FsvT5FEEQJjyM17Nlch4ssndUhljg3eVuAojDLYMRq7TEtXWsSpxHx+XontNd
ZQl3wQNFqaVF7q/Sf3VVkH3Ww99bCQaRsSASCazfvN3AOdUm20KcHhDFZ4/8TlHEpygKeIcPQxd7
3JjLlSVpcXrFof9eH039SvRaLthQ2rUtvKLyydUAyJQ9oA35GOg30+Nvkl2ljCeAGgO55DQz8XkP
pQZQtONUtXC1vWZvhqmVJJFtVlKe329KpVIcfR9NyW96ATcwvzqv6WwEV0daDggeDNjOknVm6Cv4
a8K5KFOACtZ8EjKZvCfv3JFPZUeKzG6tL1gtyHfiK6sQhuhAa7zOpa24ugh8e2R6itGnNoEMZh9x
ximbNb4hn6Z37NoByX3oFB7aTsXFqJyDg17yEJrUKxuyRUl3+dynVVnxLt5ngDvDAQv4B+49A1D6
/X/VQkC7OHdjYZVtOSjtlrOehqBubrgDQ1Jm8Kfy+Xua3WSnDhvPIRraX0jXTq5rDV8qpYO9zUIt
t4QyAGkICkYLviOSo0r83IHjcOcCj1yV2XJbjui7TMabAenf07U4c61Mr+vbKWKqYyq/72WfeQiA
sX8RpNKKX5/UjiGhYdY7UrtG1P5G38+wg+tSH+wABWFDZJYlBH+OK4yh5l4xnAjCzKfzLcEZbVUn
V97TsFWL95R4QXBplJW9loYxV5CkZwLXwATOSQf9BPIs8/8od47+xGc0yc4b6DbjbCt64vDnPjt3
jVli0r1EldTSK2pp6892si+cRgtqQiB9fPCoW3LzuaL1/n05OtpUFW+0MAnsRR4R5c2IP1FbFqla
pAVu6aLEK3+DMy2fDOk9xFKI98blVIhQsKm/bRavPx13DF3y//YVlETofKLxiSC4Q7CORITMX5+8
LLP4MvK2ml92GCQfVpTP3lp9bytenkmP4tymqJPtMA2mA0CKW0O+2aybVM11q6Db6qaRTODj0pAf
mAJ30Tw/PZOtHobt9j7b6WmMeie7r3wepxM1yM8kctr0lMQBUSp+NEYvH8xSilF3aN67e4HioJ4v
aAiDDQB/bIS+53rIwewBIfWKKdUZj8Z42rOsjUKKyJguWyvNmrj5X1E5xGQYSX3V+5VsOQi8d9cK
LbYVoWi6dSy6mTMco2CYK6Rp7xgrd5kxas0mwqdaruw4Src5sEN+9aP9kA/JPb9kDbLgLEZpq1N8
TtIeSj6G95Byr+Ea3a/JCKXCgpUJ2Rdf6n2mnRGoucbov7v/F0NspNIjtATC8VfjG6VO8FKlDlj+
5QNbfH4O4yGdpQbwgBNV7m5UJNSvDpn+gQTrTwnxOlNcEwWJMIcfWPMdNW2Yggxb7GBpRpGpX0Qu
dNpwONnHiNqq8QRCDLQzjQ91rkLRNCwEiJxvCFma/JwLp/hzJRQtSiyjSORX1gecmLIhPQiQCw0e
moS8+GT3ZiCyG7UpI5u0TuPQjup7z0zTfwM0XOpq4yn2L3ByRFfqFthZK8EmxwyQSF8C3T4A7Blh
XvDnl9+YES00ooSxX0XQzNyp313JLAT6hRYAbbZ1YB3ZI6KR05kOgxvpuloIxfTorDvFohUXZqCF
k8RyML3jn7T2cOYgNysKUYKWpD9H2k3sA2hMpJBLmUQmb3HLSDgJSgl40aY+jsxx9sGihewj3TUD
VZtfv/7TXlQkXuALN6zREgfz1fwjr1JMV2gpMNBVtRxRP1U6Y56hsozxuWLpKQRW5ichk1fM1qal
kF5KMtk7B+v4MQXjNkal0bXP8slO1T3IDD6OKDd6oF+aT14alfyd+oavSQu4z4y462x8QXTPzFJZ
chLqTFFpDZ0cT8NZ2LGuq51qd2mRGuDlHGxweI/N7HZ9kD358Hn/1quvJOSg2GRlHc/QmyZ1YYBN
ElViaEQrEUeJK2oJyxhO5Nv0XMJ5BdooksUJEgPsPOx2zM51mlrzA+G8iFeNlABMFRv1mlPXkNnX
Y3VM8OIKxbYivurp6zyhJpy6ke0iO3eItdLFKLObLIR18rvSo57HXcqhjbeGAuSUdy75iO6ULw+E
Xzpg/SnK5GqwZnr6PF2r9cDT3UX7mprP6Bw2NT6RWeMVilVNhs30nZ4CIScIVsSNMUPRwlPPNxtq
NhhxXVWThpWPHtDBw7eoPs5WHlB8A6qMAUtVkYw/9NKfCgm3mVw7oB/ph6ZCRW5ApPEcIuvBT2af
G22xASbkNlltNuryn1Z+fjNwnKnuzapS1I/Y8Pyr/u/wJtZeEGxuXVv8JU+pxqMTF7uTWBF73Dx/
FVF5CmyPONS42a9kjrZghmbp1vzaZKFEjXSOZSE6nH0l4joPbBdO7aC1WXemx5sOXcc83PtoJ+eR
hEvtoTksf84/2xqSXLy71VeNNzgRWD92IFaVn9G6HNjMhhEJkgG2sFx7M1ZJyB5+ZMDbvLqgFMzv
jILE0LHk24vIoL4AVGUwjbDI5zesptzOcb1IYUaoK2N9pH5cLrB0uGeJ3Wb+V0UCMH3Vsy6Y3Xo8
rz8PtbFFyqh6q/7n48asjImWEuWtBhecNubIB3UoR8toaDDe54YfhFBwPh5hhNWNQm++rdP/LFxs
YqMSecZQBQwJlrfsPu2qH5jFwCeeptf5l6Z3ViH0XAmVz8aIXfx2UtbSYPYfNDYFWhV/djDPJU2z
vaYf8OHVDEDmoLrZSrvKWtSTweFilTeRY0exUuI/eKwUeLOIV5xWocn0cuJ7UTMip4nqeu5Vx3rL
tVbZnl9gzn6bIoL0LMPijDDMkxRvExiflef3J+SDcY0WFx9UIZmprsxNFzlRpxNK1b+MrguCis25
igoQT0jkyvXxzrdSWVXhqXkOsbrOnTvvFo2fCYtguFawjVHpKXbR02uBzqZNHOB8PpPeJO/McbwB
NR02N0J89v7o2k1zTBxQ8uKtHQnyglliPlfNjR+iGbjBtUtrdeUAML2lUWVQMH0iexA4b23Pknq4
Y4zyujjqiPCmkcsKtlfiU7ctBC2Aul2NNv5yfqTKcYKhlEd4sgxgeYfxZhJHEsKgAUye6Olb0byo
02Sze3WQIEqCy5ughd4VbcogF1OOtc50uEPL7tEpBawdAi9NOGnbHXawr5vYaOGequtHsP/QKac5
shoVmoGwZ7wAI5g+6+AFy7P+Au5+8cvTJ/qj3U+6EVKVMNjWJOEQGXAwhPsJuaY7ooL639jLwhDX
jNXLX6+QwfY3duwY2gh6OGzuDF+DP5D+LRp7NutojSbaF8aJICelOHxWumn3QAOJC0p7qRBGHzaE
waauUEMSCdzAQEB7a/NK8nX+EMO1IzPAaqJmBEdAvgK5ZoKHXo9KyABPh1pF/vCbM166PFmUJaI5
Mh+vgsJFr5eR18xYwPeIRYZ413nazvq0j+QQ5CB7etZZOrTDQcptgZ8aM5OFW976NoYoBqnHoc2L
onWltQEWFre0KSSdBfTBMJFXS5QR5foYWjkmLZx9iGH5mNxwwVWQZTvWQFnctntxD6ZeSIhhGZfR
2pcnYMzNgJejcCj9vrM6Q1mwtT3rKU4efb1y1r0g6fxtgRImEXSehJ0nUKcJd4e4LEwxsnND0VOw
r4egFGTWxL3V9Ua0fnsxfcQVmAEZo4wGdcUGIFlvVlikxNHpOZPfc7p0nqbBfTfalk3YWqrHiY2v
yewYZz9zOuc04Q4AEhvxUxJ+ccATrV3E8QTT4NKzTTNkuJVqv0VWGaHImCBNW+UchCFVEgqTquYH
Y9TDkKwSCG7CapWF06LRKhYYMhTrjYeBLJ3d7pnxlTtxMloG8tGWTqbo6DUA+LVkofCk7R/uRV6p
N88tNHxzdonT3I9b+rV68zDN4zeg/ARoqL909pgcxbaT/DufQ72PfszgWakIBmkZpkGo08W0Fjz+
XlMUKkr5t9b0WwzzlvtlQuDuqFx/dRcRLJAFxuGw87sgjryAFLtIwPCur8QUh1qWvAqlMaYIIiG8
mQEMuQx/xaeD2BWxp81ceu40RdfwUXhgQJhaCaXxvbc61VGBQ8V9m47JLRomVv5K/t1fe5c4Ymra
tLUj4KKPGHqGNA2ra6d2FE2kbmo6Yq9BadoXgba+velysq3Z3jniUi19K3jCRp++6HXVoE/F4Drm
RvIYe9Lk59I+ukwZZDk8dMaSxVPfoCiRtMcms9jCHNebFx5BZYcUfItL1Iuj49dEyZhOATJT6/1C
8HLYsWqfZgAJ/phSU8any/L3/sqQw7ujnns/XDiheEzln8l18K5EJd5VIzjORSHqAf8UNiMYOpjT
m31czcUk+Q+SI4yiKFWJ/iE/nRO2SRdU43TknR6UbkwrCzMOa1mV4WSBT3j/TKBiw5fXKOtQGiPd
6hS2GFNrWi2ln7PeiC+Ajfse1e+1e/JfPc6lng4rQNDMIwj+2/zR86roeiYDNqNNLdKJFDK18Qux
1B03QIBPv6txcdk/tRZgmfaUFRw9FY8X1QTHM3L+W4/0MBvH9SpOjHpa44S3E+xsPXqJpfaNVerp
FxZM4W8BXBQWwdFKRldmKHElKYZ/NmwcVIAH5Vh60gpdsopP8EdAV1JU6lBXmF0GaLBRrAt8rqW9
egDKx2ZVFqkCDeYVOI1AM4RAkakpCSUY7NftY6o/87SHwMObdrUEA3oRqdtKj4+zY3JH01hr6mvw
k1ugH1uUuNjfrDEFNYu+7I4eDFC/p1H4P+WMOlJzRmdL3Q2DMDzXfVuxo/B+gItPqjjh7RichJn9
seK/5iTQBHAqpe5gSyt5G09/W3hefaIGyDcVLRx8OFkrAGoVxFmhtdSqtGUCN0iX8SJsww1Q5j/A
4P/ObaKyK4B1S/aBVvP2dYkrrLyoPzG1hhqiq78QW8CSEl5AjM+5qdSLTJfqQAD7bYAOr6QIP3UJ
PtuVsDgdzj4q50S+1IWmAn4UtDS7HLJh7Phx3EYk2s/rFo+aowMaFWOKuRsfa9LuyjrurjdYhshu
Tpe91OnmAOzs2gzVryp1iAxiElzpHifQbHFQjiGmpgsgGq7UtOjIXGmn9Kadgg8o62Y4G83TleBR
EfeXgpP8F0bGKNGR5883f/ooRog2jvaing5rpyJo2HGyjHK1aFQqNY0Iq/lNnms8diUrRM+bJDi2
YcRUJyJ7pJZfQ+dHhHMMQUFDUEoZis+ABDoujE3hKwixXJQcwHCirsrPqfCYYVwCBiZI0uo5jnQn
d9RD+UbBpaQIVwUKSLrO6Syyi9Nvq8cxT+PdfWSphXRNZLMYUkU8dShC+oQThrAfaQCNJwTYJYmc
v2Obo85Hz0qc+uR5lrKghX1dledidtNtGhaiO8mBWJkB/jdOeoN48F5ZiSoYFOZCKrAKxpj+J8lA
5Qe/PmLioOpWWZwE53IMxsO6gmln6v5ppWe++aOKywlCaW9+QvSPlIpxg1Vgdckgh7AljYJWFJIS
LEI6GBnCxX/o75qPCO41p2dMpyIuhbrEu0rKFSnsV7iZT8tliMFW4KkhNvQj1UDsZ7bidbErMJTN
BijRdsNpUlfqrHnxBWY+G2OGVtcm89ZVtkmwNBy/yy88O4X9kXa1O+y1CAZ1KK+sY7FldUP45cQ4
6Fs3YGnCRJDI0uqR7X2I85Mxuo4+XEocX3dzHlt+oiDCtYxKaMJBaRj4HJOvtog64j1OwIY1Dx+W
rGe0LmjLDZs74c7RpdTFkJMbYelWkUtvYliiiIRTDoA8/fQHGZ8lRLdAiwYb+QtpOnsCEUatlvBc
wZDE06iw+fdTYFQq8AR8lRv0WtjfuDPU2f8XoZeQMuw04DHgeCUrzzWB3Ul86m1hQ116MOy0bqZY
xYIJHLajcSfRsg6mgG94BWItGGWmXeOnGI/A3lo0mbM7QTTo89thxBktkhaVOTxYajAYUZ52jasc
/aIzWJV230BWRlVFAyDeRuA+SOedDz3+3oGWWPZ7gsrgRT6Yi1FD0Hef1jEQANh2WxTVe+7a1R2e
4Ywh9+Qsu8CQEmK0C/SadroMW+NcNu61N8Sl6LjLdUmjTUFtot41W4asXPZ9Gn+LH+M03DHYBvEz
XCauRKnYglEx4UWtfBq/7QSNS6e2UXcHHzbQgLM3sWvmZjTbfqpIx9vqrtZ+sktA5OiBbHPGy5wE
rg5boLs7OFtNkbyd1Pk8sDafyTdaXzIydFVJYvESpJvVEc8Xyg522HC3s7IgZZgOPPVfre/1Ew+T
ycl7SnrUr5ucuzwCuHGLAolCZBbCPh5x3XecIB/kias1yCmhyZ59lJIvcf8xsbL57xWB3VkQCoUw
5A9hAeUDgk5na809I8MiGVWFIHB7twsqzCPXVkZGvbJgu5N/EqVauSmHBD2HyVb49c2MF9qM8ZXq
hsvZSCulgYE1nTEsjvTa4KaCubqtxJqeef9WeIRTUP7Ewe3me4HBhkdoVTpvlzzHI/p3jSQcXbir
xEH/9ypelX4A0q8rmfmLCRw0q6B80P7wwNuDUys40Ndom9ctM8szI4bHc+PyGgqtFERcpAeHRszO
IDyaglyJYfcHgAMhGbbjq4ELwOEMyUP7MiuMH76bgbzzzYdNLyPhHaYg5xHLByt3eGubMXUCOc/H
nP3TrMZFhZDEFw58OB3A5jGnBuqvGM2sIsYSaK7esro9aco7R5WnDKQGPTTGgSGHegXxUSSi0K1M
qY7LKLawdpOt//G7+tB7ihQqaUAY0GwHHVEAn64hpPvgF5sfzfl4CuvRCZU9VoAgsik3Dm/YjP5/
/Kn5+e4S+DXXNIqWdzg49EOlFnh64wkxJTrkM+CcT7D1GOCwncCcMRimRvJRNivnXltuMTEv+W61
N9zF8ES1PY7YVwmvoCAVwLGGfr4eEVZ3hAFOiK+3tto7oi22ehOvdfdPCYMuaLeQj8ChLv4veVnr
jFrxrkvkGdR6MpGZ6wuDvB96IWVle2Xbmj556QtFwcFN1Qgt0nY0GFSYGV3VcmICFnoabUUjQO9N
rNA+PZUKPXcU7YW0Nj+Rj1njITBUCUrozwjTJgbWljEi5vjfRNV0jDaaMuVyiE7Oqqr5qGLH6Dw+
DCkqJe8R4+uJeRgJB+KUwGApS/RcFN5qBKXYllx+OvH/n1ngaVL8C5CXSEmrUEvezy0hZwUn0ldW
eeDKMMl/RT01Ib+HXh3oNWbdkvG72l1mbPvY7hBKDNK4TPYOCgfLM2vkrnDgfOhMKmJ0StfgmaTI
YXw8sXCi4KIpFjYrLt3fSRUBKK9kkMb22vkXeIslQPD7u8DBxtolAmbJME6N6gdl3rTzJGG0DQvk
6RPQ4LeDzRL1Oca9fjg7r4Fe2NZu1a5Tl93PSKkuS2GFMvZ4VRL2j73EE6u8xya+PiUzglONlvv+
2BAidlYqUi/ZHHXPywbUQ+nFxBkVJdipwj6Pz/oCZoSN3D7AZZ8xFu5nGFzqkw0mZ3wWqlWXy+F/
/EJ8g+rXE1JdOrQSEU+bpmku0cHkcq/dXV64E09/1tlPkNADocTE9ZKUAGqflduo1Ulj/65dNUkn
0ZGuNBtWhjJ9ZA6Bksz/abedv/H2wInHHTxhAuCVtAWi1V/SR6aF9hQ557DdoxLMACNj+YCs3LtR
h+L1VqrsIthVf2C93mxusjk+nX4huy8whR7jeXqjL6KPNxB57lU8E/3wsyJQ5zgwxH6qPMo1f/RX
E4g6mEcN2eIxZvHlPsYkTk9RIRgFiB+ZjwXUdFQXlLYOJzxcNouNA/phkUep4MUkvKZS8+u+DsQc
+5zmZTOdfb+bb7TmhLa+tANKB8npEST9+OI9zpf9Cnhk9ehmHJO1QbEFjEe0r2AQFcsMdVjfc1Is
33Hy9CK/Li7JxzLIkPxgHFkJ/YMsQfj1W4Wdjc65S15Qa/7VslJ6vWL5cZYR3wO1+n6JkZ7nsC7s
5/u23WQM5cooJrywaZKghqsZTrA9m4lBk41pD8fmhQ9uPbBL1f78f4aWi24w5l8spWebdfxvEyi0
s9zhxd4DVTgKPeKPiSmlc4t6upahJNxR3rOCFA8ZIOvRHgNCm09DTUvsmXimQJb38lek/rqjLVPX
1BIJYmSnb2wn6dZsFNkS7JdwA86GGKUoL3RH7s50cYOOxLWlLnljTy+YYa5jqYX0wKs8Du+1/6Po
tuCHXq+Q6xWJlTkNffE1RtyVRwa+Kxv/3VcGTcvJXqKSlWkqrNnTb1casqZKNggcg3kMKR3Kv6nK
rFqhjuvKWBhTz+fS7XMMEXM4xSW1K6806vF9PUsUbDESYe5iTEbIxeG1dOfZd6Ij+He5rIM1/LhO
SqI8yq/DmGnxo08fFP/7EuDYTUxwcbPKVhGd209u/NSYniowjCO4zLA7JSL0YurEnYHymclJGbWd
yGWnL9ianAYAdgNXgiWMBl5ZvsE/Wyl7nYLDqgJ7sfltxSbWCO7l2WZv1e2hhGulfjyP9Gjx+VQw
tOjbYlzIQcxys6qf/bHUdetrg018ElAdBaxW0RQxBAJbGmXjVb3YhHGUp3T5yhhjtjOsCFgTlncW
PZ1OZmAg4LcSURVEwhf1BnFhqBJmHr/bSpwJzTItx6mVmM92bBBnt9g6lPUF49FBAQyAQUJN+Cp7
UlHUqCW2ojJu8EvfGFj2PymFuxyV+sSkQT02CUPDYz/cZj/C7J9zTb4I2Eg+57JQc6Li0n2GZU9s
W6a1ux/5T38vOKjlou4RqqCXiNNtzpSmZxyEJFVSTNDofPLMtC0vL5vkhLN29xFVceC1WgLE2jVu
2xaWWvvAmT+MNCqM253eHNIXgBlCI0FZ2Nxm5cXm8rpoe6YvCYBDEGhNmSsxM4DImwyPYfMc5i2b
YWugu/0Z4ho0UKuWwTGcxNbFfxG94RmtbfLlKp3pVEaN66HKwUfru4gJ/Lx0OC+rqZq5JohRsbeX
4uWrvNDIYrfoagjbwWtWAgsEpi4hSinUwYPX6GKXUWPuat/wnAv015Ze72Na772YFn/LI6P1NqmO
75np9dbwh9fm+9/jzta7vvquK17KfUQ3WDBRz/YNz5tTByjuXmIFHerfrlmSMi45hfuChC1l45mJ
fo7SEkTbwCQ5HtA8QTWREMBdccNjQRgX4s6V42l/br1KZW1u3aqdOW6pTmIa9InzzQdm2H0Qlpf3
+I1waC4DQtJq092RQirPfeI3xIlAAILl9KX4CPRfvcCGwgLSmY+Dzx2EFtEDllQ+iKQia50gYpJ/
iop/P3p2OqomRlhOhRqvnCX04hr1MvHwNwrUQLM6cCi0IHrDHQxS1VWUQxYrfc5s2K5NY/HpxFw/
aKE1P/I9FQJcjPO+M8rZbCPifmDmZmyXT8uRWxr/1zva8YqRZxg1v3WON+KsKWeDX/beuBfVl8/L
fHj75bD9yp2LYXPB8czM52tmfNlXrzmHGYKhqHGguIkTq+X7BXfnY5NTwQ3LYSKe1Zf/1YfZLgft
Do18bOlltGyXTCrVaaC/3pSavfE53mDpSV7Baho09gm5v3FPJqcintamYayoFBRivgUVVKfz9AsG
0r+f+JaSEdl+AVtLj9oopu8exjBEDB0YSdLrL+wWVPIOs6huUiyEU46Waznd/E6xR0IdONKes3kL
WtbzxrXipDzdFhTwWlXRiLJed+MxJ7tK3BStaGyFjgkGj7f2glDzgG7qbgoSP/nxKOk9c/+7CUSl
4YHiK08mDZ4sk/fdEMfEcQmFS/G0zMvTEMfGvNLXPI3XaN6gl7yfSUmr1CH1kiK65/y+csVM531s
kORkueq97x+qp8FxMTHkX7VUCKawM9PBc5vcMPDN6vRDZ5tBBTt8dCcaFmJBKHtgyVr2lrycxOdc
nk9WZAJzBZd61Bdz68ZtC+Ps9mZ7ctS4hDzqwloWp/Vg8aUQpJ+xoE7vd8uraf7qgL215M2+10VD
B2tR372XgsRYwNwgAIC1FIC0rmgECWuSr588saX3yj+XSgrAE56v7SZUxDPr8wEycQS35uC6YKNz
x1QYjB6rxmMnGCXGkPTi9cMpivaxNwxaDR5Z6A8Uj49QbXTmAG9TyM52TryhNGHBXwCnebM8HbG4
KlYdc3IpQbCap/Np4QYSd7Y0TAIhCQgW7tGcTRnw5whX19RdG3Zji5xttQqG2TPmOyoXxwz9GHYj
VeVB+mVuVbVoxOE+mvC+XPYuVUqvTyuVPgBUFTBOj53QudPYAAwcW/FSJWKNgIPLSLXOfmdtFcT4
fp2rvlL2rsmJv8eUUBd8cVOly5j+ef/YSIyiPmU9vIaclyp8XMzWg3hfcVLTGRd+xWWQmnhi0uPj
JAqX1cK+tgc58/foMe4W2Id8ziuej1mGRZJmeujsJ50RyYiLiKIcmwDD37Hq7efbQpddsO/VRl1r
gxNItC1DfF2GZA0VVGZlJbAnCpLGCmchVuIaQHh5NdvVGzL02XLMDDnsz8t7b+7RaFJOtwMKYklb
NxsbPvOYuIPIrP/1GXt6wC94h1n1ecWuVOfF77EBiUQptoaNvWCVz8EEt9xJG1z1IVIN5BomE24n
KyLjl88PNObmNU3KB0t2NptcF6F6G6f2VAgeODfu7YwYNtaxz8gPGHShQFLq1AIr30UmP1y948k4
ZxeDwdD+Bx6U7d6vEtoAoEDP64bmWr3/wwjTcal2N1m3Oyg5crhHnB7TAegYMgntUATv2MjPx1bk
33H8D/uW0qviENedpoXVt5IuVOleSBQwrJfYe2btHBYPXCjC9g/EXk2TQFKa5UYNszZ5jnI1wNBM
Ukf/1uFKLUHEGnCckoUuZgSfg93E6+hGJMhNOy6afDE9riuS6fkWrfPN6acqPOWdj43JtXUlQZ7G
LvomOS4DYF66hOiBpnqxl1X1kvGObcfQAHn4kFO8svZCBEdW94YSj2lybT5lvz6F40JfqeUiMLaX
RCBpb8ydbiFNB+tC9CMpjDtkFiKhfV/z+svlu0NmUXvXXcIY57VZFYLc95iBRxUVyJq19IjZlu52
2M31sL0NL36QEqEXkcQrS63NDPBXODPEGuBbDPWtLYN9BDOiAEES5o59Cg/40Uo+KR+9FNwkzPOF
wHBhr5pKe4WAqRklkNj7k5/Dp/Ku4FielL209IwfK4/x1KI+SrJLiGRFByUDnYC4NEgecMnymQXT
rzC8NxM8hgu+Ea/7su8046f4UKbmhjDamVDuQRVKEk/BNtmHAmLDp4nnd/X1v9GaSN2Er7Qer2xX
5oNGxEVzLP/rqMRpc4Hd/NhN/PvH2jslZVkh7qmoykLCA9mxGwqZ+6xK0K2zWGmTZQmBwXR2Pvv2
NR9bMJlptNo9ovOpYw0My+j0VpUfVQ5a6VTnUb5QY1Tq0uTvQoTEBaYftPEthDGlYOUmdS4+pmuf
9jvNp+opHBYeS1lSooaBSh2cV3DLWOT5aPDzlnF8cjthnEoDsBI7amGM1VP/Ri++FgnOhZj8/SdC
FRXFqxc8q4hMXOeAJ3t4OpxE3eHQ8q2DWl9hHiglcpgQfTpFaszt39MASc2b2XerUG4o+UScVv5D
KSDvT0EzQnLIE2Jrw6jSZQTm/E1p9z1E1OeXgNsUjY++NOtrcaevvfSlLuZqkA43/5U7ppTey/vk
0HFGLljKaK//A/FKE4u5NtoPRsuTfKs3UeDHSVhGpFu+q9aCnFURM7dhZylo4xCBj7VWVegLhju6
JucuVpvXTtN9WCymLRVnBpU70rGZTBbEAbtKvBCEDt4Vk7X64FaAennOVgKBEf6PlhdhPPIimIuz
vhEfBumHP9d2ORASkPrVO4DbRfl7vFlYZdRP0bmrXX3+upzw1HBOkPC0BVKcIijQCOnYwFFL6qTD
TRn1OzLfS6TZwgUcYTryVWW7KuVKC2lweW7+muky34t/2SJnK62ags99woWtWXNM/LRZsfei2Ft3
VPqKKl35cX6pLaWCdqFR9WEx3GeMlD4Msj4u/QtEz8/kQTjpki5SOot6Hu0xA7CGnaw2QXtfId0V
bUn5vGehSixrmMKfxgaa31Clb6Qk/VxfSVg2C/TeFTPcqHTWYCDB5hMg8eAwQpivpUeOOgaRJcJH
yiww+bMKUVWyJMOSc9BmqSSgWYH7PAq0Uvwed2uXEj+lvPy0+9GDisyup6bi4snj14xzAGB+J4V3
omrJjy0l3xqg+3/5IzdHQ2O/X6zePuNfeHK8F05Y7NdCx5824wiv++Zp6updTBSCJOEo5FR+dhOq
8b8aPbmnQNNTSZGxGHacs0f2BwozW7p365E51gELr6Qhiclb9g534L1RevJfnUmVbvdqZU05fFPA
NKLTsBGTxopZy3uG87KP9hkgk72CZChLmIZgyAQBWiIYHDeFvwOuisVblzuYNZyDIUEoQZf+1ZOM
eNS3bpQFEJR4gKYM1w3J/v/bOPmViBimBjYtZc2Xy1zcMKyzQlDbzaK37ObIt0yJM4DBAg4s6B4S
rcS/bBFbD6idpqdbo53eMY9xa7QEwmChpDRDSAdpM0v/BVE801K8LxSLlrSmsqS54V8TTtLNu+OY
BOCZ8duJ3Di8jDp/yV7plxzylydYnJHgAh8ClDMJpEqeh2HrJX70WW+ZuNVBiyjxNgZrWNvMhD2Z
15bhd8ZyC9AI1E1aZhieWcnfniqICF4gq4ZxDkuA6N3p4+bNBCKpAcCYdnooji1HY8FmVNoSI5Yd
IwwqGchx/qN8X7Ym+a3A2uwbzoPMJZWcPH2hECUIFy75wFZ6jAk9Fav6pZ//5zuOMUTqG3trZAr6
su8UWpaynFH32Pq/pz/mNoo9Yeb+YrpGeXivtekTswJYbw2/X9E6DhuE9rOzQcPR6clmY+lDgz/z
hXxbxXUfbOBmOuppqIXHmydcp5Ig5HcGDFnO1wWbmZRbk75Zwy4pa75WmOGZLDcqHPDIPp/13g40
EORQjRmzv5s2Enu920LAywZqmONlGR+36zr1JvvVmp5koTv/N7r092xB82t/zHfScSlVzDvO7VNV
bRUvXcznyQaIqv8Z2HtNrerrbE8XtsYKV5VDNZFX1hU/ep+r5JD0E22OtVpxiLmYeFYBLrbvEL+F
VI4yV28bFoqHyPsZrUTcMQ5M3gpTdGzZtZr7vrHEMucwzS1uhM6ThnyzHqnTkhZq9HDQY5nmGHAP
/2OBwe0uFzkl+rI+KUdCHvFoGn3l5LikMVbM5rWvndCIVTm6twq/BJBT3gUevZE0lXww+ZZXvpmn
kw9nkAVkxl7O6pdf0cCMS7PxgrhpKFUQ0r2TznccLn0U5YcUbtkwG+sKoWeXGd3mDVB7KG+VmlZb
W9NHRdVTNmQMhkQ/WEWw13D5wpFChJkLu8eyjoLej8r/jkiXBr0FyI68vRqVbFF+ftVMhlJenREy
MNSbkiZpdeURJcz52bVKsJ0FPT+xtkgSG6ts4ZOVYeMMsjLuEEYcFDAxtl4O1zaa4d+r5Nbc7Zww
V45LB/lSqaFtlrBLWkG56ztAHiLa90TNYALGwlL+XZQc/5OdTlKu4yz/w+dXu0tQEtsyoIyB2bFV
zHC2m97XeEtc/MPxM/0ThgOVEY7qCE9MhJbB8BGDaAFt8z2XcWu4sHsBb8BbN26GFkcwTsWiGQ7S
KFRHyJuQll3uDrmSKRPdcja9TlGej1H9zIsVO15MQ5QKnQrwacDDKPfVCGAXoBWWfaqGlwYTAxiM
SGHm2VLCXdfuCR44eo+q9K2ng6l3hWpMn5uOCOhDGYq76hpoBk8nxrsDrbE2TfTT4XmmaVxiSSWk
Ljd8olUZblxuM+Vt7N+D5fZln54S/KNHQd9NxKkO9G0IEVmFQHT96Ss5B7n9a1rInWrePU8D3QgY
2Fluj/OqHqtokTCvjtCSHku22E4c0lFY0Ifve/CSBWzhNuHgLqNSVrStvneDWsudim+xY2WAW/dV
h/fgmUcBdicLDii3CqZNE62dPSIz9g3vYmJ4lWxjE6pgsM+8dv24/WF9oavPXmdfaxSJu7/VYgsI
vxHQB2iH+j/o2oKUe56pVj/Bmjb7Wph1fOaU2XBVBeaa5gWDigu1B2UwowNDfaFuNTfr0X9oLu3p
EOFp5JkLNUanMFOM3YOkAQBYAAzCmZID8cR7PMUns1ifiuyjR2nmxbQXOWH8+svIslmbqrhYlFLT
7ZtgnCY+8BfEgSyJCOuP9+gvne9bgjfXLSY392nfxbovqOXtjjqSoW/4rAXGdtjeNIoQVF1CP1aF
ADIJtwkf74BSAl7P9NQhmnisGZmtwrmCQTFE9eYdj4KBcDJlVrdropcCGGNC3Ywjqw1qTNTGK5EF
eFOHk7swMDbRQyJ0g6+CL82pSIS+vBLW/52HY5Rpdjb+CcIR0Y4taJMtOiP1ACGKkmJrAOa1tb2f
/7ZubYlG1KSzMDM9FEQJfrJZPD+vyTJuOwcqGOis2+BK
`protect end_protected
