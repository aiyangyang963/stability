// unnamed.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module unnamed (
		input  wire [0:0] probe,      //     probes.probe
		input  wire       source_clk, // source_clk.clk
		output wire [0:0] source,     //    sources.source
		input  wire       source_ena  //           .source_ena
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (1),
		.source_width            (1),
		.source_initial_value    ("0"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (source),     //    sources.source
		.source_ena (source_ena), //           .source_ena
		.source_clk (source_clk), // source_clk.clk
		.probe      (probe)       //     probes.probe
	);

endmodule
