-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
D37GC7WkCtKgibDEt4diktpNnZH0llKDWnn89I2Fj7XzzVNBGovoPSJMnRufmvq2yFBhJn74lSwG
cWikzQRfg1qJozN9jjkYxcMjk/MDINYzeRKB7mtG7GGFq0eb2QbdMPPQKi5x/PpW//0z7aYx1EV2
eCMgAuqyW+G8tADhX/zPZRlbG4ebB/HgnaH94pUg4/o7Jda6+iT3V1SmIfJt8tUVjkEVwT3Fl/K+
jNt6gSeOvOYRGFvHq8v+qi6MgZZ/vCBUsGmz4xhm80iH8MyNNILJRRMpzmbUYpQmib0ev6NYov+w
+WFDIJxtFrS7CAr4WI74ztUhjBTvrbyCKG+r+Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
ZWbeutyfhoPU+3mA5fugiRthg/OMuwPrFZNzjvmWcq4W7YUGQZIg573K1o6XxrBFxYE/KwPur9rW
ed4L4BbaAAAf2rGvlluS9MUdHFSAdwXf18kKZAfiIOZqIqIDAKalePXPQmeh42rYFHcEv6x96WBw
zSgq5lYIzRlrJxsQv7kusqlCwyfxceVL1HnNHRSvhd0ThgWOe8/ChfnY8ZKcuUxokfjhWoVlzF6h
UqwaNkRHJIfpQOQamWE7O5FgdDgE+PO/N6qiAjPJhAlg2Pb2rx55lRDgsrLEJQ3XHqOZ+aXKKvjs
7+MqL2RNZj4MqL56h9OKA39Pe268erBunExI8ZQV6BLXN11F/tcGW8Ico3s5O44ASmji3lpW5fkl
auVD5pJjzPaP6xeGBLEaO6+4TuRakcdv3a2uAV8vdEoCFpsvC/3+hafB59NwtfCJkjhYe8x8OTVP
jiLvk6JP6+vCL5YfQ1/d7iZwKPIAepu8gQ3oIfgH35/POTunETBgKyKRqfvLDn9kuaEZ8/M9eqWB
rz4vyGkbfc8dfGWR/dUDajM3J3thewD0htui7x1bsu9sIk8FtAhnUxJbp/1+KNNq/3Mu6KzUpQYQ
ZbJ9qlFbcluOlOO2fNdfEPczbD7KwL9SzyeZkqLy40nw9akhd1kuv6d76B+hOJL7CuhAmsuR1B45
WZEN6mYIC08hKXHurhqW+xwsebqSGIKK41IoF6yLRfsdcFob3YznNQBXLyVsE4OKIl3xtUICYZfM
oTeXAzdZIuA47ZdE/nTqxC5m//VJFi8aSVAh6nc0dejna27+BSaMh7M8k/AIHToVQXi67fgNa91r
0HPTfOUE0oLJZUEMwXMLBAWIY+gPMYt7hJo8UDulUWVXID2gYXqUEcsb/r+x+UPf7GmwrghJjFpx
RK6LJctPGE4gluZOSE2GF+1Oi2tDV7pVCcnuHPn+Ek5jRkerONUruuEHnOo16uS2ncXQqK3/Mu42
XnF+jOmh05ynixXI7zwBAaWRyc7Bj1zmE0Qq5MVfZnqeQ0QreADT3M0Abhfzz6B+yB9ullZ59AQR
2YauST8wpKfnLFFp3mmfEcLctARr4UZjY0rky8if1McNZ/RFgkQCfHHBLyRCNa6HOYBX+ikPnqz6
wjLfLZoul/fzetAXgY1e3kndO0IgF22eshFEq1bd2XvtQG+Tc14TacuJ3sUqiNiLrPmco31YfLKF
YmG/Mg/NMprtcy6hv5vstdGjHwZ8wuUpwsQyjYxy5Q+T23rg3RMCeMss5C5HY67YO7ECmLyEbb45
tbc9TsO9vF9fiqpl7QtIWE8va6H+KJ+tWh2ezg7e/erFnzWA5xRpL1SN+2bCfADp4VyBSSIJwSng
nzYZxuipLMgoxhM+deUjgXHLw78mE/wKc+xKKHEfzOwYxAPsxYYCvGkHooGFWMLaMx+SJbzDRkK1
d115gzLlTuSIadxHrAak4dE6XZf202fFeBkVSGcfOsINRnjT8lsGCevM7C2xhK6uBxOVSEh4iV4Q
V7BGDRsn0uBJsMDz1PQ2WZ8zFAVEWLqtl9bc7SX/KVdQ0wLGuegW0754yPo0gWZJbrRZ02ndgZsb
i9ivAZeHZXhvDNHQsAsrwDFtKBT9HGG2WxCptRkhJKvFIkDc6si+VKqjGh+bxw8EEw2F4OJPiuSW
sl6KapfMwPdcakkpb5QdaBs2EDzaL2+H6Y6WRbeNpBygIoNJs+QWxRECcL8/B3VAAfxh9dv51jaR
Tl1tJQGOgeRhlNxOdTQ210+ktJDvg3V9bD+qBIUiSySkwEYfustxlEZFQTgQDATsxbcOLKCCyqIc
rYCZ+ShVIqkkHkWw23AewBnQHVLo+5RKk2IrBW6DlmvRV4SEjN+V4TlCI62KrCZYZ9AdtdjwDo8H
lEsgsQFsro1IQwhgsq/f1y/wyc2PVwjiSlD7DocbjEzK19HGV5k/oaJ9DTp7xZWCfYrusEs2d1z8
RTM1MNAb+x+8oCPPxQ+vW9Zvc0dly81PhAGEfPwPknaUcJPW7lzj2Ceswxh1jdDfD39mv1gfi2+q
Wgx3K2OUuKop4uG/9aVraS6tvuTBpJEUu/lUujSqTME9eTc1Pt6iL46+3LNC/RzANEDMVX+Odedv
Ozx+9opztNwQ8vYTvefLKWwL/05T3OL4XpXLBKXHl5aQFYznDWeVauR1qBc/zYelgqYQKE3RV/eJ
jZcMdZQABK9R+TIqp+CeEJYDDSajSl8/GF9NY7ao7VBhiWpfElYm/fi3NJ58q32KuBejlOsMI9ih
wVwfKAssEDoRNVdTJ2e+F5IQidmGsbC7VLCE1v3qsu2Izd5pN0b5hrVvqgPyvLmmmCRkFWvaVKg0
nUkPz8Lbw7NKeFEPSDmZAxOvG9aearJi4uHWkV+qcSXRf3FFB7ogdBRcaGVAuu3VMOM7jHnRA8SE
gngs+j4m541buKO/T66B2pKM2p+F5XqJLIXIaiRdjZEAKoBKvOrV1QWXP4S/YvWlMrYOzVOLPUom
xOvKlNtB/mcUiyXUojImwFWd98w7ugyn0h6o5NC7+xChg3HyDprx1NcUWaGa0AoO8Ya9AF2Y5fmc
mItTEAZ4RIUJM42oWFWZGhRZVaaDfrk3cT1fkpyqSmDi2zzIKwXY0XB8NkoyBaI3+FIMX/m9Xj6M
5udf8vcwgQlHj4h+X+AuVO6g+wnF64o4MSYuXIcVTHV9Ej1/iXPGgmUkzcDo7DnKrmAfZJQyiwst
Pr/WQUYEJOQHGkEPlqp1AgujZLMUJRJsxPUkmf5hZpMxCes/hEgll33j3mBZUU0vDXjG4tBeiquz
LofRRvHnL2gV+mUFZG//pf0mU+AmylwCo+Y7SLCSZMk3/EVjy0jL+wEcntfK5KmecSMQFJImpzFl
bKudyZWwrP0+3exEHO03nXeusWTB7aUJCketOKjbklZUbkmfJtDVyPp8xz2p4tLCrl+rm1p7IeLc
rETcbqj5X7unaofoIJwyw7+8kpJla7T7l/pgrXWKgkJroZFS/hLJRlIAjvFoNTWqODdqw8uN4iSt
ktCbE/puc4QDsOzVTEUYlfkWDxBnv1PRkkACYFX+N5k18Kj+1E1VRZ094O8Qxea9ytG9MyMSWUpx
7ZJmYBVV/Azmjrt90jY45DJE4JTZ/AEFwxJar1w0kHCGZogxg28XKtE64FcE5lRu0QUFWn+xGWiy
7kPPO6EoUrL5Lv0lLmpS83PcI1gW5Grl56B3uPAD1/IXjqTZgMJhn16ybpKLeKf1WyL68BLfZL/2
+D3wU84jTdI/WoxYZxGI+OG/RpvDnmUCF+i5lt7wG/HWx5K6W3NM/ScTOTG6cT5oP/G1LDtpyrq5
RMrGCRHGFQNnyOmfQ+hlaeHuDvtMEO78dj+hLk4KSmXg/xG9ub4ajdFNA6w2bbyFWD15C7El3COz
3OAZyRMMFujDU/n1Cb3qhfL660dcOlikpMVto35Gi29ZSnNaDsGhUhmUJZB5CpmpwMJOHkBHewAE
HAWwb0raKLPFokbDHJOxltuHqDuvgDpNl2D2ZmYdstqBaXJHtLMEcEHKhj0bQPlG7t4Is9r24SQI
8tTDyp1gNH6w2QoTYXgm4WPmE2XlOBPU+rDjnX3Xv7TCGxmVXs1Lv5AQp3jwDFVDhSKOl/Jf2VnS
VQ4StFkQyivCNo0PYPE6yqzyvkrDSzwJq2XljoJaVt6W38i71SZVdlJkJ8ZwhMFuA2JOBMfIygKd
OcXZbe6zlSqLCc82rY/xypvCcZglrVELH+svY8lWfu7z0eFf+o2O72S7KszR1YAGOnhWJpUqdlaT
HHPXRYFJJLHt2DOhSRIpAHv7wSMp6GCiQmiUq25SrehcW67HRjiMz1iy+RWJQhBmgG1PZJ3XS1gq
0YXTZhY/FSo/le0ErN/ntE9HbCOMgbHWdtki2IZMip2pb6YYnzO6REIJQW67RdEK+OPDA0uDxzC/
AaCq+7He4jVaBKSzBERrsLxX1R3b4KxOqLR7q1PoaibJDuASz7+NgQAxieAHnxEvD5OnIOp3q4c2
3WIMlYNcNBvIuZhd94e0t5hpwVN0jb4Imks3jleqlns/KWPLzLI6zTO4Enx8K21gz7BnHT8AV2l3
67hmJLOfAUor/wAaaMiHoqLl1TGazXNvGSufXQ8OadpHWlSXOZ5mDHXm6MW9N90sUw6XfI3WDWHZ
x4OP5BjWPipR45w4/DRPgVqtE/UGystOwopkxQo08++aU2/5NbAhvujCMffkUFgtgi4j29AmkYK5
bNqKUeV1ICgeZXb50Gsh0Vpxp7M6bJqp+Oyof0SRZ5/uLx41w+d/TxQpcPgqZS6NdZ08NSdTdaLN
SVUJt5ZtA3OfTDpBrx0WBt09lFMxWfzCTm7OlPDJ1sL5viu14RPANxZwer82qkftJZwfKzqZwFHx
v3vuaQ3HuYmtIGEa/BDnlmweTTY6M0+HiW0tSTXYPJpv8G7qw8s3iaP1atdVKnYJ9nbq5o9QFnAA
Ra8/Qwt8s0+srWIr0KjVocYejaMw8kqL539yq/ii9ReffAA2fBj1wjx0kfiI43iZ/rGdgRf1QO3p
YffFUWdfXaY0paV+ml15IPlVYKPcF11978n6+qVyhSDB1b2Lla/WdQQVK0xECLw1/PunZtcwHsXd
R7p29DArpx5KYpMAT2Yb+SBVO+gMQ1pmlaMbIyQVqtIXeHXH7at1IGF88bZDdgwJBb712jiG2drk
ElJM9+cQLteEuWert5N6BIDXlLMzaOx5XNaHuZCfJ66GPR5fjOnd7mXxFqd87X6IdkN0i0ujLSz7
V0hd49LgbuPlGm8JoagvKqFfFtHzdbFxs2+IZf/Dz8KMaNAlmH4DeF47TDCUshAd/dbQKf3+DOrt
b+5V5m/DynETAkQa6Wj0GuiMpbNixXkgxVzxvpxVGA6OuaNH9NmLWzBM0//o9LHG4YaVE3nIuf8l
bPeF2QiTvZrcxzVeovGnVb1+mCDAyV6Gg3TbQXmpWnTcqLApwYoi8tX3/m8c+78rTPOvWFDUsA2z
NnBKYIk4qk6YBYe0ocSNuWcq5BY65WdEbz7JuB/MyA2UM8HiWf82xhnbC+M8lBWk/17XDeSkaQuE
9mF6b4UY0zkmjO2TMbhixGEtp4f95ZvQrDQtPVv9hdSn/QzlU1zC1LCU1Yg9nty1v+9DhstXKFuR
M9yezpdD58jciyPDPR5igirg7ITs3t7iNTjeQ0UdS2DIOUdI8ExfpDsMoPjrAbasLM2yGLcvRDab
SkSuKlqEATVBOiCt6VldFiFqtUUu/T5jKPKv/yMd3e7KE8YMi+nfiV/StNJFPX2C9FWmho2/56oy
PMjrifgqQ1Au7g0y8V+5FssADPFQn3JAV+itilQUxlssWBb2xhWhbz/T16ophTjDQTeU0b62EmBH
mnqULMeoVD55pbLzvJspndD0iv0pW7b9RGpd4sIOUSK0QqxLELNoyQcOQqaF0cBRlrET57kNvdTZ
YHQ7MKKAjur3NCSNS6/Mqj5plvO3kjoiJanWVV/3LB3oUJVRdYVVoHggqVz5QBeKUKz5/FZGcbgG
rdP8FV2i+FlyQi0ZqRJjCimuYWSVcGAJl6pgMtZ4eU2W0pncUeP1g09gFihgysJee8vFrpUTt+KN
4SjjDZaX2an7YTkM7pxLreU/KW8FLzRyhpLQh+2TjVVYLMDRfJe8SaYATFQZ/YpybDONzXfzQL3Q
TWYmfZsJNI2UAtMuDH3LXYkDigZXkq8TzUQB+2LKI/djY7Mt4PBgv39T0RKzcVtryU/qlvxeKApR
/YK1q/LYsO1F0WsURsaYiI2zrJnMsffLBz2fvZz/o46aD7mCxOQfZlsJlaBetY1VyEZlIFhJR1il
FgvlmeAj+oNVFP18SNe2y43vPkPsUoee8nlK4VKLBs6uyVB1y7MKywJ3PwihVCFzvBoSJVI3TCFv
0MBCAEp+zZrS1sGpVxGiaDjrfFjdB+BwB8wCtceDzXbG3tyLm4qP/d6L5nYOm6caqk2KiSHkeIa2
6IacC/izXDtFwxhBocAo6kC7bTcyK9NlwvR480nzaJMdTvTL5m4yyrnU5P2Ovcjba/yOHuGroHR3
BplfvD3imhXDTdnlt2juGEag5JJz8u2m8t17Blf4MWGvSra0Z4RTjcV12kNS6TB8Hj8R11Zk988+
nlBvJHKmYpv62YKBEsD8HMmNepvzwABAu/a0hKf5tOBfQdo3paYTXaCxNkj/vwZkKqhDgQhkEYaT
oph2mhUCY3C7oOnd+XE5Y6MbIR6RJvbcpHSohP7rwH7fU4onM6JxcI1L6/mDHFNQ/CSm1f4ZVEMh
OU3omtcBLu5RVVZB2TWNaXkvsC9TRG/t5sb11frrXeLj8jizqw00j0QevmDmaKW6LCFN4ncZqtvz
mUzSlOBpPAOtNdiMNjP5JGc/BbLnda1GIxuztnV/NrnW9tYKWa110UPTmFNbL3rrNSj+DrcqeLw5
9d4quw/AgIlI+MRKJpbSjHYDSukqzTj1149YfO28t7sBUbfBl5ZPmHG9R02p7XCEm1bTuqSsR59r
c+I2pn1sfMKOpuuju216BAsuneqKy558Z/+CV8i+jtkjfR+D49E+e0Cd+o0mHUfbhHIcX9CAe+Pu
uN31E2UQHVUYFUSS/lUF37XVlGLiDFaDd9X+JfD5yCCROKA/YTpYDqCYxrcImC4bzKcIjqQaOpcb
pLvb5y4O9HbVWe6UQrBh3l4Nu4W3wqv6cLAmkHrJID5wNulB6XiaGcyYGe0CuYuWwhKE2//jaFw9
U+txy5vzjR7CneNpoiR+hh3OCNHvoNoqXWexbRIuSKcThaR15Rsds07rgX2EAXUV8eN9yQzwiAta
R8SFDZKeVKwU3fYqJzeVgC13tPra/B2YsR8wqI+54h2r7nxQ3Q0XfKUq56Ss0F9LeRgFQBQwfVPR
u0UIyrIkXZRXlIOMgdldum8WvxqekfevXmcSMXCa63KBNY3caGEQuzOw4buGONOLz3hzDklePG/b
u2OfOCnyfT11rhRqzmLFSUc4ibsD+pLwQEtND9q7j8JX7/tYXAca4t4Z3MU7x0QxJhDsMw2bwZWo
FnAD91xB8QqP8g6ST4t1htmOMR8jkb0XdD9iRLYb+baOb9EDzX8HwaA7icKx+QQpjjmrGcBgmrJM
w1gvMjffH4hufh+HFu6YUTmnugh7/k0llO8FYrdO5pegLxLwRd0Ub4eCy9rRRfJn8i0TtFdvH2mI
RwBOZ3I78EbkhLnLANCvfJn2m931oUYrpjzanls6T2xVl0Ek58NoOMVxKmydlWa6svJ7CUZDiz/M
4yL/r/XpXb67gtE5DZLqY4wgk+x8MxMyZCmmsrB2esfZcwJ2XidAyK85e6FjHeMxBZe+2VMdbx6T
+pkLD0BW5ntoVus+OPvk5e2nlgFa3IkObOGd+Yu3s3/PlH3v1jF0OlOzVE4Cpz+yIrH9kBIREKnk
L2MRnzbELBPZuHuLBWSEnD9lDDpj0EV8ud2kYUnxXqFLr29CjkvtRASV1dDM9at4ZQZVzXbV1xLY
sD31r+f9rypuizlo3hBP5rUhhle9/fVSWW9UvZXV4RMj8qHABLEeOzmq/Nn+knMz05TCb6Iks3dY
Djnk5ilz8N04vueK+tmYSy+8SIKvp8/A/4Jd8B6KrlgIcUhEgdf6iFBmJZjFwCUytd9pr6T5d3f2
q5ufkxyXTg7tQjjXtyXvE4fxPQTC+r8UQWDfqGPVtfs5IY9MOe5VnPtEglY2qdo7fufOXa4tgdHP
I4fvknMGSkH9gPynUh7Ptm4vLVEoXIcZW7V47zhk1emNeDCwChOOvSslsIzwswY5NkRsw5J+DijU
2o4/LwdujVqWLrtV/pHsKztVm8CR1B1fMv9VxaL6yO4pr4ykgW4Dq1Q3p2IkKSCB7D2MZxDuTqwz
A9aU1b0ZyklSuWcQzQ10esQazEXFXtO5zb3o+u2mbZJFXmb4CU999nCoksXOjLuUYpyKVBExwOti
NARX5H4OBSe72bQJqQbcUgBSyt+TKrxsPAtXMoyWVmdNY24Sc9g1sc0aipz3ArZ7QlIRtOk4UR2n
luBKQJGWgX9wQ11u1Cs0O0dypzEUM32r4sLQ4mQS8s0L+TIFbSzJQRJ2aHBJBmJ0AgeLFfafh+Pd
oOnLHfWuxBYU+SUfACRIYyFeUrctliTcm7ONbMvRL+DDB8GADaq+6BE+V66ya0pmFzAfNkS8hMH0
NueETYxjueOl2vv6L8MELDfSRZrK/JBZbruX1ePX5gutPjRr4N8W37Pj00N0prdLupZvnvnQCsYj
P3H+yIy2G1/Um0Xk0ITljdLkRHa+xY51nE+aGIxbSb3DnJ/xOEl/uAKN9K5NO8KpsUbiYGXNaji1
s7vFsex9H1knll7Wiq7vMqRsmfdC+9LQtnMu7mC0wnIB524m1CPUClseQtI5wUX+8mo9B6gtasTN
FWr0KfSUTIoggAHDZhlK3gFRFu9pfj2OJepJHiMp3J18k72q9EyIUBwjPn2DR+4FJiaD742qstv5
jenUj9myj9VVaLWpbyUEuFfi9tspxkxfLfjme0T5SYeYuvTvAp5Jdph7o1VPLJKIyuKhodZm5hc9
GatUxwxdpzXVq2cMR1AV8pQY9Ef4wLnd8wPI6b3HlwY+Q2M68//+N5XVEDlsT1LXCLYB6p2twmSf
Cx9LNsiasjTai1n62KcFJnEX/Vacey4LGIx+7OqaFYDfST129s8AvmEN1cw9Ffm2yVczj2f4131W
NAKlEJf37ockUQpGdf9Mtrl6eqMPg7JXpmyciI47zYly7YeXK8LN53vrwyn1h+/BwphJtvptbYVh
mV/7uINfzqCRajQitGuv6GwlsHBHBNFb6XNoXSLjaEroQWGErcuLH55Xpj371yk/PtgreMMJmz4Y
b4QlJfvrmPg2ZswFyON0/0ISgTejeS5qaTm5Np9ZdlQH8PwL5VDC0evEenP0A8SSBLIwTGj059Lf
NORHapInHffhFqjHdzYAvOvMCSmDt7tsmkWq5j/mKd59vTLvb966AkmEVRhn6LPWvfKul19iiFAT
DeIsAr6t8elo1ObgP4w9go9SFzrrvn7fvvhQnakW+UdsOKt3hKk4n9RGqMhv5s1uwudkIGfKYoVA
hM+Pji4REw14mnR2O/B6x9gD7jNv/MQO+XVxgPAn3B+HamYgH80ibKVH+joauygHDhRRJJIGCT4O
lUH7pma/5OotjjmV3Ay6K7TrWNcdHNSsAnl8xWwzGZS8pOLyxXwAGlSluAb+oaZb8fUU+BmCt5LY
DcSPu50aHOZ5u4mMTHEJpj3PfUE0UjrUseswzSdZ0oQGJWJOnJTJ1+grN9zQ3BrGaI0+3kacCpFk
grBqAoDnjsQqTBPl8MRynNGO2x01YwmH6gqeEiEmJfw4B7lwhsfdgsAEreqiJSljmRTGBiiND1r6
1JioXTNmGh+faFylpdppR2wqiqN+RQigWaZQknxRGHPE/MULbq5o95OXZgKa8ZAKMHMC47azkJoh
PL98g4HfPNtGJgfm8+calkd41yIyh1E2n1XqBftuzz0bvhPbJm7LaaIXwjwjbel0InhoOKoUX0Ds
y29vXPaAKkbO4MECX7i/VGamTdQrWx7LIzoc0eju76Yvdg3n+R1YZD5N/fOSwvY6ySiKVGNzrpxt
YgchSc6JCya2m10qON6UBUl7kPNgz8YYF+JGujZ9Xc2FgN0NujSFw7Ay697UH9Mi7MZvOkhrw49u
Bh42+exNwZsSsm9vigbS8SuDeI5pgR8bqLXdb9fFcUopdBT3xvyVNj+CaM/QP1MxabmATS6JhKmd
sAicDLqFvE6LUWBnpPpMnR/deUlelruQ6/UtLwL8VXxUT+C6NYKjEH0FWzYGs5hmR5D04IOaq4/R
YEG3/6+VlXfZLZUFuqJx+gcfAAGZc7NjeBKMbFtqfNcgq6bWfuDFnCSxk1TEXgf6jyWaVlevqXL5
vLcjdtXsvwOwZ2MJ08nuZAxQ513bCRDC+nu40JD/0g7yeFqpx4S19TH8TgetUUpspCIJTSI=
`protect end_protected
