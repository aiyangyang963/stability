// trouble_detect_enable.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module trouble_detect_enable (
		input  wire       source_clk, // source_clk.clk
		output wire [3:0] source,     //    sources.source
		input  wire       source_ena  //           .source_ena
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("troe"),
		.probe_width             (0),
		.source_width            (4),
		.source_initial_value    ("0"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (source),     //    sources.source
		.source_ena (source_ena), //           .source_ena
		.source_clk (source_clk)  // source_clk.clk
	);

endmodule
