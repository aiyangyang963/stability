-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jKZBJbU+o/7n6xjjf59QkUsb0tEsKbWTOoXm5CYLMTypWOWyWEAbEtYpFyLWdcuiDxuzTZsMRg2h
PDq1r0wcLSIfzSNDcrnQgzSJC8FYkg5emsqPqlWDFjV4Cdvj+6u4XKnTNu+uUmCMJyW1Q2N4FhFq
FbIPDwHuU8c3yob1nr+YC3g9ln+YXlmoODj99NBuAF+61UHbb0iHp6uuLHgZXDIFcRWwsHuwDX3Z
I+rKxoM3F56JgZ62ijuhv6tau0f38Gyc20z5uGlYkZQjanKWnoDQev60xcXvfcvUxWNh0LkM4jaO
KdWfO0ojVKsjsfixU9QQmmeHbzBvNOxKGZb+PA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
eNLpu9VmCpjdK1QwfuSCrr3pQl1o4hdLo1b4JOovR1+W7aPAZWZ4Mf7RzbRC404wPkpp+C0uVN5m
9qzBCVjRaOjxpICJZyWGLJLOsrx642Do7c1N+xdVnXAnndrXexg4cieGUHcfpAHjBVb3EWZa06EZ
JNKCIsm14YGC/A7uP0zSM6JIiK1tdi2RMvugtnrX02C4Y+GGLvRDF5y4itBgCny8OBnTgnFp5KlV
1QpTLZeytXLBC445wq4HNOydYdPhHJM9cSQ7dcsNv7w7uTJh3F1PJzX7cEC2XcGs9EU9SrCvmrku
vsMuYlF65PBr+AcUxUbEwWuxewAfId/uvDfepQZDYbHyb735hbETxh8ceXqlGMPd2BmCyF5A2qCe
nJ1wN8QPToHu7mwIIoTBaSjCCkT25cT2K0RS8qKxYcLRwcINsFbNk3H8CIv39E1bdr4wHsUdfGCh
9Fh+g2TnfDw+4pKRwMS876AnTw4UHtcd6kf9G47bRAjMxnfPyUSjHd2OmdB9LPWamHNZTbFzl60Q
tBNA2IQx9PoElKHNKgJWjhGfoXt3HRKUBLNHgeU188/FtXAxNBy0AeiBR91eptyAAHOUHZRXU5eq
Yrp7ZqWWKQRPrXfyW/OzR7pqwUwuXrU21uxh63ZvgfddyeIQoUlo/6a8Px+ndm24hbjw2RulbqSG
Fmy2S+YUcCWdKrji+dZGfPrmF0trJy7P5uAkE+pJCkMmFUbSSMeoAG2jEVWIRkq/Md6Yuxes/UPS
XprAFtHXZIPq11FPPZymHq3GSAR9o/jLKKRRv+PY4N/5/JNG2RBHXgE+TIXrLJVunnG54R7HMxEh
w+8jROeH6TZhTZeoz9JX2edCXQJBxyAwtN53D7LGl0Fs9JCjuaKQp6QhKn7z2p6W0zx9lmKwpAQJ
WrxgE1zvSfwMeLdmFXuOey74GspQH3LFQGuTubf2sl/1QDHiaFcsGE2latHuH9XV1WDIKizx2Omz
jQw/JT5Djpci/3cQPmTie2jtJLgjeVbRakMZIs5kEEaLZi1RhKeVt1pF9MAs2WSdacQKzK+Eerfv
oktxpGGiJJo7c5CnW60At1KN5ibqwnH/Oucv3W0j7VRAaEUF1UdNhj1VJtEf909bxblIINHUgNoG
dtkvn+m2IGP6ii/GIMR5p4ZKWoEfdLZJZ9tgpcgmfZkQiEA4E+JWjqi7sFg6dt25MVx1FSDKQSqq
TM7e6W6U65Sa6JeW1BLdaq8j9ftC3P+tKm1I6Rh5NYk4Mwydxa1ISNlS0eHy2E2j9/KtHiqCbHZa
1jnYyAALCzMKSaCB6WMxVD8U07OYhfwSbfQIy6jYKG/opKMHwN/xcx/bg8vCtqXVrUv6zaxx3Fd6
b+wOo6hncEY37zmy5/oGqsKSwwQOGdbpSp3p6XLwjg2xsNTsARHoGr82MuWVgRWQBgW658/TEjGK
x9lFDP/cAP7UpPKg6MBwkvv1GQkCqq6HBujIJrd+kO1Dwb7X0RWbK9ktJtak/5zxsh1UFXqpI1x1
xGob1m7qeo/B0jWwy2D9SgjpFRmPi5IR94tbokejk6AqNbOgqjgr6/xd8c2F5Zx2S2QcW9l1N1EI
LdTSVkochG5XPy5UCYuMDRR+Ts8TQpDjJwUXqlxPeShyhLwr/jvcsMBwG0or/1dTB2qEeuMwsIfx
dZTqygYfq1S4mhWTv/cbq+XP/yfFLehlkc6TUUO0JAhpPcxPUn24+/RJhkOC8EoTcpAmppzkM0YV
OJaeGflSgMnKtlvjSQFourD2s6t7xXZsuVjYKDqP4YmkotKi2dmyE68YxW6qS0wokNtxU3N5kjEu
yKoZ6buXgh7isWPNWOCDIJr1CXUxjmpzqUCwjQkKM1oITK9mI0NI0FDF+mujshthVVguspHN3jIk
f0QulMyOwmxyA3sLJLiiWwPF3NcRhCIHK7s8WwDH6e4M1O5+dQ46uHQ9hUapBTRNClUKDhtO4qCe
6jWwlgT6MIFqRjb2eDRDniJ2ibm5XO4wCLsUkke79CNlNEWg5IC4WKj4O0OPqknGM5R9oz5o5w/c
9KY67cEcxurjxIhhrluMzhv6mHaTXw64BcO7k3xtpQJogWrC1ribtTSo6RhyhO03RAQoOo0T6iMQ
uif5V1N9IIBb4M19zsUc4OyB0LVZcnlDogMV0Gf4R7Tyo/e98hymWZmfIjZStRmL8kz+NwUQctN3
NoXUaaPp0Ak0m25OhUI/7KjfDHx6vlk8hup3nJiv4GGeyPXOyM5WxeFxIbVK7/dubInE+/ai1KnA
oVm63ypZ9ni4r4pE8f74RceInERbHAFiKS9Yq6fOlrdD6KjXKLrgOkGIvpDWjccF8zZBKxyi3soX
lrGDAJoGQNQFJp6WqF5G+bNUomlgnwSfBwCC+/5d3A8zmZAK2Kffb1rgghiWtRY+JW32sfBrDjkk
2GfNWeHVwfS7youwPfluuT6u13YMnyajFHH8SoDvDRxDurSzvS2t0oClU8h9Iyp2isUbpsC8Q+/n
5PRkfRfN2zennRPqHy5K500nAN7mUD72umZNETOnvb1RpitB7QXZ76vJbcRaRwyXccNNnBQbMFzG
Fh+zcrE/XpSZkKHbYuIFR1kkG5AtIhhW3BN/gLsH8XdUoGm0RqV55wsXqM1z1W9aAEw9t99wWZfq
Q9TV1GnOF2L1Ie7z/RA2AnFudHccdgb+0CiLxhkrV2AMrcPTYpuOB/O5wz3HmL94xb7e+YScb32y
0njNbxNfvdeszAjT5XFu7YfEmeF9KRcGXi0ncCq6+HCwsM6P2r4iv7gNaohCrL53u4t0vummi6dv
EzItSxx2s8ADoV6GftCAhqtqDojYN8+MTBzjuvU0y1bDzCfePdrZG0KIAmJvZKtwD8UxE4Vo0P9S
JGxJcyVRW3zOt7TKsmJJOwSN1HbxVEUcscR6iqc7zR0j28rbXTSSf8HItq6L9wQDRERmYk0F0Lci
rSzEH6knadPeOCIXXDOwlQHg5ZoZ/isRLHGmTh7ywqLj8UyrNIC+x/cql5nKC4QjFYTZep/LZVFC
koAQZVU5gsamAAcpO/db/cppQYQB/vVfGVBCdMRpO5mPJwM3/u2AhQltFrxBPqqQqlOmpzM95Naq
QiYoG37LipdqyQfO0jwDiMIEfGXa+/KVVz1U4KejnZq/DSuAre07ZmpZpbtICaDZYHR8i9TWiRn+
scgSa3qOHxsPyv2cOBK7n9QI6tELdxv6wYYUgi+gotqkxClepCqA1Iw7efuLc3gUpsKd7lSA10dp
awwp6/o752Htk70M0wlMX0uXDf7MYcKk+bQDYkma3eUiNu+m9SREBIctEuIApU9ONpdinqzRBo5N
HpQQXuX/tb7UuzqmWScuKfkxWH1O9QjnY4BRjNINeUwKv55CWFQAvgBASFBeI4u8pEI7C1o+1UwE
yIMwDAQY4Z35vUChq6PgOKSMWWi87j4jqCv+R2vZRmroJ/HNkvvEINLM8OFt5o5zDYJPin6lfndx
+xPxl2YbOQBfuikevrbZmkqntwo9VwaPjEv3jnY2K5x3nZzQDpSWsVqakLctUoBbets/eDNOql02
OFTdOI1vUnGdZ6aMnXsygM2Qk8MXOVT+heXTRC/XYLmP+cTsttssA/MPZKqjxxaAiC7PCKhTZkHO
g5PdObFn9uAGK8tRiWAdtX8QQKJB71DA73DFslHU50tP2CFsF9JxVF33dXIMRBQKu7/upPoQDIie
XiayVu7o9IA21n3PBrOy3Q8/4SmKBQvCiHoyDdVZLqcjGgZjL9LpBmO5vaxDTZLiuFswxf70qMFf
j1bUggwlVipEUIVnxAyg8/7iJbsDYN7ssPBLAXDfXhhG/mQGGstVxt/SQ8IMnaMrJle+mrRUthH8
xv5VpHotaTrIZPabfBsOmaIqoRkl1oU7o03hW0qgsV+57gN21fTwujpw5xak6wGU6jC9B0qqcTzR
2DOtp12EmtFH1oTbPoSA+wu31rNtg3mWk6Ixwu/l5R37hjd+7lFKVRfCl253z0VZTKYFjWccRxew
2cwsvQAGId5RnWHdj6tB+6AyUBMY08FopmQFiGBG1mpuCwTccNHSQG7pGxu6xuuxi4o9Kzn2mDLR
RU3n9f0c2qvNndyEBfUcK5pNlS2JCrY4l4Xx8FRHvpnstj6V5Dn5wagZM9s0s/lRAPJ6uL0jyhLk
rsV/MDCY+sfp1oaGM/qaaIeTN2dJfoulYxNG9YU4zfESTUgZEEaIbPiHSrl7QfTELJ8SDCV3qpNF
7Jf7ryTc3Rk6LLrQLwu1X4f6SVkAIcTobQmZT88HNUNdQUCZT9W0wECU9lXj/rSAc7ijdXbJRonS
4Ttx7s2kDTVMtWosI/+YDzC/CpGKJ6wZjKy2NxlwCnAyYbKY/xfeL9xb2PPuTZ0oeQL4gORb4Cot
5D71KhXE/MCit9t/ke7lmAIqFUlJKPo1TZYdysDDc7kxPlttaqvOu218cURpmsyDMMuKt/aNJeSF
4eoAiIeT78JU3OjGOi/EQ+Pe+2onhNrV3jxhUGQYZUX+ic0GXzDph1cID027f+FIv5zAVCzVUnKq
KJnv941V3uYYw+bPohYE7Ijj0YCu9AZ/+9KLw21Yq5HRDfDi42SthOZkN9N6KNZ2vT0AU+LPx74m
KJyTTNtQE2lRSboMqDr4lhIrYgscJJxzAT/tD6I+3jqL0oX1aFuXtyqMXy3ihtud7OIbpENQTK4X
WSTy5fV4m6TQWbOuTggQCWdZtBONNvZvbu7zJJgtn6cX4Z+tOEqUQe2qAVl9U+a8JmJbSxT/wrv4
ZNMmh2QyPuHbxx7FfrwzxBeQT16e02hgmacpaoszSA3cxtW2x3ar8JG19UlBrgDJLpnXxYmUgk17
CbPVSt4qu+9q8gbVL5FpeiEHTsBx0SRyqT570784+mc3B246Bo5QzcimBoTFmGbBD+lgny0Im5Fc
c770PfQSqdJ+5rXjMwhQj7tqbmG7PiVh0USoS+LPbWTjF8X+UWBLv/xUkJZJ6yYgEcPtI3/AO7k0
rhcYdiEI2NS1NJ47yOsjakAC+b+gIaehYZXvOWJMzqy5R35ud67mwMYODaob1/MjJEk9kxQF7bvZ
VZp6B43afAfhuRNtBySVF7q174LY7Pjz6bdjR2XqHRILdku4v1bj/Cg7IKoVnX6QqCMOeEXB1U1O
YLa1pKrtOYaUHUG1dUYPKP7+LRY4nMAkhHyRcvQ67wuD/07F+89TY1/rek83gdgEgkWDLkNcowRO
f+m6i+2qHnLRMrj8PlicBWr9gxFJprv1ixQ94wBjj5DeHFYmjeZP2wFv6MN/tDBSgY8mFEUvPP+7
5bj5N47JdDyhi+j/YFuspWHx1a7I31M//88Vq1yexHBRmZBYv+KaRBf2YSgggW5thbVkF+JcQvcv
VVwgdck2KfzhKIqh/iW+YeiwfimOwJpjHaSQtScav4LCYCbizJsZIhWmEZGYGpvtQ+alMohzXsci
TDO269F+TACOEEwjUyd6U1H9Rqg0x5J7u7bOUnL+SthGZxfZADtRIuJuU6p+ThUvupxBBUVbsnF5
vJV56meuI3+AKk9xb3XGKAT+Apy0cBy/YLo7vtjmSY+3n5aUUrku/g371K1FKNWt9kiI972O1Hj7
zVdhU4vmr444y8+VJGd/lZEsrdLLw+mtDPMci0UMKVCfGLYcPwVRvfpAJibv0vHfVTOSlPRPrDcO
d7WjYg2dyeXtczVfgo1Z4wDMeKY/PI8kChqDbT7asfVntBmv2zOPq7rougYatdfHX7qqF+lRR83q
p5C5wUclVxMUkiXXUGmGB+O0bU0IroFnoycAg+bELnBfxMzquJ42BK/U/yeH0K5p0+dUhIlv1hk0
3238lk593GP7IhdJd39tyjAWAgNJrGr7r7Cdf7v5yLBcA9R0I4THZpa9NI4FM0HDGWMh04HhFFXC
wBEMDDZfiLAmOcwzrLmx9iyVaWzBKI32Ya1oEb7i6wJOVqfoWPXGAdzv2DoFJ/1nwM40p7KVPh3R
wIYiMI8w8FVzW4/8aCH3sQhFrmFIj1ovKuk24/6U0yRYvBU+dGvc61dt2acqrcbODL6c2UBKfBPh
gPBUnpV4BzcRxG+J0KfOhJTkya8jrm0Qu1z2xhvL4bHIZ/n9JF5qcO3s6U9bmyygnCJbchr0UH83
C7oQjnHZ18Pupq+ZNnZPmGMPLP4r9o5xYGyRru4wJQPT9QKH+ATmPGfLpKa+eabduajqo0GEN9gb
kCdUgLG+D7+qqAy82wSezSNUvJZlp9bhrlzZf0/8oZS+4bE1EpwhZ3sIaA7Z6Q60udHL1UihW/r2
leC+OmZeR5AEXFMllZqzrn4EZDtff5ynctuSq7tDrbIRsTh7c5OToJQV0qLTscUvSbs3VxzZ6X2l
99ULDCG5OIK758+++QWtS3RbMVBw8nksKyqf58NmfB2ZZ8zxiJ8hoVy1+tq38WHsYr5u4O6W/ZtF
jeX21yvDoGkecRzMXgxW0DrfPvNYA4d8U+cyNovy0TSxM3IBb7h7djSVvaAZb0UzFsBhGPmjueZt
jimxN2/JS+6bZQOMfq27L3CveEfJ/4Q6FE0ll3AKZuwM6qJVpPpFwtmZ9xFtf/t2KbHr6NMqozhm
8Wp3En2s6SInFIiIupDcof3Nnf8P2ewfvar1O6Zs9iUOR77aV3aPJOd+uLl80vO/k51MGWGBA8tf
Kz4v3rWT0t+z6e4HGkkNcuQl0HdXhABBjNjoDBTnGrJHjL9BGhlBS/oQI9coSH32CD9Yzq/FhCw5
GQl4AEtdyytVFghm5o2tXnHOWIWR6XrNN9Mg2Ba6xPcv0rKaWR5ln1T3KD3ltRnuyBE5ixf+ycP2
MFL76L0+n9z0yKoB6DjprpxmU3ac3VpGCUB5G+6lB6+UD+H7c0jVuL7YI/IyfMVdSZ35s5YD6riY
QGyBY1WtG5uwxGpgZwr94D15Ij9MM6XIzCRZv8l1Ym7xgcnGhppYh0aYI5DieWcils3bXc5ko2jL
wW+IZBJpf+5yKcLBYkOG7N4qTqUSTEkz6ZHIpsxEROh2yjYyC8SF2Ezg0wND0W7umLW2a/ehQa1A
KaJI8pRC9QBQECYXiQAL+wUwQY7IQwi2V9mHQUR5mxg5VWP5p7SoLPKgiONED8EnUOCJ2rtiNBVW
jF3gDWZn3m18OU8fZK7tBFbfOgUQmQacFT8KjpVKr22vLxgO+957d8iPybk5wY2xwxrN4cvZ6/mI
Ty3J6zEu3PFRKF8QAUXMFNUfaRRrVP63BAe4whRs0ARfPNwDWPrkX+ogbPtaIM+u7u1VZ0qzqePW
/I2pHu3Bqjl7RpGeawOBeYFj34tWadCobwcSerAKWc6Ilm8zZu0Jr2xgdLCRqdf+fhZW9+REdiwX
YXrGvxWkjToQ/ci1D2LilKfPBq8WLyBW3AUdFvxWtNMrBZkPpCcyNtN3pobSQ2kUGWHKIYFU5f8G
dbTuHmeFE4voIOBfs8YQwAlksqN9oZuJsaSzj9Cn6lHo9OzBJSv/56klhBtiBAyvWUg8O5hYs1LY
3/0uDRsIP31QsTJ0em8lG3ov+qcASAUv9Xa94oBSXzMz/71G9iC5nTyejkBCGOADdTTiym66gnrh
rBSYCBrgaofacKHaOMrq/V3JAHXOOo8FVNaCDQ385xrLOdJdus2wkFoMSSyY9TkSZe9r7NOu21eM
WC/Bcq6oBq0MYDweMzlKkcbBohMzLt/i0pDPLzkHqxgW/mqMcTsBCusK5XgjK98S90f+74AIXKCP
ARPdXx7QLTuLYhzCC2nDtWbiEZAK/VO9iRIOLfNKQEGjEfL7IyJmh6kmBB8MsXPZ3/2tY9VSMSPo
R6z72uF54KvHpYPOfdkaPpTZyIpGQ7nEd0238Eg6gmV5AWXZZUX1sqIUhskyJoNkvz9CdUXcSwFJ
FB/3YNTmTjLUwfiQ7R+hFdDab8BDDbaE1KbhNSlqZaViLJExVXeRIRRsDC0KmjHsfh1kqtdEEqZM
rSW/Y5YHrtV8RHVPMqJfDCriA7tCjrKokjzKDBJmik8DO5sojKhlaSxX7Zt2Q0Chf5Y0mBAUY3qm
/26Xgf4DUaVU/WeUMmWrHqwV+OAtFQd/l4uoKK3p5vxSdXb3D5/awb0+7qXnm0g+L77PYe0f5GJf
xdeI8IXPa36b5aaggugl4spZ2zMFoBg7mjCnulMIhOLyhNcSZwzPzlsymbVBDjABl8Ogsxc/6D0i
aGWycgnkiTs0dCcwN/fHGEf8BqHzmtgun9A/1zw5Ah9dI6+XVhGNO80gnsXD6UdEjHt+6Eb/EkMU
fUDWxQS/uHTkkQUPpyBL85YN9FzBXF0Rf8sjsjTSeLWOQoMOhQmk9UsiA3skI+uDKPbDUFu230lg
PdNdIT7Wkzo9n8Kv0SMlRRleDRp5gGsElNm8CI1FxuV84LnJicW7d2AH4GvoXct4kCkiD9QhpU0C
UYNRVQ5lGNSAX5kynVQQ5M55e5fvUTYfGrMI1hPu9yol5WgQfjK3JLxn35uV2DONEzejU9Yfr2Xe
egPDmgtkbNP8lRWJMIe7pMzUfLkbAHlJWI2OF4iAgpENCStGResAfz3vGe9e4R2C4hkU0t8qAPJ/
V5Fx/cZ+FXptM1DkrwJ1RKkICKh9hSfHS/0J9UjNWUwqhcs3ZfdP6s/K5pKfCj6/hyzr2kulZaMx
jbHzUBZRQczWRjQZwoyuKmWNB9d1MLIRt/7egZh4EuHifuiG6Bl7njIvH1DFYbDVAWrAXLYFbjUQ
MIhynju1O22l2u6Qo6R4J+1a7BdPnNX8FbYsVg+Pygqm5qYTyqq5OJnzg9PDHnWrEIwMCUfRDxGH
w2praujXFuDggMlSdTzQQx0KE5qSQ9a9aBuTNnjbmSXWTFzBUJmp0gldn7XSSbnH+KbIvWNAKL0r
HNLw3nsRJFapElQDc2wBfWgd/zJtAcNbQXwpF10qedQ0VqvMqbCtVUXgOvUjqWaty+MUum744fmO
MEHadWCavYOoG0jfo/KmLj7M13o1oC0DLZr82//K77NEPeSMPXwhaGjIm23m1bQvknfp212LbMwo
TYJ6F7Ez7QMl6/KA/e5FLxQ9mARZ7sucsqy1jolIhBXEZvVVXqF0BPNGlFGcOgU3W4cbFiqBNFfw
6iI9uwvdn9SXkxqZFYe1QRv4COQPOIkHXzIIVbS2gSr3QFsThHOAzz5MXfu0i2AksH8VekU5+81I
WmEo5i6esrs5dn4B0+93seJUT0x8rC9uq3ZiFT4Ej8BIWK9MLnkfaCJLmOwBR+HbJ3HtQEI15spX
X6oOZSc89BUQN+YmH+rgJqngs1NkXJc8o1Ws2vHghqRYYAL/1LGcIXmIWe56KJb0PWeI/evV9luA
+GS6ue1qSybIjVzqJwNN2Df5uHvsA2cp+cCWbTKayq2Qu3/kzsyCfyY12BpsGPsF4/xCM1zmBeIw
Z0Nv2Zx+1Og9tBKtt3l+p8/ZwqgI+o0CK35BKSRF3hIP80snzAKfYw1lNwgiUGEpwF94nsYkYCS0
ccrHYL0HoYb6UvEBdfTJMWUpNhGVV1AqEE05pBtXPkVEH8mHYu0UWuLDrMoIZjbhZl8T+MiNQuht
qWEZT4czVusmx9VZOO4ZX/1bKhtq+uK8RPO2qW2RLSlCxA9ei0h1I4K5A2X9HkbTMsmpvtegSCAS
cL4UX1M7pprVKBhumcNc5fGAZZXDEZGS2zJKWtJsbLEDfXCO5zhvkW4bE7fOBK2J2w8dEMFUXVCw
tcVp4KFUcAzJnpCD13kbNgLxwKQZotaA1zLKmVuvee2235qOTH6d7tSsuP9ZPrYwS85fjhXVwAEY
0nizRkbFOyy/vMirw0/mutBrFLMbkF1UiWlDGC0s6IwI1RTmz4GIEcBjpRHjMCWxyZb9gYtKMs1O
OS5QR1A62REkxx6zzAr7BKkBGI8guGa+sn/9hPxl0PT320BZHUHIrMADZL5/otsG/4purHejZoE4
XWnJzharav7pLvZzyqQAztQIWIH1KhO19QZ3OXwxoqjzF43+/1z5bdV5TF6/iBlcqJLpe4CogeUp
KmTsK9C6AlNYueIfQsE+Ec6cPoONPfYgRywzK/ZbSq1NVcr2LZqcCv6XaORixV58OsWltESkGCNw
rCJuqTO1d1bSorDWNpIPrtc+WJlAQlYdws35PRpGmJ9q5KOyV5l6K3pCkrMm7znBXcLCIxuirLR1
Axc06lz3lvVZTb5pSHRIptrrj854WDJGyouRnCSNnH1RdsqT2YdUx1QZqRdWi6cgZrimnTQigHXC
UDWJ+8roLqbZ9DyWf5gonGWexsSMtrdXtFmBN43UI1sDVDrwPvGue031wX0US/VduLf6DhBFfuqS
1J/1ELqm+EYj0xKkvbxvcHtmQfPiSjsovQ2TNZLqJCMJcWLyhtT23EoDpJA3nixlQdk1ruSIwuU1
WHZ7slXr5dO+oYVZmpiJS8qcE28V4DMsdN3oFmSUVrnuA1D5J+vBbqMSdYxBxt+Qnju42yrfPzbf
L8xMLr3ftm7Yis/kF84WGqy9XZtbRFZjAPpczDpZG9wKHB5Pi+DMIkX6a9abycyAhGzAfWicGJl1
VqbTaxVDfrMSgvrvMsvp43APheGPr/A51BEqQ5APmR2AErEK0MJ6/36OdJTUVQFDkvxXPZt6fWR6
k1rUA5f9p8hzBIS+JRDZ4qxIjNp1QXoo/LjxlZKUodQaejedGf9/BYmLZp15ujtFMKp+EGretNn6
vKoesvZ6LkzrBMwkaB6PTdv8DpvajsOrmUqYvRWWYNoC+SOXE2fCREbHFPpYOETfZ2GqjFF/RA2p
Rf07cvnMLpU9fOvr2Y6sYySYk0breU5vrgdSPsXKj0WXVm3B6n5w/ZLylo8gzJqFDe7dLN762DEy
CDLic+V7vU/rYxTGAQ81dswB/zSKAVFYjpPQXAlx3e7allKDIKx54zKsBgHClP5MnSc1o3VwmGuD
y0oevvbsr4swMNW0hdhxc4qj1xns6z6z+e+MTS9CapAy0QSpRfAhQCboa/StKH4DQm6t/gfLv0tt
WN9U1EXsoU3I3df7Tg42rf5wHLiCUhWeExFCRLqKelNNq5wr+45mU9s/7NJPo7YRaxZvDIOuMnJN
4kE/QNiw6C1p5LCyF6y+Ypa0L/FKdQOdTj6cIgKFqChmJaQG7B4HoT7An8jTH7U6h7F9FgGerZbh
b652g8ZwqDcs04t/6NJ5kb5HLBfEPM9eJHKnuPaJi+GkxIvaw77+IrSctbaJTEZGDIG9/sCjS9ui
z8m5NRfgJHpVSl+BtUwUGvhnBPr5DrtB88EsNaRTXi3y3g0cKJ1PLL5bMunP0r1xOscGFhjsAfKv
8oz2mqwGQ1+0AVznKwGYAuCyGaLpe+rd/74PHXXWir6tB9up2vZUh4y4Xzr9Se/tpBYTzZ+WH3fQ
xK/7J4YsR63Yp38sCGD77r3QpblfUspW7jfNpDI0SM1AYl6xVWKYQPgT90kI1L2KrwLY4JOtnsCY
ZHAaqJb/3fpc+D5aNXNSbl2DAqmQjb3rtpuxv0twsDFdcsYG8ocROuErJiE572ldwCtI7XVi2IMY
9EwGpzJ3+BWIEk4S/x73IGyE7+D9csmSx3fW3YzT0+cc9Z+8qiBnBT4EMOJtvwYlZvmdd3C67Kau
SpNiWKbgfaLMfxKrr3DdYxDLN6M9fj0KFCljskTxu1q5XmmE4Sy784m5XW98KiWgobNleH3zWrLc
/cTC6gOuG7ixLHkLiDsug09Q7rLMIdRcnDakzT6T7hNb8zzh6Fm6gXjAmTKD0bHRHmH2BhDsDwkd
zTDd95HxEt5R44ftu4pphphqv89ta6UumHxG0dODexdZL3kIXRsL2ALY/fCOKuWAfQqdtc3nLnbW
65umudyY1Y6qCbEG0BDGKlwQJ2ILyVVpBe5hlCMGc9/9zW/ufBTaIzWbT050NO2JKU9SUL/pbpNs
tuCyLyKQqo25xNifCcMdLdGh8DRaIECSpkAtZU4vsyfgY4+bWOEl4dQcPaTM7D8fHK9roVzcVULE
JeTW6lqsajS3aO5M6OUQ0BKS+SiDfwuux6U4JnLVP2MGeTn7T/7V/Z4mY/31O48h3GkCEdJ2yh+0
niV6NWhXG3dLJU4qzBq/d7O78fNCI+jeDmnOjzjI4FtKpO2uLg8Xjo82hFAxn7EaiPXdCTT+3BC4
KZ+WhV9BLE+ajhEaT5hel+T6fLcFbJ4Ug6VrRCl4+q9w7/HCQ1zyipZEJMWoppfamsmXZpsImn6h
Tfi6ARnt0tREyJdl1RCK5thiIG+qireKcZmVNQFuqrUvnQZ9SN2LhBX4Y6huSG1TN1Q0KmZ6MjMA
/TxU35HbFJuwaxZBSJwtHPGxAiBfCooH22gmpjBNLsh/d98d4voS7dx4kTGM1k2VHthIuT+J10HA
uaeWwWeDI6uxNj7p/rpxtpPG5wcA97QXXbu+hrihiEHlUW5jtV3B798/oP6VjcldyxGrrgyXEVZ5
Go5ZEmQyzvLt7omVfMvs8zc/SXWbEDNcSQRS32o9DhLNGNcj1ZDZ7wFi++DOlQjhg0yNZ3EUBoBG
SHB/p1vTt1NY/aGO//NIZMUjILCKjwxBpLQJbuTX4TNZaLicq7sTyhSPx4AViODmo4UFoOezZ7lB
m4Xv8aIa4rqSRgxq60WV53W27wRi0vjk7pY+p868Lnu+U8XSvqhYA6oSOd3CAmVff4l/3KGAIK2K
51sBrBnSPgqGsHW1ABmCZTyLA+Xlg2goKW/rMe/g7gLxF7gV0ITl8A96xza/vJtSSu6pqmikSVvs
uXPELZN8qEMuXs6MKfRfoeLr7WnrPDNZcvWDujAaqQtvFvwM7HKYiiupIrryLgElZ/CNjEIwVd6R
1UB1Dh8yzAoOgQbogFPJVn+wxMcHXNO1OREs0ZaqIy4sLEJHkeSAY684j2HbOdEas3eb+cgUmNQl
Nr8gD9M+DHmOdHUMt9PxFdzMUxQsVan51MUdwTiKcg5GJ/4S0ufCtTcGOlcPSyehiLyTzVMdJYNl
+i4r+UXUy4jWpYXAmV1qoWVgN9FAkZJtuo4tBHeuGBxQYKvGKXjlLWCFSK2pM1mdIuULqt0Mg95l
es69Y8XjrNH7DkSqVTFvPFiq+X7EUZq//TakVCVBJDjmJG9ucne+FnArtYkcToBi71GsgIQtZDRO
fKUUTNdJZBNO32nJFLQ2RzYKlPuxqxmxg60w54kpJ6Og6JPYxsArRIrQEG0vkwOz2fHxQI6TKyGM
F0SJzfUHmGvAEKQ51gSwQZm4HDUF1vSIl63M/qv97EG7D72pXgGvdipKajYe4EIT8GEJVzZLNUuA
hruCV1tIwkJDua5FZfaAGK3nJVFjTf6RGL52Jw46tTrAue4rMwSS193whC9Oz7UvFNt+CbKiCeTE
kcRZ3tLD8BaHFVlMTIzCsYEUpNEXF/mJc1jMYeHhBnL/5QEt1mh/d3YaDt4MFufqVCLiOZRjLNkV
0lMOEHuoS7/OzV944ZNVbBSkRlyp9idsFkMPz7X3SIZ0RQ8X8ziov0ThB3SPdyKViOF6RnVuBPPM
8JAFx/d+1zOqR5C19CEm3y9BMLECe1a838rO3440+Fe426E7jctLd2PtLrtQgXhgWZzzRSPfdhSS
CcEjEqjRUiWrwJIqxn+94wXKkKw+uUYR3weDYbsE5k8KuqLinW/VArUM0KAFmFo0zlX/YbehKpru
s034oPz02kEecW1pwjrD7xUqxnv/vu+l/TMtRbhS3YuXUOwK95QSb4SujX8A82CG4Ba8NYEC2Jh7
bHaTWI9mZGMdYgWcvzeBNGqlnwLvTO59SxQtXEu1C9sQgHbgb7Xh11DQ/qHTbBXkMsp464zP+ve4
uLsoElw7lJomQLsqBMpenwnHAjN3z1ruWVjx1Fab1Obftko/u/OSS83CoIOo9l0uVyht9OD5cDiC
+HKxvOkdyxcSQoB3VHooRoc7WcoBGkatYshSeR882YZENen0F89+RYqvtt8rHF6gyrmu2SAkrtNN
BQ2csiACOIFDNd4z3Nah91CF/9n24bM5snR1LGWewImcBFc78JIFYVJopLZkdn1xgEWhNDp/ohFA
IkTHQj5nyxy6UzL5/18Av2a1axnrlLfO0orYWCu4okeg5xLB7avjezZUCfZZp4bXpbCxCGKoFoyb
Gj6fmois6kAhEPbI01J1ntCqhrkNQezsR60ULQDFuszpqr4ZMjV266ARatYrc5utMcndYB4j4FfP
Sz3nYSKFE8G+IYalVvj0SF45lPLfsHZOxPjtz8de3bieW/V0yVwO+JO2JpCGahkjipN0Zg/sQfGW
N35diRLFSo2yo/b320R10nopEK+zt9jEzcqk2gy9AUlHepsdoyXGskPNXZ7xcI0qckmjZQpsJC6r
5oZpFXxZ34zNeJZyUC582nIiurBbJ8kapK8Wkp4nYfZdI0iya/1mmvXlPVcr2s4EUW3O1KbbPN4x
+0XVk+21dUajAH59Tj9y/Bws7PyZEh37QaElLgACB/Tdu3xi21UGK2BekNcVAjFajacHNPEjTviK
5mVEgCXOyLdcKnZJMpIVf7TjQ4e1LOhC39ha1JF8j8XpyGYekNNSme18DGP4pX+5R3QfZWaTAx6Z
mHcxMlRRWaFBHqP1+TD4ju4FERDVIv6tbl/ziAFbq+s4m/Pd4POFYo0TI4/zbwTLBi4fxDx5Zt12
M2WAJnlf9qG45xTljoJ0dFZXjOrBrWDe906i19m5ETXphN7jwCsERa0X7JYOL/l2ONwnMMkwYrH7
urvfN1h5b3CLcP4btZLdCKS3nuopCZgVFWF1xQnPpxTdsNb3ufy2DEP/8Isw0GUUjkDOrlehraDw
mqjyj1qdCSZfoV+BTh+x8qntShTpk8rDXub1/1FteT7H9KcRRaTapt2ayEiqgB67FsTzKJNTz9ny
MSKdSKUPGvA2mrqZsTE8s65H0Yji/Sz/zyoV/iTnNnim9p6GDKCr4Wi2FOcprSTc7Epa0TGMMJwT
vBZNCpchKj1HHiBvflTDidXwNz69hyJ9IokE8XEbeKttLQ2MDfiXXcIJKexDyP59W08YihEalf0n
0+oJxMA9Xy9/6pd7huM4RJCJxj7jWS0pqu0FT7hHPDrZLh8DSk5iNOaQsj6RdwsFAklYytEVk73J
sK+NJYiqOHlsZ5ON40l8MVcPqHF1pxMtIaoXhvYNSEX78d8hpkRy9fpjKqwklGTEmghXu5slysw0
s/7P/QyT+7QubgNfgVMTlCN2N4S0/U6Z4f0aoIStLy5sOXFEU/wS/wU3jt4asff5uxzYpL7XTT08
7N07JVY9sQXyPsUlYHBn8fCijQ1WRbE8QP8qO7YZb1UEl/nLlGeuq9VpUymSQsEf6d/KzBol/DhS
X7YC03hBhtz2dpJLDmxIoufNoq0nPVNFRLURiLGquQJNERB5toe2fOVTN58ojAAuLknElfRjFPre
AvoMq4UYx8UZ5gysHsnStb3QbKlOnysJCX629O2CVrxSnUArFvAz4LRFZUT4wEYguzbwZAZB97I2
mHWck/GhWFFg20SDperXbHOfHaj7fV2DlsSCro1fradqcjidijHX66MbRN22Py3ka6XlWB8gY5+K
jCTkadC91JQ3jvcheM0ZRGVzHV/ryhCMn6PQsYKdMcq0kkOd7KKQwCWN9gxqBVADYBy4gEv1MyD4
ikU1eI1mdxt45DzAz0rRqSM88gzQqRSiIbhcxXBMno6ZumshwqHlmdIjmh0lJNY5dI/ASq9y0RS+
p356IbcKaTYEQmtCN5+mMYSPy5Ti7j2UyRu6OLgd0NN8QWqnF7PtsCx6LqqJ/vU1ahHBg4XcvxEn
+xnbvxRbJdrHzbf3YBvr/t+Q8nGaR2MTIP5yMaLuNveUM1nDx9c7EnvGp7fdFubMJjQM4Yb3+Nxt
97fdWC9SHjG+SKk5nN8tEbMTv6mFMFsYwzh5mXU3M3kWKozzL6K+iUZh79LvJptLpu81Gfi+ysp/
FdPO9Lo2VjDNxwTkGLphQsrxNS/m6VS4kPuEpKGi7+UzzBXTziiF41B0xsOll6ldezWssRor1loB
lAvUKKhmpFINFmtDu49hGQloErUP+6bNC+1Zvs4iSaSyIQwHWuOmYc10HZqxxvOlmCj0ZA/heMKQ
yYHdQeRnkbnntUwO/a+9S3V3LMGbjI7lXw7TDmIgljd4CN7Mhr6S8Pl3kvMupfnYN4nGTJ8+aym0
6BLIt6yYzdlEivgcYJN9yQZTw9yqiyDzu/XxR6/p4B/EdcrNgMq23S4ZLUpzq0jZj5cFJpPZmMqo
/iLntrgFiW2rbgFz45fGg1t1AjJCSRiIAbkAb0IFlTArKx9M8ilVIKuX2XMMYITngLp+nqvMGWFn
OLI3vGACjsJQzDAaF8LXe3KAAcjEXdu+AuAbtDAJQdzS9nQXMm0/wa3kvTH8lZ3rIIaGzkgMF/qx
NqhjZH2zaIh3IY1Nu8oIysVtP8hnL6GjiMnzqxlfMs2OFJ9ddJb+1YxplFR8ApXrxabRlcfp3x6y
nBC40DVTdezmtOdy8nSKuWv6TZKFTcFhhwmRej3dBU9oeAS+y6+QoJg+mcf92qDIoHqD2NTPtZaD
7rZkLfyyZv1S+R0K7Ld3wC+FXdaOnnmbRC6b1GMasXX19N+yIBkCuG3xT7OhoPIdindtEI5pUq7a
6Wj0I7BEDe2J6HJ83WvsCR7RcoDruzj2/hCF1Agj6F6+nZhUGsdzM4654kB+Olx19ex2kNniYDOZ
OZ4J4QnGegnqFdTYjSuPbWFrJnR0k1v0ux5/iYTCtcZgmOIXar1rRQv8lNb++XpYhbdVheH3+ta6
WfkAB0r8qy0Yw3nVsoz80Ex4MYv4qBqgBKBXPfBGC3niC2Z6WW4pU7JK+VR7ufeYkyzLguyJFcfO
ixGmLFlhiLoL+RLc35oFp/oLQ4ikdSiCU18WljyyeI3msFxsvX9uEId9m2SrKuUlGdoZWnqshLtE
VV9qe3gQoSQJVuKsZbvwlJbWE4Q7a/3oylKXEQLyJP8K6yS4Eus0VOL3WL6BKh2OY3lOPeK4P3cI
u90QbN0COa8PeJ8NZUSeXbVG8dndzTeRGjSOwqcnTbXuyPj3GOt5Ya1mnV9Mk1ZTiPXVe9sGYjlQ
BvFpOEEEuXCZleIW2tuwEmfYHbAgvu3Bc+Q6oQpUSSnsdS43f+Kepg1Zg419UhdTkT8vfulwEs/m
etxveALWGt0tdyowzX0WGqFL6VzW3iGEYVCCblrYsGQhzZ+OfWSN5wWyGIzOvkZ7OHFm6QCnHSXL
MIuTHMYNfvgyklvennXqGYdHO/XKLSsHJfj44MD1U0YNDqBLI6LuEO3xnkDhMMG5nu8u+GTjVKdU
4wZwXMuP1b/QplflC10kSbCRCpnlz8WsIx0Ejqvx9YjvTrQRxbwKdCs4DmtAm//X2DzHoqiZktfd
Kto0+OaREs2qw3fVBw51SubcGcZO35mE6/poEeJtF/odw3GiUaXA6a58XcVktH6zFJK2v4zZctWo
ke7WPuxAZ98arYZkGXF0jL7x3Xlb+F/75lVmfT5RxOehMjfzao3WfTNysrDxyO/21jg6ZLor7C+2
nAs7hmOSsb5qYgnnlay/5ctVTb5UDJtoP+T80WvPCas11CeI3K4jVnVsp9vZRdX3sIhE93fBLvls
yE34cB72lafK3N+aukikeJg4kdkJkuVkwpgeXpJ4+f8ftZ3VKCronQ3Pmbo8BKnmBNxrofHTNUff
3UHSbVIV480PbDBJiFpMRHWrwQRmPXinzbQAiUJ5We4RlL+gJuQhySPyIRCrtFLZbQ+7Szekk/9b
WyrFoBQN96Y6TPlqcSo6/xcKXaXMjz/5u4ssPSGXHNmhVGihiakj10WejqBPllwhrvYJ0zp2ZjH/
ajugexji4H3QMTRvHl6jnq6kkfI4fNw/ia57QC6we8gIQ4d9IKoZIOYCEvaN5VX+I7lDEApOTRXD
ps/0SeWKzTPsUA08oOUNJNA48TUQQEGgX4OaXKVbNWSpAd+QnhRIsvQQjKQs7Y5++wYNCpE//J/f
r7hDhOFOgvCkc6ut6bfrHaszzoqm3POcJ/2AR5P1CUqOiEvQMJQAwXGyjSJAkU0iSCcse9dt3XcZ
mC9KQxtbE4awzSO+j7dnjA6IdnOjxxGpLfanjzO9WVXr1S4eDamuUu4rUFZD9LVCcx35mU8Y1g2c
/w2ITrrfF4NOE44RAYILALR+qsi+8rcuNmQfpUfu4z9T5BHQmCG/3lT8g658kDOVj/s7AyyJ+JE3
vLx14hT5IsRg074Oqawpe/Vl0YSga8yGDCZ5YBU6jXsJiaTpjf0FmOxQWoV9rLAWRKuWF99dH7i+
x8yGNBzDUMEpn+lJQUjBCJ5AaZhTDhAGSw7b0MNLulsrgaG9/zhR5NkBFFaEo9t2aLv5q/FYC2av
HdFt7XCFEci0wkeBAGkE9bD74EXibzcA5WckeSa8e6UF+2H2ijgq6i6tvNYGbEfEDsO+kq/y+CSE
RNhX2WcxJYH4tFyZA6sbcosOp2ByWb69rvW0jo6XzznzOMclXyRtjoliRj+9k8bTbwNxYbjusGpC
seq9FXzJipmKWKr4+uBZW6p+N2bsdIiUPC/DitzEUwxZMWGBqTv5Wr2Vn6cnDaqFvusmG0N4mP/B
BGFQ1KU9zUpvRacxvmitK2g1nI8T8RWGu6808lGRa2950SBJM+tMJWqIQm7R0g9XynhwlqcMDS1r
MV1K62pGG8uXOXOzq1uKy4UkTmbydFEojU3Kw04usXD9Ht7fMYp76UJNUzy4foIoDqfvsYJ2Zvoq
pqWTLuOzXv3HHduBJ8jmLVi1yGkoj+ENZQ0/w+nM24miGkxeyY4GsihKXCRdBd/+NUlfW3VXw+Nk
VCu2ALsTyEa1Ptik5N1nxG7IZI1XHeYfCqyLKYT6bKEDYF+8Q5FuQ1pYbNn5qFyOxz+gtNoAWJzU
7N/A9KvY2yL+8elrHKzC4UXzk/nJGLZW/GKSbFhu2vdxqW0hXAUPyWS4BTT08eoJAD42DXN4UPo0
KYCdsS9EYXOxQyfxmRg6YVAM6Z3j41Et9L2xSJnzgT2uy1vnOW7Dj7Xvv9xWQa+UZiW4zUQlcY3b
hW6a5LFSmfvg5pHRj/9o7v2kPNPV6znFC6lytV+T9EjqtpAoLqkbRkC2ZieuVbrMPaO0UDQYIxdm
fq08qV6npcjHs+t5Af+jJZLU4dkBZfI/k9D7PW1AgoUutvfhe1ZWoYc/wS6I9+X0bNNP3pDhzfT6
itSP1iZuzO27dOGpqJd1N8AZpfH4j8ssDTx3rT3oh+GBb98NF/TM6nAQYZy7IetdYVAudKsfdMt1
SVHwrrOxYxnMgUWvdurCv/pUHUfGPIMeyhP8X51hnMCYsA+i1uuo/RdfT22/h6Rt5JmgpMr/p2S6
m7WMsW6q9D91VenNmTqHAKDr1d8PCBzbmo1mFYrCMf0Z/zlNagcNSNOtL+9jZjQZEDstZpQdffKv
nmLNoIBiQIn9DAYtGAW8c1o/ILBVd8nu9nraw68bBb7KTtWGvHG0kqplZyuNGSFmzZDwnm73v9sM
6kwSOtCVYSsEalVgzb3lOaEuqU3gsVq5devYXGBbLm1HgxZwSIJo+0BYzZakr3ymyJfgHIeYalcZ
iQF6aq/maI4ae/uLr1JwXx9eU+fF1X5/u280VICyw+1txchrDX973jFXBd1ZphysyLHpUe/tkTOO
AInvDONNSReF7ogd2oaS4b573riw8EOl4m4zp+7WyuMODRqtWmIveXS/yn/bVDh/ppcu2s0+xGgX
0OUDm86ZavRBHjaycBMmtkQtlgMJqIIP0sqzXNy8usUUR2S83/C7m7YA1I21eH4Fg1c1gxMyK8L1
1zldPhVj7apHrZ7YL75Qsf6xuiTfxBUIPfKQNgMk0Y1F7gXUfTWav/q6BTBL4ovOw5wQJBPY+Pxj
jz8RhDEFInRSphaxQbxpi3QuehERExXmFL2jnf1Q6BtHaXW707BnfHoCecoyCbHqEU67Agyk+CS0
gszy0uAMZHzfdbEB5k/GNW0DbIAgx2CF402HwYxDPMNOhJuvr/czD1HH45oiQVlMTarwQWrOkUQp
YuolbbZC8cKbCXssm1CDqSnq7V6bUFkK/PWbUud03DaRgsBtDXDqgY8XVcQkvyukvXpyvHJOod7k
BtWYj7GnADZ/Gsfbuq2yewJqvdbzyZ4KDTgTqFq8UExk9SG0jwCms5YkP5Ma9b3xWR9kNUThrMPE
7xWeeXlyi+qVVJOS6ZK2oA4zZ+bSSMga1yOC3gIK8niVhdchhYfBV+IL6E99XzSR2zVpmv1RzEpw
xrHEOTsPrxUEi2hrHl9sEWUmyQEZnVZLbgHnQFHAtKAJyCZGGr2SYvsCwguc733TbmEwrxMMmA/v
6Qm2DLSVbHtWPXBiPRszs1I45EdPKNhA8MgAlXKpuIy1UFgzQz+RibDpX7sU8GFoeDEbHzydDNV3
x28NDKm2yBD7w3e67BxGVFGRc7UPT5ZVs+m2LqdDinHg5Y/S8NADN/FF4CF8rsftiukMZQxx6gPZ
E8Bhb3vdop/NOO6sb7fvjIqCTjOJrNgR9wX10EeqfT6sNFCIcjHGTOjs13T2lCyqp58xYdqkwyam
usJ3BtpX4YjMkD7xSx6dN1tDB+IV6sTAVVHmNlq8w9IpfO/rz2D63SEjNg9+cvaDJf+QEm/vnuYo
nTEhk558QWgm8U4EPC6ZUhVrWItSCwsL1yjSx9DDeIH5ia4nu+KU04YXJEMD6sndGrs1SwxWJzC6
vccbitUzMAB2BRpSNn7WftkjVUGekO/1YsI9pOj32YetYLpXExUnVeIT3QVeYLKhCQ9586jOE6rh
o22Cnz6U0Hlxa2XF8LuLoOoV9KQ3zQ9LUZMUz88Rf5iR8NM3JMT1t9MhOPIJxGd8jMsPlcSPbYwY
8dblIZ943pvl8cYWYuZmfxZVNNVTGeabBzZOVSRy3C7bTLI2EBkcw7wI6Ccgh0K5grBY6eAGYRny
xoYIGFmEi9YWDnQWYAHlPJj4st9tWyqXa+ARxsm1MXgC/hRlry5qDCh9s8rtV0Ih09+PO3RdItEn
sq1YUfv+bFBuhKu+e2vyXbjFhj4I+xKHlRXHgoi8GkueCoAkdgtmvS2OdYu2hsF93NLR12zUoZKc
/f6hhJ33tRe9gZkhNBkMfPgsT+SnSZaA6Zm9ahskxGTl1qRefrc1rnMT/giv+QK9tAQM7QCPaxTs
NmHAZrMsgJxPlCawYDcJiSU0AQNqzFfseVj8IfN+om2KBH45tIQM8eprla0t3lHTNnDXSln7v1Bw
IvaAjw9oQIXhYwwYy1OLIoSLTENhg99Xjk4mUrsZr4ic52BoHOH0mwxIW3Tk74bwkttiv4YWN/NU
7LPOShP4nDoarLiVOPi4FmHEqoqkzuY+MK8iUdjr+6mSdUnphsrt8gLfoLpEi238cI1cLU2IVRcp
yxT2paf2V6UEREcNMQCXhvXfpVhG960jkfyVhkuD8dWecyy95lU4ZA7f273peeEQJCERhEudfLY1
ZNlt6e51HF1z/Mzn7VvEZavmckr/8EWcPWgyGRpaLSC1whahRTy5KHMmsgMhxpzbIhz6y72ZaTL7
B0XlXgbji0uhou4Us8zLdA5MEPAvaJHmccfmQadqrolOyV/73AE9Qx/xn/vHDG05fiVm2RHOqLrR
pmsgoBJuRdIEVbJ/vQqj8cHM3X2JVXVpoY4d8sIyS3sK7nixV3DU6mG/aJSBXrvFYra4r/npEc/b
8MVpwRchKq+Gp/W1TFv3LPiWnB7FrKnsG4hjZmdnPnusHY/BCYo3dACDcx/GNaGMBcX9lVKgPsnm
51u0BWvXibIvnmLXdmhaFVd8zPxkwv5jPXDKwDy4O/TjTDkDb0DGD8RTlaxHCinlpnDV2bbdJ2uK
Ae7yocsY2SdPYAqro/YQasTzyIQ+QhYIg66oJq0OcnMnMVveaCGLr+rqM+Ku8++8W3ShF1w849bb
UuEQQ5n6SyE/wu2vnMkK6uGf1cNIveM4zBqv5QlMLmbLcLbPuHQ6dLGk7qk68VtvSy9gIYlAOYHb
3ujuVnypwW20ouhveRTFXXCXnx5NNWok5BWX4bdjnM1VqwK7tIsDGw1IJgA3mnwrgY4yK4lY70z6
60F55D9n0CCBiSz+j+r2hjXqwzkzlMVCHnLrZrYzoSd5QNKbsuPGQS8cyPbfhKoNpatIajN7CBFG
xdNIXV062oW0heDaqez94BegTYO/FpbFCHH9+44nRPq+FbEcrvEhv/NDwj2Ql1nv66OC4mEw5n6o
UbvsAHm5CUhYEWjvtkjW49Vcbfxbxeqn7NIIHEZmVxNAgzeSKc/1WmY3Zt28FFndiqqrRBftHlM5
n3SR82KUdJ7WQJwV6uc5OnV6GrxcdX6Jw0s4QtJNWRRxi6rbU/2b3BmR889Bfy1VETvF+Nb7nWTt
CkMWfNvz0ieAFcC9EwrOvqv6xhKSo3zk9GuHw9UrYJdFDHhjZUoHYhk+/MuVN3CyzNp0Z6ztLxcp
tK0rYOAxzsj4DmWJ6OSsr2jEQcZSScHeJZwkRzpLIvjzmv+YIBkZ1bXfg+ayIWwJ3HJtBwh2XeuK
gHpVdNKbnNNlTYpiK/HWO/IdGL2BP35dZA5ETHRnzzdR6A3C2KSdct/60EGRdGcV7nlMYNnkziRv
ypG4jHoGRemH/vVPb5o4HH6Fdeo1BYREmxNV0fTPaRxOb2Jwkt/fjukmA8cdgJ9TX7mb4cz54ubK
I6OipzI2mrfdpxZ6sCdGAwV1koA0dxhjgzWNJQn2qPsiVHzHA1tLq/UEB9oqMryuenjRZRZx8lib
72PmzU7GeHsBAIvzV2gVfuQRX7ZC6WSGAqMKGb0YBve/5GbrlnmLgsgZ11dbto5bKzitG0KcxC6E
3uCTt9IEGMaL1p/T8XVIQtvrEIpcbes/FM0dJlYWzPPb5Df44YoX7O/muiHysiW16py/SyivPwpu
jWeoNrfOZeQGdfVUVCINWdMYJsoENbQEzK3wl9VA7IQznBF8wKqmYxZtBWYNtaolJWaHKmAZpDDI
ZdCpdyBsO0SAaLTujl09VN69zxguQi6l6XbS2jHSfVvdUKmOWeKUUU6lmC5QAkd1PogWntp/6gqu
899bYzNfILcmQ/A5Loqy8U9UYruDdF6MHEUE9pgKUBZ9m8D+LZHLUtBtlZPvTe/AXY8b212PlESF
PVrZAq7TfGPezvxbMLLxjcf8ZIn/EifsIgokAcQ65Ho3WCggWS51cWtwTCQZnZLr5MlMfJku5k1K
QC6Y1wNOw4wTaynJkMyqayTddK/D+0drWM6OcwYncflgwnjFsPfS2C+Cp3Nsy8RQBHLayP5BBNBH
3/r0Dy/2J7YB/62frNpcTF4CeMG7IV1SkUYag8nhnIuBXRefo8LKJg0Au2FShDLBTQW+tI66NOkk
QyhvdZyrvMiBuugfDH8LND5PW0wjcF11HuI0BoQGXcHQpkFn2Pq7NEIiKcuVa2sxnMV9OBG5N/75
ac1B9rmuio7iN8pNRiA8maR4smO2TwKGpTAxtyzWrZxnqpHEF0tX7GN53+njb3Lv84R/i3tYuwGk
JFTUFkXTJoM4uSRQstJ6BQiYOuLLEDP1lUij2N/d5Ir7QodhU4ot2WL/14KEGj6DoaFplTm9yGNO
kMmVxKdSLe1kUTF9/zfLHmHsel8+XXoVSorPDxDAo6zRRnWA0s+6Ow+KJqlHZ3Qu6t+33cKw+Ec0
1Q9kYqNHC492l0KiQMJjZbdWSsSAxncR/KEeIUcHVLMtHHHkEBdV9c4rmBwBdJ03KtRG37L67GhC
C0O+CMuWR7FGkwrGQQ/WXJvKdmNVqrFXXaw941NDt0uk+ugC5+Cjb9hfXv+YHXpaPYnUfLpIAoiL
ay2/oOJ5lcHAIj516QBvgdg4Cr8hZ5dGqZ0Tas6RlXPStFquZ6iF6cDzfpnjqv4eVg1tKSzmIThG
Uo6s3Gr0GMfKnpUV5fmvOtdkjxbT1ZRMhtn9XdLK+Ay13tZnJiEiJo9gECGYp50dzCPEpqnU4n3x
00Ugz3GB+3pFeGS+ubJymLUCvpa7RxHEM1XQZp+y2yGwXc3l93DPpRjEHSJVxYL3OGqPFRTHlQzc
1Mxiux4If66/m9dapk+JEIU08rwxIfTA8SDrH5Ji6Jg/mUTssN1lHv3KLnpFEqR/x3sn5YZwKW6T
iyRCxAVub50KJBFaddTu0Es4fT+SzAgeqslUZq4cxC9PtaEqAd5KNUIKXaLJ+9lsBFUuKY/GkSxU
S9nTqZFShBVwZfWxAg/1/OrONlIFuoJQQb6ihAJjqg0Rmqv1CsYqVM+IMvLej+rbNz04lFk9+WuN
QNw/15Dfa8CsiHfc9H9QZZALuvsk0+nhUMfunn96W1Uv6ED8mg8kpnCUs6ca4jsmcfNPS7IjmrB6
cGyaykk/iPspy5AIHJratHmu1YMP1FUwq6qbzBubnoAEsSYIaA9PZujX4QesKqOEU4wEH/ua8q5P
8qFn8BBHJneJZ3pg77zvenQCFLVC0pu0EL4HYr6q58nRtnNDo4/NEY+G6b3CVh0DJBgJurqKvUD+
w+v5Z9XstvXW14U4uprSXeR7E+ZYrwKMmYmjEHJiBZDs0d0hv9qwgdK0PhsnFGNkb7M5KGmBDxLn
de//UEPIXpWg0xmL4Gag58jt6LB+8aN76kqwMtcm54XoHWdzs138tCytRtg6p9V9teTdXuTUysol
dD4+x+Jh6r3W/v5Xbz3c7WWj157Y1GisqLMfe/3IN9fiZ/SYj4Jj7P/Wja8bagvpXlc0RRbTraKt
+y8qGFJC7W71R8+LmSowyMxStL0+42iDK9rd9dVD/PQddOFs+qpnbahP4QFhYhmfJjJoSMpqK5I2
zz44DgYr4ZPqVA9pDI8VPmQjqesmdVovCXi38RVdoGFGgJaCjHY3IjJHrXLpXZhBfpe+Au7pDfE4
hoayvQXpEa/+Lq0YFcwSZTEFynjO2pSVXvEX/ImIpv+Tp9XlYXEH4gc/Thji9/aAfd87G7NeuUZr
/EhziUwNx3ZwygmjYItGysLX+vFS95CSSWcdR0QFIxiCu1ZKO2M/pm2VG1hsR9yfrpSL8TITKxUD
EhRkFdrLtlhgm+ad7dOIpinoN3Yf7y2UZvy0LEi1gbNujdaiTMqKzARdelz7pxENAqEsKcDaVrOc
9cJUFeYoGjbeNpJ2XG1Fl36DC3w0M+0Rkw52EPsOWyFiPnJzBluCXTkdQALtSWuAXjGHVnUb712G
+ivh+ThecdSeyjE0O4iTjZJdhkTKZMavpjrzkOF6dyjBnNTbM69FaFl1sQqDz+S0c6cypwxo2PKl
A89bRiV5hIWmjHm5efHBAjvyForputPNfNEt0RMCA3uBYBh/k3kzrYC1Lou+bzNBg53/nH4q2hag
f3Hd1o4BZhw2D6FLzjGMlEFypIjW0BxHcavARSqokhkSGfPy2bnbtRCnAX9mA8oQhDXRf8f+OF8P
lY2SaYc/09eq318qVHeXFtGWi54rsVvcH1gNuGumC6oOxyhHXeLpD5U7srgI8GvnbflDy22JMLp0
14EubOuWTWblcO7nZy0jyBHKJBK+jTAEUoURR4nJC0R6n/H6SzcPYuvFlEhXKJ2ieuHuGJ+NLF5Q
LoCmaiG7lfLkT90/fju5vm0hSZ63HSFEy9YVXTDjjzmFu5g/LJf9RswHSjyrhBCkx4u1V+aMkeIW
hV5HE6XcmbTyF8i5Cy+gevYCSA2apL4IVPyUka6MXDWq13GnZITrl3aA9TtpE1MgZYAuaFPHOQyg
Mu/lYwDsTWd3cdE+h79ovwAkzNskGcNtL7HUJ4tRmUVOUnEl+FAq2fNRNXSCPusbYkOdK27Mm6Ra
kjVfGVszR/p6jUjLyyyLxZMn9eusveaYq8IuWJQ+MMVSZWY0RZXipMdnDb3/4CVUgsvRDKH+7Sq8
KDo1abn8u+dLgEUOmRaTNE7R6QzWtKdcOdViWu0xcaDHVEeBFkIft0mBA9+GZbSL5zPvA9EHmonL
RmGrwlCXRkjFUrxl5TIv1ikRiu5X5OoBLTEOegdP19PRb7svUUXiTImhi6bOQbJA1qydkGxGtg4N
l6J/ORWlzvZjGkpWHyS6ykTRfyMEEdELHjzsybsTtt0jSx9D2r2qsRltN0pt3sm4X+yyFcnR3qXI
lLw8F0BxZKD6/2rhv8/cAJ8DIa7ivMP4gOaHq0HnYsZE2F1lAlspzofo5YEubl55iHdbR3kQ2Tzp
cDX1g4cSR/58C+OUl+yQzWV0l/h4p6jZGs4wVI0eF1ISq0Y6YdZTkHrbD76qTvKHSlNroMdUuu5J
a/Mt/QiDktWz4al5B7TU7Ijan3K+lP1nfSPm8H9hu6kWoNWuZIKd6pcCN7K7aDWuJ0L4d2msIxoL
RYf1gNCE3HtEAEJ+TmdV8pBEld/QLabNjHzqT+CHNVZsTP4xvPoaST4Y6yeKmy23TonukD8zyEep
FwhmDt70MpuJQB7QPIxewWIbaEA76HZLo3pwmhaxyGqwai0BLxAjY1q8XsfEyujlIRBFeYW/s0uz
CfFlyFimAhkIyXN4s0AXR4Ue1lyy+EsSoGZ0M4ujcfKMHu551q+bStf/eT26trOBLDMtXCxcZQuU
wpECeGNp5FKJYaRzKIgo1Sccq6D2oAVXEVDiNxoAvs8YXMDZ5yekWjdS3azg4BQUagVi74XcurVr
h1tHr9VLzyOhB1EWhixAnqGtOIfTYIO7r/gWt8YvhXXmGn7jUxJHJ3T5ksUmo0nHZn5RDPlLfC4g
cv2ZdzCJ94A30MtF3eHoFhPJcRq6fCQ0hZDmiUqiWo82FjRgxQDtJLTk4Np6CqfHD0V1uujeAk88
VnSsPMtiLCiepz+DmDIgFNFwJBu5BNYc0aZhKUM1L09RcU9GwADLSxJwMLXcIOWxJOTnvBW3im8t
FWYSKy9DwcDOkOa9AZAdAJ5fs8OYuBmM14vF+yujKwfoENyqvrACfHwgYDz9qKqkrKC8Vne4zI+t
04x3xVFrZYTZyWEmclvpBKUFre/aLoBEStoyicH6+O/SaLnmFuBmENmV+tBWu3yjNN5C9Cj66VPf
qGZLEHwaoToftBOefsWGc8MfdVrWRYZuzRU+0wpryAg+OWtwABBeFaImq6dm/IRs4TftiD/r7fkt
wcfiq7v6ScZlaCVOSO9c+GcPPoEi2fiEq2DAZRbmXeYS6tEAbtN2bWnCPcpX8euQIQnhtKTABVkK
QDm0rnpmr9pAVnUPTo1kQo5QzLZavcURRsTKg3IoCVFOPocALIvc+QcAhcwHlLOpsQHAThsMrRFd
BZhYLzwEiNarPpdbkCodAPvkhCR9bRA2GuUszDighMKvNZDamBWUCMCiOr0SJAuePZBVxvtwjAyS
1fC7aE7O8Dh9aC842VecqjSMj2HyErIaYPtdufyXWwBXniGyXZPb85oDz4K3AsVZCqW/wPOtGmJo
ieMt4Fsg3FeqsJsZWDwwSI2YEVlHmuOc01cwqP5uBGZ8CdgYDmZHINAdO2wsWK0EhCtzvYh6MTrD
FKQRV6bA7bwPydb6s+ROfSKk2CvTVsZmwaYgOuIY7w70V0gZFWjKxgn1goe5N0EbCeuqIyX3frmt
TBJ0HLSsbr9ROkkdIt38nfoulXknKVAE4GObealHGfIhmYAHoySNCDqUufA1SkqhPnB++OqFVys6
OSv65JGzHVKbkrHoyavJia3O2rTkSHf/wGouTdDEap1amo9sl4NKgHr8AIGspaWMCGWrGaSxZtuQ
CajixbqS6JcA7v/7O5/6GaExcduLtQjCuJWuV5JlxYSPFwIWnrExk58U2zrTiuciZhpuUABGIF/Q
N/UfAWQKDqf0Q8jgk273fhOd5n4fZCZaA6I/ARzQjEh98jWJHQaFUWGZMux7JnZdOqrhXXz/0hhr
MjBMXvO/O5dnBuR7SLc6xeAIn5teKRkQpvmGJyofBFwuwUDcOKO5oL6C6e+N7BHDZh+aBAim3QrU
Rw3gp38qE1ZWei2eOEvP4ycJSGty+5ObG6SXdczG4fS8r8ou7pfwBV8wm2RoMqN4sVk+0nczOWs6
N2b43cf3zAWaLRImz+J7cKWuSmWt9aWz42/0mmx/KPwLS1VNYI7lxlpOJkECgnPOpO909Gqw1TYw
1JQ9FzpblmAnBrSCu2rxqBJyCwBNJ5fpxxEO3rHtmtDL8/WEjgnPSbllOPsfK9wvXB396yfGSx0f
8wznDcyQBg7IvPjKRxwenn0ldz0drTbRJx7WLUCbBgk0VNXLPQghszz8isDO68TiR/1avTq/tMfM
Rc+V5ZbmjRTBpKV1KrNb0X2YdDODcHre05THSlnJY+TT/wvGa6UFz0tIwlqY5Q7YkhoQprI27uUH
2llcIgxiTSOB8NxfkiKbiMxdXl10EYPtEYELdu7pc89wD9+yAKOBPax0mcy6/xKoZ1KKlGLUQSNs
QQo48GMvHpG7wF7RPizKLsU1mF/dcaIesTIVEyy4ies93nmLJJFZWo4sA2oBdSN0DRcVrdPCXjSW
qXFwuDR5E3Oo0Gxt7oYHNgFrJ4Rbkjn5Ac/5Sp/xO01QxTYPiFueWj67CHxc4L6jeVv3k59sExBh
C5/GaAkwWd4qJXtuOZZ3oZSHOJGNnh5TXWY3ewh06blss2wV2hMNFAsnjF0ab+H7NgFaffVhAJPO
NnaHnH+a8bOBEnf4mE4sqdIjUszZYA09s3FrDEv6VfxSyo4bRG5bVEWY43NJad4sBZsCp6DEYboB
a8pLpe4+CVbhbgVZfkVTo1PXVsly6lBsVtKw1EHdfSBjRdcD0Y2WRe2lM2xu8ZtDZ5e6p2bPHXP9
J1ste5KzZp3vvGqbfYDIi6pJ50ZsfFMRQKkpvzse7IaQOQTQON2SONwAWMHek90YuOqvAZQ5vhTz
Qno/tb1L7PIMSSJW0jRXRsZDRHd3a/p/eXShYtHSaltL8xjIDZ05GgOxMewnuE45nTqRRoFgh4c3
kZbk3/9GE/yL2Kh36FyvqfEykBOP5DCJwi7vs6vr6UaihqqY2K+kpfojn1kaSncbRnsbA2KrwnRn
ixaG0eUOhlIuYyy7x+zh4Ad7dHbTBLRt6vrdiXTfwYax3SDih73XavIOcKed0kWZtFS55DQPtrsW
VvKLL7VdIykwc2/+ISeDApXQrkdN5239Wvma4eLlVnJ8MSpSsaqmxwdzVF3qZAKn22Fz1XCOP+Xh
ByUVvdtPYqzSeDgD1VqB8/9JM7YPvAijR/udwxnw5hVnQcXbIKteRAQ9KjuB0HF3nxUVFDfV0XvV
BybNiTdLaD1visa6h7l4clH9nUTcgAejTBUWMQYjlPXS8Cghf4rGstoWCy6lp2a8/Hzrg5/lcMGO
8jcUXBkr020jRjeJ3iCOzxp/U4P9ZEIGLdCmEiC6F6mqBQwqpzS1y/SlDQg+7OcmTwLU9MSGJeEx
1htReRSsNqPLmYI/VKznCM1CK60oIeBeCGdsfdZB1iQtaUgU/8i21VYlxKDERK74ql6NSYYOCjex
gApjyNR1Vgc8ZYE6rUEzKRisUtDrxbyRIi9FuI1UCUkGXDuWp+HgKiu2v7GsECraDlLqQQfzNZpD
joaM0RyqJcUS+5V/mTG/2JBSs2NHQ5VU+xAzl92p1JoJHiNl9gzswRYQB3SOlsDXCRkMQ/DAGh7i
/2izjbOc8fsIKX86MmNf/jM4UKrJfFWYdvWKV4M1ehlt74FhADLEefubmXKserWk8FxyNxdHKOAR
Tra/IwkZk4xSkpE49+jrAT2dQmJwlpU4e7PoPltktZ2G8kdUJD1ycvSGiziIz0KWKdzSdKb/9ViV
JkPk1JxfyNtO5+O77jw1jktedauA3pIiTGLm0YqMMc2nDyKKsT2bKjQnNjiZ6RVl33YsItNdO/+r
jpJrVEx9dUKy/JDk9rtx6aoSz5/PwHJDVrVAnD64pLm/QxcOI7zIuXWZ1xHUnsDu5/F03SPImJYn
FcnpbrwwhybVz0qRHs42d7322YF2GM8Vqil2lfCuU68w0rMzfbfzlef13kKzpeLh1IbvOlAkddj1
3wBB/wxXpd9EL0UqgzxwJxb32zWvfWdrLvO9CQTbY6VmAI09XA0lP6ZzlZzsPqHoc3w/9EIDRXBn
azOfbAGvdGeo7fvTtfIZozMEH0gOX9JGyalBzYLvQGv9Bd1RzFWc7WMza/x6UhaFyVSy/UmRvnBZ
htiH+hNm5+h7e6g1wMDV68S0sQpQ7psC22I56rVljGMW/7cdVvXMeE+nQzWN8+1AkOs4JvN00jXw
EduxcITPcNcY6HF16yrDiGVoe6LgpTRbReKvXr3E+9wmITe20f1gpgrrTXeae7G7eBV1PjikgGit
MjRbjaFej6eMqe6Re0zlR0E9VU0+gXEIyPmsIUe82dow0ijUtdEe/TKaAxFn5MJJARoo3bYIuVL9
Ge00ra30gbFtBMXAohCb/RvrB//SQGsLiraxpiGyqXZDcaB3ZSuKPg9Z4Nlw8N+RhTeI2cm3gYHU
9SkYxxVczaqKOfjNcWmYtHfOZbKFjYJUA3TCnslLGNV5huHKW1vkKp7YuXitlEMzs+4lCwV1Wf1m
FODvwczeBoBDwsFYRre9SVJ2HsV1dqjqlOSgi2Dm3F8vGJnha4QqQkxd3GK6ApWJU2bTP6wvBlKv
c54m0evLMXm8CD7/Su+BNSnSqGqI8VMGVxdUUGaPOYbeI2xd9+QvIFHg/FXACv/PaCFnTPmRCTml
O7S9fQZs4MKpsEPVNi+KidXynk3/lVvJoDSsyYk8OlneKWVl4yAcCLQm6Z0hYe+saa+bFoFubopv
kv2tC201g7iJxjPbqoVdpudNtII6/ZdS2hbdxC/fWmhEJwA3JxKTwWgF0MymW9ecI09TUNRS0Wu0
+6YPJ1LWmJxWtY3umCrqasv7LF5vzVPhFd+A5ZChhOAiL2FvO0Zs5qx8A0YXcZy6A6pJDqfybzv4
Y+eHVsejnxHweBKGr6OQGz7s0Fj/WUBPP5NX4brdkHg+N/RHyEYmzVZzw9Ea/ZGpWODH5sCDIEZb
n4bORWRe3kFXUZCoiOFBmv6QuPnU4nAxEjmJAG88WBrSwV4XcvBuQoJ3pE4u2lYbdUIEFpmViIgO
ltxhhMwIdg2tztctyxKCVjkk9earQxZpqhVqDtnLnW1pglI5ncIz4zXxvo5QvYd7LuyCurpnp5LS
jZoHN71Mb+af/sM5cbpxLnd0MMhPzeZBhWUPxmz24uyqce+GpHgj2JIq8cr7e8ZjbLBjpkqdqEFR
tnzN5/x96OXZIlFLPkcN1oB36tPqBqwRnB0j83DLfWcLab0EPr9VcGSpB6R6l+znW2STB9+DIed0
ofAo2tIG/F8FSNijIDvWvCl2xiFziJth443zzbWWag22BDWA/teVZ6BLh+9aPDsTi2bMiWfq4Z84
rPAZzpGNNQa731bvNQ9pULAOTuMM/GsydNh9pCUKpMDcCWtwDgueUOUMRStSj2jZ3lyfPNiiNNSM
ub/L5dL0ifCnfn4u/PNMiZc8yAli+PElJ922bbSqMvA8s5xWCaRyuNTI2hLOsClucctBtFtNmu6x
SPnFrJug83nek/FGSwbrQJvi0EqDyBFdJbsgIcGYukWy1sP4Cw4dG4pjT4PlYo5InkQ29Av85nTr
4rLnc8/Mnbi1eUb+0MLrvVQVoeCE50OKpn+wUTT4eUXT2F34bCPgK4wjjDZmdlkXUC+eCa1msonF
of0oLY+c3Swla1RvpKc18TCNyyDBOJP8uXFDG+pBt95JIDk6+dmhVyRvZHABJ6Tj0dT8awGIxZsd
GBu2FGDpNHftkQuf2imseEfqluZKZRZ6jdcRW0M2WpbY080Qlc7QkFlzcs8nTOq7Y+it6BcYBHl1
HXxTNZxiCwX0qgZ+ZF/gbDB5GS30WtXCGlsrPKTQRhaWNaAsG/nQ5mKfU69PT23qoqsoLpse0Mlt
1GHK0lPzk8GuafUd/1bxYeSzFamQiZjxCn+BH3kL8qQqBgejB0ZHxIJ784ZarLrzgVr/TJOXb3z3
Pg3/ht4k06LQXl2ffr7vxDyp6ad/AOK5rDTaD9IIMh/c/25/wbiuscHaJJjwJwcdxDEijpiO6JrW
ckxu/RLmNbYIg4ssdsmWDsr7nm/5EXLHrkyVnLif7OK8gK1tudnZrUdARuzh1fJotDlZRb+8YZZR
PdjHaTC243Ta2t6zfzK6fFLWNQuDlSf2r4VyXEWsmruYkRrwhS5iR/3NO6tBlgWQ00Ky5jc7GSzO
N5vwMr3Yd1zgnmR1f+mHmFqXpD+EJmZ0nUCUvj6tF4+n9eUEwD2TbgDG/qDVMPGhZsG+7l+CNCCB
oX/LsXudOUgrYDtzlXfcWleVBDYVX6B/ZZT5vG0tJNGd6feujEw6aAkkzcjbbSWyhDX7gaHOgLKa
vZlg0Ej7xck7smkIUshrL4BSXA2THvr7LA2uN6zNnXYg1LSAPQ5jjAJD/aYz+JYuznL7s6Dg7PPM
CZEb/V148w7uWeKbJBU9JNIOewqU9+ILfkJNfFo8RNTIiJQo/75oEluSMcMvMS/CWOCtcsO3Z5h9
L15lVD9qN2rALIb8tnmiShEqoIkco4ApNnIfC4hWTjapxKgBO/ER8na53D7WRVmK/CdyWjqituyB
9ZL7RwONWVVJERwOHfXTwEs133PV88mRjmvjfFT/d9l7WpP2YS1PA+a08NjQtHb+dScnp5or7T1S
94L4EOqDHjZlpFvabsTdN3xQSWT3RFuKXff/YP46ESh6V1pLJB9dc9Ud8pvJjZ8iOtbiHoUQKZDM
mgGVK9T63zINP5wvCe1Pp1ftTZvrWmf2IeuPHBIcKeUWX6bTSeRWbFl/ovFVCy49u+GnA7uBRkya
M3jY47IQKhkDC06MHO1gIMl7drO+nYfxPfu7eRTTDrwDDZpcwoiToiWEX7kYHr8bViOb0UUbEUAD
LDM1+GfhWjBh549sFOI8OkFuJA3loSvnHC474kpt0lE2XBjzMoex9Cyes8w/eOVJEgACMRW8C8IP
VhU1FerPOSTxQKH4cIdhFS6VRHjIClUDlOSlRvQRVsmAb0HXtBmnQdvtttdr/YMEUlj40wDLKLPt
BtVdx0hTNFm81+u52xJ1a8aJbNjJQzfcVFyzRumkRrsuoUCF3V07+nELAAteXUz62DoVl5TnLIuq
xFfEON99VNvDlRvN0MBn0v7/45EkvD+N1vIcFNcUpnID4PKGHaEuSsRZ3zEFvo9gxR9Nv5ot20bB
Z6Xwpn+pnP9Z0nENibnXIGXTsL1l4hBZHFYRhBQo3kusocp8byr02LZ8qCb7ei09k/ZLO72X+2lk
KYKOCMnlzqbpG/gyF+GEM0JaNa0EObuXB+U7cFi7ii06icE8aBXoaFlTJChqfpSPIeEFAzqLppPu
DB71sIjUAEQg+TUpYuMbPg/vOxrT4b5UZv1Q1VQykm0gxji4xvLHbAbFYNoRUABes06GGMkpfMvi
cqyW9xdzPCiNwkhoD9w2J76S7J4N0H+h1FQLyb6eXVUWUGRSpEQV6nFyUXuk9Uh9mx44kjqKl4TN
fd/VAOcWMMeXqxnAjVI1o0RNkwXpHjP1ER6YsxmcfOQRRHcBySNiEYMRAzpDJdKDdB9pl+Ppch0H
hm2v4LxD20HFnLnAmE7RIuIEeFln9dlrQltSaFkPo81VF8yyywkhrM0wxUCpgNq0NpAz3s+eKEuz
zA9p74Tsmm1A9fetxPnca8VY+hVDW0w3qQGv+krJkRpamELM/w/5Tg0V7L784wNR36fQrijIizs0
Zq/X5RgaQAs4wS38IgrOLe/U5+Aneg9ipn4W5cnMQENZtkgdDrCH/u+oc8E6UQ3++b46Q6ibhZVR
CvaEp8oXapyTViy+gJV/i9twEtt04m+PqnShaEKOyN5B3JhFb1Hpie9pupj8jRVgkf1Ypq21lanc
HKTcHa8twQXSk2hIWD4gFBT84aZdTr8kJz8nuv6NR0Wy4Qik8nUiKJL+nH6t7Ag24uDMrJsiku/i
yZCuCY346BoovMq89pvdmQlqeCfyJjy76klwT65ZxyHB1bI/AOITnB3DsfGdiMkt/UvT/pFyPsb6
rXtL651KWpXqFssYMrTHVnWGApuF8bT/te5rdD5seywhc5skeJOmbonhJcdV3JcXligYTVJxdhWz
ab8fS1UX3jC5yx4mCwHW/U640AOlfqJWK8Lezvy4o8xmoYICYJwU2t+2ncVKWigwzeuO/4fW/1T7
CqeMKWsHPeObd4HMN3KoVARobnwhZ6vejMcaBQFuvuQKbhgZXHXO5Ve91jW3biQVl4VryYDxdVlB
A8VJ57YguqVwHzGoNoik+tkPDfQgIHJdH9dlW8qlYidgej4BPcsXpnJo5M2+MfbUAbOb5tnn/lmT
ewBUQUrEBOpxCJ8/38SNQo5WaUEiEHjw5y4z8909PNC7QeSmegc0y7q1bibM7KK4N6oP+7ibB65E
S9rlnHVMiRFqaUZCxuOvZKkyfKlRm1bAqPh5ARwnyWNZStv4RC2nzm2AO6CU2oPW5KQHIeUfv5aQ
0u6Rhf6ZO5Y6CIDtnNG37UemF8bzse+f0PfzoN/0NxMeH5KiqAl4bI3B7MhRoZpuaLcfZBaY3gjD
px8eNcz1cYCGQrgP6ohAShwxghIZt9xpuJjTxz6XUKbvSSAIqSG55j/1EnbBT0z4Y5VOWoGUL7en
tRI+2Fhts/Z3zeLmse12J2ony0as9gsdwUYqfmbvRe1iqyMHHmVX19oWMDBBF66/dHd2z/Z+EEaQ
l+A+t2dGjfDdoC3VLaKm9xto3xRH7DPBd2xJ/40SL/ndsFVYyicpLvnY27tC7BhXTSTrLfGqD2rv
yKyv/PKwVjZkjrtnvFbwC+uvdK/RiBdPcF0dsF0wMejcMLYJKtfHZuPm6Tm+fo8TUUeZVW5fq5ou
gZrsXr1ul1qK/OY6u/PlcN3wzJ8k5/KvYNUhfMAAKQ3zbPVVvzS7iipg7w8MGw8C0D091fac2KvD
qO84NULIuJAGMF6HEZwh5xad0/V7/I4HLiE9/1jliv2aVlO6FfUWS0AoKuC8aE6292N1ioa4N3c/
7tatQjNT/Rjiqt8CKxZh6SFZo5N8PGSu5jXaEg4/yi/doUrXl6vHUZ4Dq0sBLcvCnIpwF6A4ckVp
7LY1XGqnXhpupvXfk2FeftzGeizqtH+HtO8fZgPoh9arf+1u0xB7ZWShFIKe5wxLM9+HsqSZB7GL
2GmcKDhjlF6ffdfOBEFeo862aOHjLik7Cv6v0tkJYvmotoro+F4MPXHWuNPDdUXzQupDzNVgNZsd
xSGxkuF8zup6XwI/5cfguluGMSXCZmEh3+JdK2uub4JZPdfmLA3UgzUbafpgeV9diM6MP+soJoT0
wUgbt6MY1/1/osvzV6FuRLI2rwfQiqzLkEl/bprYfLCiwa5oad6dbPCIXcBMBrtJJXUKwyRGCOcp
mXsQKVjWYE+Mqw8SSMBM7mDBJrHMUVFofugCsGCr2kNC/uIrrSoVOWS2Y72BzavcuO+WgHw+hOBt
/AeAMHfPHQ4o2SqkqBldor99342BalPlwAqVneTwovIaFRC5dX2NI+skPNxvZqDLT85Y4NXIZaY9
seg2c46psvoU/Z68rWbwHRRULtLZ3DwoLxYLpZbcZFvZ/eNmzLdgNdLKoDwAWOqttPGHDoY6qWnZ
Etss2W4rIi0Hf405m8mchQ6WaatEZ4L+kDyOCH0Z7tTTH1fw2tewfeGaM9nf2GoUwYqpefNOixX2
xxHabJwsnFokFTyRk5ciE4jn+A/66gv5FRD7W9Ghs5JE8AjwX6ObZh0Yu479Mix8Fv6nCKsk2fpa
kr6fsq4o8B5QALQiKJSIFFSkDlMmLv/mrYeNgQUcD8QgNvUiRtOyPInvBuz0+D0VTbR3D9sH9L9E
g/qwUvWeanNgzHCsiytgdB1N3rGmdKjtHCZ44h45YC6KaWuSRWwdgGTGGzlOc+JqNze+7K/1Fo3F
/gfLhC7+o7cOm91i3Oj0VHVcVzOQ6UjOhccFWizVVvJCZoyEsrJoQL4vQdYsRIJCMXIF3IBuZnSk
E2124gS9NOk49AOU0UamYwZX38Doi8oEXYSoFxnIZwowd0700qoNLqjGKRe/apcVRdhL8NhJFuKZ
7ELCyDoADbfH284JsUO5MyDHQXOGdA1zGKWyfGhCKsRsV4/NhNSuQwsXctZ/uDsBsdYDVr6OMVE5
GAsSetyiooftXPDluK40DACAfzM+OmkjKY6Tg+t5rCJXSQLmBBQhYGudTLNnSXqeHgSXxTj298+r
riwODSgfjyQ2An02wEUc4lRa6x864tgC/IIMcGktDuewgshvZittDgQ2Sxcz56LSFEO4gzEZUSva
vVs4ySUe8HEdnhZULPomGtA2lfVGQaDYjDLmJiNnp5M+mlf08tINGGEtEKLvwT4Ksf387aymXedD
Zp3YhblRIuuDdHbiTlLukBOsBXAo/Io4V6ntLPiZR+M82CHYBPn1zDNQfejocmC9tQ8T5kEuxNdu
MgZYUKAOps8zQ8KmmKnQNfdRd+rTbnqfO+6gczEIlbll0VsGrMBXLoMtR6vGUPHlevCCyTD8cirX
ZkJ0tZ0aMIwKDYooILFQ9mrwwBVxc+NHQ/DEAc93QQdnAnUMaMYXU6KSy3aASggg7YbAuU3FEfBT
RP6VEalgyPTF2Wt9uX8qSHH3fzFlHluXrSuGTd/rsIueoOGgAtSqTXLIbPJDP75g+QbYbfbMrW16
KTFr4KJ4yN5Wjuntud0fwaoamBUiV2llbLletOLTo2WobOEDJrmxpnx1p+/UpxGm+XEaMAK6peoF
BL5Owxuk7RYvK7uaG2GmAyuBurlYyfpzrP20X1c8BzGwbCxnRw+BcJLMoYsNEeldO2TO97XCqqft
uoU09J11Km/qkn3iYq4V/7I6IF+jB7I30sdwDmRyD8H57ThGJUfssT2eztIRzd/zyQL4BQTqAHdJ
HPar3Y61dTqJRlAjk+nB6fdOQ6wHVyQ1D5FnQOJCAz2rSi6jFj1sg4wWbTzkiQB2gncwRoZVaDcH
PVkznv2XLvsZre/daUr4ISvgMHhnzifG+Eb0ct0uP2kdBQGPQ1ADFYnemzj2WYxjzMvK8sitgmgT
1mVAFNIf7pLy3S+tsb2nYBlJgzqu38jB7mJbn8/YqabXJr7/N3qr3Xqa5ozUJf4TUCnPlH3mV/hk
jWJQ4PZRvwaBEMurnsl9QF1PZWWta0frZ+gwtdBcpG5j7YKbjoFAneIo9ZOYpqoJinJ9MguTQBPj
lkkS0JjC4HRNbF7lqCliK2ReTvq+qGgGKf4Mzz8F1oBRkzZuCaq0krZ24OnbMFUtAkgjVPrVQXy/
20/uy4vw8s0tOi5YvZM7WL7qhR8qrP1sggeCn+qdR71ur+FDIMyTWiURKgQW+dPaSNdoEgdalc4l
wqbvq0oibbUNcAsWpYtO288T5GVGhYZHoP2mn3JI9yWtAOKXO9pRdYUPjSFFs5hi4G0u2sAsspug
LmQI8h80lE1GTFDD+c0NxymEYhYZo/EBwGlGdzGQVGcMpyZcOs81HGF0cSzCU5bRnWV3q1lL3gpc
vBmMXH+yAceUGIZwmlTihI4F2Ujah2KY1U5hnab653LfZB7djB6IXMoKwWtHZU6O/4PUpnbknIuD
n5U2zLZJKV9stIZuEevC+KSsojEntUQsf7HuZkBEU3g6FKREdqzLWc/x8FiVR8CpP43ySTqvnRbO
2tkKYXXCqMKTzXSrNjAMoMXq1TqFWuoQl41oHphD6bq5RG0XF8A5x3t189FdQhDIVwiokqvEJzNq
7bdX0Z31zj1dlaH1NmwfZbKz3R0NkB7pNYtcYFensETlIRBd0FjAIZsLO/QevFt8JRALYJnm1TKq
ARsyBDLUwBmmCJ+imEqGUHSK/cWyzw5Xlkg7LT8uKq5SCj65fYYp0MjQX0oDXmIZZ+i3lye4eEP6
U6mc0gefBK15uyXLkE+b0oIVk3mlTCC/cUtI+5KL7eZFL3wn7+3B9XQ2hWmx4xB0t1eqwSkYyXfW
NNB0WSHq2QuikU2nzHiA4VG2TPR14md5FtRBPsKYCA9QtIEbVnGYFMp+n+5g1ySCM9P4rkDEofwk
/l7bQuFF9IdsKdhlGyJMetGIuwgoJRt0iN830BtHWovnm72UckRMG2di2V1LEvFSghDE/MugFFbe
A9rPmsjg9WRiCp+xpJ5VMy/58NckZg+lHUJo17JFeEDfQ5x0ZzDr2d0fseUcMWoX2TBJYT1io5TM
UGtC9XoSonEwAZYA+4zP1SayrvbWmvuHIWvvojz7mwX/5/UpLMPX/R36gZbqNGi3c/crXyxK+3Dd
/ZxUrrxUr3BelCwUOuEPnMd3k4se9L/nkb8MGxzEHPmLKm3tlm5zz/+TD4/bTJjgxj03xu44fLGk
N4FPxidwZYQlkDDgaECSsWgAT29kLkjSoUKAGkTyq0oQlUpA3mAGD+qnRFLfgEOYsCRRfs40UMYZ
S680EH+tTZImgicJhi/QSbUbJcZJEqSkBusoLKZOJh1V/TUoWpNQg092aR07/iLegsmCc+RFOFy3
uK3TXoOQn0fAOIgxGRpXt175xbzKOV0SgdAPlazUelAGQKiR20UVhQtWKDpFV0YTcw7bTDhSt+10
JEILStP+7LuaecILQGws1nj126U5mt0JmqK9jIXzI56rZOxI6IyQWPa/wktzdYyEKGMM/t1WCrmd
z0BYhm6dHSZik1DMmUeSzAnz9L/XixztcBfdPCTaD6H/0vl5O33pM81pd3WCyU2hDK58BfS4nTq5
CDFb7vKCS6/SjgPK2LzwL9o6WHzy72i2k2sNhq3uyE7+xvKh/5TQhhPM7PKDpJkLZkywrre/YA2W
Kd1Fq0Ybxc2XP4eVEieU+kRb3Zrud1yEXv7Zoeywkw0Xs/MAaKjBswt8vZnhcoef8x7KNuNQ8d2C
RaOX8WeP1EetzzSQl+Wg/0ou+ECcJN2+J4yEAeMYNqO3Aej/tMlvN5mBmmMN3WtiwiZE3fGtWHss
Rekistz37AEsyaCGpRYOAEAYx2NxbgT0AGSRcXPqkVvvyTrI45y783QGURcSNZVio2+H4ehh3mfd
fqKgEatFVU60jQhuk8W+2G5GZWyXi9Se52eAOXUS4HUL1c+asr9miWOVBg7ZpcSN7PcQPY5cM5nH
+UgSLOiiBMmIhDAEhRtCiLUHzz9o97h/9Em5EhZ3FBdQ/lhcK2ubL9qazrBVHuDin+MT3VX4GdJm
g7+YG1pgHem5Wx/+YVVau8Gof42hlwVDmiivxE+v69srHlCCrDhc0Ut9QNn2Bsg6XpF3Wxitabz6
Xj9rZlPeH4hh0MQmY4hRM7XTFaw3/kTnrejYyX4mmv4zjdldOYsQk9GXpnGd7utfBbJG8dKG+74W
v5DaDasbDJxWzXW9Ue4XO4D4KiXX8TeOkSakRbDt/VgoZJ9FsdyY3FRqoRVdMxVFSdGnSx5n6tw3
eUeFVExFUhLzZbyXuonYlKtFnp9p2QjVsmCwBFbRBJjhpi+UaCdK1UlRr0dfjzeaa8EAWTPXlg8O
MrAkDo7oi1u5vs1DccHQdEeh5VdQPUYaQVu7N1LqThvouGMnBOdLJa1XAcP8Pnq6/E5NLdIZ0DYX
3VsSV0ci3WQTWNh4qqb4K/NtLU+YojYgWGizI59yVJjbZAP8FN4K9up17cTX/HPPuQjnt+VEMUn6
33xEbIPRnRYR5Skpm5us8GZqSwlBTNpWNPl0pAHTiVfE6HyKadFLcdQVnMLRhw8AqGRB3atH7YEd
GynlI4+C1dky+w6wIH05TlUfdzV/wWElA7skup6NObEuslXaRUmjaEiyD0QWT/IDEGAdFJTQFTxO
+xouu+BIgqymmpU0bg2522P9SLNdhWnnasJnVwaf9F4sSawEskqxKhIN4Mih1cV4Gw9XrPIGSCFj
90j6FuhCXS1mR8PdAPhR70HS41WlpIvLBJAxHd6V8l6NwIylZyC1xw5ASV/7dVTdyLiXVjqQObQj
bqq6MBBAAGkBwI6wt5laS2pFqP6n7niHuI2uJbmrpQRf41GAVfecIA+EKG1nA+FooKjjT8AwKaA5
TnmMuOCUDtF9lLrcf1cH/e7n31pcNCUGlRd4svxyKyJHKz3KqL/45Qte4pfcy2jG+PCnRMfq4xCc
cj+bxTLiQaHjwZcdDJXB2lackHQ7f/Mghg3Z0UTT1W7BHtY3EyhF8ZT6vguphjj03/HVV6oPTX7v
1CVJo2ov3/t6b9U2NtBPrnKtoIYtZ5czEOFRrpgriRjSVQI5nrrPCFMivEIoAleqJ9Dutx5a0sX/
9e2lxlphMetxFqeyWR14yGaBMFe8IcZUQpBpx0yObEb0Wg7oU+kkzDzo4Ak/Qz/F7LqUZYXdQfxz
QjXYDXBmMyUDn9vR1LgdnUYSKNzWC2nGTwk0tKtgps+V01bM2MIF7iOOvUrusQnDGuA0MGiunYOU
f62h/l+doiVrPCF4FQP/HKvtCLadzCm0eLvtOfYXEr26T82tVx6lzyWZ8DCg7hk4QKYStHVCXPaN
EOOmmXbXbD4pnkWmzvRRwwR2OhrrPxbk9Ob74z14UkymH6Mp5Ls5/RkfWqtKn4Pq9Ho7laqo5DY8
kVQxKfryrH1M2hE05pQCGRCW+O+aMe5w2i5sVx32dGg5nxprnk8HPZYZH9IjilIFfi0uyPhMtSUo
W2LRf2LUPEkuUDcvwHGMEW0kXpS0bOAGt9MBGshUwvj9BwNe6SBFOdbl+wVPCOfrVKstj/PtLENw
iLxOKmb2uYEiFwpeY281ET3WYIKUuqFwf6eHhd/dPoawk0fCwCjiURYJm0wHxiiTd+NIDJLBQxA3
7LRH02MFB0fhpkb1B6UxuxQuCvmr1LOg4aJPGwdmOcba2rMYYuFAG9FGEBSlrgu/hacupjY4AmN/
akN/IClbHa96PGrD9MgylgB1qKFI1bDSWO4yJ3gzmiBq8lmZQ0uq7YmdfpHak2J7leSHIxwu7raH
w5ZvXjUwkxGoSVVMVtZxMPeSS2RA0EnCXVAiXd71kbiRLPJ2tEpPCJUqB4LsipNag8ZSzFWyP5p9
8bcL+8HOSWkT58FNLL37EmPA4DzKWw0ZPE/4DqPb3OxXALLqqZ7IGQohbv8yMqmHS1iBPgZ9I6qu
3l+IpX4lErSo7PrxNS3cZzfteqdS/ITRqxpomEFvyEoAETbyfAcszc+H16ZGp3eZrlJJrCZOtA2v
EAXGyTJuJuRySTyCUBTyELnmhhELd4TFMgfC+XDi6YaXwNeNTpzPqN6QNZYRX3Iq+5clsSG7huer
TRRTnAw3QFA1rH0P26iejMHg1FNmFYlngcLA1CEop1OIZH2h3jyCS4SVJ6YOx1KWFS+Zi+t84xC0
F/co/7wJm47NvxITTdy1TGCuBll6JjSiuYLdQjqoIEGQN/AJsf1QhKg2Vm5nS7mPe1X9RfUHCbH8
9Z8sOp6oNMAXVRXx5qwf/IjNDq2wMJrNWOvkxQLcIBuEqJaaAZT29Pdz271OE9kHaaE/uj5x6pfN
AKpM0aamxYeijabQfZgcU0NcXGcga3AoTdEZ62qGFXvYHd2f7DioUhpAQXUHlUSTjVS+QCX0rfQm
Jd6c5xSBDU+RIgXsbQn39vZwGIPeKP0sfh8x1k4j0u2UJrSPerY7Wd595eH9nBF/vN8SdajR1lwi
TL1ZSJDdvxA1fp15xsuiCH2/GaLj4tefQxHWRDsENi9G2oT/4Z5yxkyllFbHp9eCEEGBdXzKgaWh
c4F+UMx9A4CK6loB8AIG+MyacLCXYp63jOZHcfcqfpQHfkaQgyLDHLFxYXq8lb+G6huAfWUWSeDw
hCIq4La9CZ9A6fNdyYNkxbFSlope9sRw3pXX1UDWZso7/nLV6KmB6mCQTyxQ0Nh9M+Xzxs4m5JcJ
IvT7pBJAeGersfoJuHQC2LA33RIgM5teFyoH6gooKJBZJyuJTiRLglY8BHauy+XkJ/zZwtd3c5ZE
+B0I4fNzUBp2lU7ZKwczAioeNqTCfctDyex7APCxF7K/jEEKbrc5/fO+FVSu5JOjTSlXj5hJIr7H
8VfJKT9ytHfbjX8CrSYOo2sWEkQBhXqYHxA9E5xQJteVQYijXVGfPMQvA2BafG/yuWz0Y/ezRO33
Hpkji9Gr5MTU9CbenDyFTWiuQtCOx8mNLIi0Q1VtDvW2tjCTpMlFxvtUqJn9tNb41+A4FJOgBqlY
GF2K8qlkDlOxGTGlj3+Q7sr/AsTj7W38pt6iDDCyxAJ4CM9dKU29HjG9PTBuJdQyfw0anc6SXf/W
UCOt095KUCZZZ65x+yaKmInICfeh0Xe3C5rxbSqlMYD23Dx8t9E1IJXN0Rlr42sJOUdiH+DqxOr9
gVSV0H1erHw54nJEC0tt67f6dnx2WeFO3/GY8ZoCS2iC0SImLP2YLxNMmfOjzRenU4YylGQaPSCK
KrUqLnoN/ZPZEyJPGtZGIXB5dNexeBr0l3yEKtEjkVqezgLPzoETuvoDmFngu9MjRQkQZMr7rFak
jvipjERcNtEjku/9C/yk+C5F+QRSm5TBGmIX0WT3Hy7KQ/8lPq3WiKQnvfp8xBkxmXb5MzIJR/w4
XR19Y/d8Lihq5wSiT4HbwasdRHmTPFnhEjAwMozDuE1znszdLf8rrXihYpe6Imb0XWe6Y1wJ2qgQ
9dDFFmoFm2mDsFcS+ne+jTrWswkprC7L3X/dQmFsJVGkuGzejDedU2THHdNE052Z5pser0t7/K7F
JiZd0oE3qzaTeqxfqJpAw85lhF1ynDK+LvgsQscWrYZrTwtkYvArWmMEO1KanxpBROKXCNoV+wu8
ZI2z8jh5IMGHZron9xt/xQvBimesyacinELuTnL/dL0lPRvl2nFKzAYg3NSi+XQFC9lnyBY3ROfc
xnAkgwHILTAodUcQF6emcP3+AbzgE3141tfAU62EPqDC6vJQl4DiOS38AAXz3Cp57hnP/fUdVCGe
uF4yRRW29xxSR97jt6h2AKGN+HViuNJ9U+cSSrhXdybw8VZU0P5+9B8rmLjvWVUEYdRhZrxqaeh8
3EISzMAdjUDKv2s1Z+t6DjIaY0mv1/qoTUqYsJflJlMekJP91RmtSCR0dze6rqG07gngOeLUS8Ob
kU3sf3unDAGWrfGOZ8zrM2zVr/UapmbUa74fVAbWA6/IJSsIjlyQnvDF9QESg2wwPKOWXpe3JxPr
7YyMStnoZYW/ZlM88Tpa7I3zL19H6diZfYu1bbwCaFMNSRGh8hxXGWMtdLggPmNt+hn5M7BMcdqi
yMUroQUs6bWNk0/qH4m0MnXcsnO3BeJlLwTpq6ozhZtbLxGWRz4BFJo5ZjPSvDgbii/TcCwt5+cu
D4mx3lhSUjLlU4V0kgfF5JL5vEjkC1hTZmNmQp3pOyKZBWnmK52Xgswri7EEzcAic2X3z94tHd3E
NWWznBJxQpBbEMJg1NBN1Of6RF8/Y+XcVvgVnM+68N/ljT0xEt+PKo2jRIQRaZsO+PnnFhsdyJfh
5MhlhB1z6eXogM8AoB2OXjqikBr4wtegW9zm86DmSSDOmqmwGHCAPAQ9GdARt9sdP/8iOVpz4K9M
i8c3uI7DunFss4elSnoSZUgJ0wUUQrQe0lVQ/r/FvTiKVpv1PCGgz40S9TaLGfyzzlBsEx9yRFCA
jypG553pqej/kyODtpGU000Xkxa+2L77lpUqvJhbiDjsgCsG466GO4CwGeVjpZuHl9BVwpwf942b
h1VY78XtOjVk9qT22K55J1lYaUG1hi5mzbEHdpxzQTEQt9xFsvbzd1eBfM2NfdaEaTrUeP5XuLkZ
lQGhh19Wr1ryTvGiZ1RXChx85jHqChhroHftZygg59Lgp+gk01XSI/es3gcnu/Cj+OyKlebN0Dl9
pfi0ow8Vad9PdMNYy7dm+LVF6aaYajnZc869gAuKYnxiHyvdVfvS4G5gZcpxlz4k3UigVvv3stsa
TzMDuRzaJaicT9FapgAJLDXWS1qADuCJMoe4m/+qlbHvj093CtTfexL2kZHQ8fdTjKFUswOqPSUa
2U0gd/WqHZHlt6XSXcgNA3XmJTDp5gLKJUCCh12s9kCQBp1ZiTmEiLIRku3hT+UkU1pNhInA+aAG
rwKuKtlv5tthMEU3xjjl2SmSTelmCz8Z9WzgQIcG4YMJf1IvBNMyb8zmZNdseBb5alS2QmUU/zwg
61N2pawGhRDSEiU2br1AFwHW2QcGaFpskRFZ8K/efN2SARKomcT5p/R3ushYlgqoVrs4s8jjm5EU
1dKF1mpW1DimQyuVpBTiQbPSaMJaLm/eKZfAFEJB6wilclJimTkFZ2bB4JPSV1gBZJJSRIqkWsHf
2gGfW1Zjzb1Z8qkTxlDtZPDbugYUog17KrDpAxwNT+PSdcKvH9i0GAmG32wYhVoI1NqkGJOqAcV7
cELH/DI5oT6tuWi6C8NPsVNytKWVPDd09K70G4/Q+Zkc313lOenbmKfnT4XNMKHTBxzOPmjhi5x0
S1KfSC1XET8dLwbME1OJbGJ/hR1oAFDl7C+leKlH45ixOfyCWX/X22xI7bqMMA1tzD6dmkYgU05h
CgtHJCHXJhBlXZw3NTlXpLnk9VWixv8m/L8rg8gJG7CWwDjH/DFWQzHLVeXKm/rxOnHvVyxvDoS8
4/P2/cWYmRqEvbW5vngkMqPF+IdRPHPehCb6nbEwTSTi+t0yRRHazOAyDZxzFJmr2GVmZP5Y9FUt
zMCxqbXZOahYEBNA2V++tlIm5kKFiP2UyJRJTeuo4vHvxBwO2bjnSpoPBmoBjQcD7hNEp/pBISQR
uQhl0Lya5wmvRCH7P1MVz2xAICZ+AwNdtRYYZNvUQdeRMNrrzawtzTqOkdMzu+ZqeAc1iXBzxZof
/C6jHlAPKLoiX3vGzb2f4TrTMgi5Og91BflzNHD4Y5wbe9QK+QBmPeK3PKSJctdlzPIgrwclexC3
9l5fc96SrdKNf0I+ygVt/2o98hziSz+Zrusbtf6jpFHdqfT6gvD6HgRy8VLKZjLgavv13fjfOaqU
vIyWw8KhA/ls5bSW0Z9eTThEp1UDF03S90Vdkrh5NSuAx+dVo/o/eQoXqSsrV9YNK2rUwTOv7ZAs
75myOUt8i4q3/0/C7YCPeDQQcguMhqYN9jXHQLZgGMNe9DGIBbT9B1WoZOkjoyX9h8ofWSJiONL/
MNjdQSqlNrD74TSHvdt1F1AYTWZ7Th9AbgkaDDT6ULGQ4vHJVgTA1DIiIDAuEhLuNhEFqu7umzR1
dwMP7+3K0rUTTZoQDClKuArjSliTU8fYfjhu3h1swZ9U1+t7ngJ8HV2wL0dRQJ4EFD5ZI8M+FW7+
OqwjHX1iAtVxZn9hp/Mn/wpqnDHLJwmI5+NfN/tcztod9fmkO8UA/fFpaYe0jerYk+Fw7ZFQd/b2
kAkDwz7gGmU1w57E00rCOmdeFhDEyhK2hJRXqeU15YhW+rv1DbtsPvGJXamF+RmP+Lik2Qm/Nsp8
0wg5P58bCAakXDSQ5IoMqPe/gDEZcs9trp3eT2Q2D1dYQx0QTNEU1bLmX9vr9qVlXTWvHX3Ctbv7
ldqdbF7BJnXVnAu8RLf/tyxZA3xKokVOm7xnd7CXawEcGjub/8JEpTIqvnTtmI8t2ctIdtg6YquW
8yenGbZF5rwF1Nf8JSGsdI2iCbkU0+EY7ByArJUgIYKPjfPCC7oaC/yJUQyX5eEydKOynQlIehww
Un13cjZz5ryN4EDArQdkprzMtUMzx5yxu1q6H1/4x/iPgUsuMKzM0+bEb4LkiMXUSqNG0AwOVyxf
9WXlZf5MtboDvjuu348muIJDy1a0iTVwaBoYevC0BgF7AyaQi2uSCSSCW+EdQLiInSL0M1Ku+y75
+VGpj7nbjFGDVmsGBsiv40X+tAeIJrhM8RlHoe5Wdv+kKZ2Cmzpn0bQ7R5oe2KXVsvyJRfuNmqP9
K0UBEDl7ZqquFK9Jpg/J7L6UH8A1C67QGTcQ49BqXwz+gdsB5hpFQEoLKzKfs6UXgwlLf4SKQN2J
vp+kKkfcLgHbBbOcfVNxkckVFSnNuFHkq6vdn45lt5T14el2pbTyNaLnDG318XRfB34kGRmNvWsN
/t34Q3PDY/aDl3oWlZ+Vuw3+ABMPokvamy5m3cyiLKgSIfntwWIl0KmJuINjmDTuhgT/9hb8yNMI
g3Uabrwj00pBuvgsrTOI7GGOR78ixRAgwP5kMTFB6JA3usX6CUdZaES7fp6OujIq4ACBnoeLq8Cs
poU3FTBcc3N2VLWpj0GCerwx28LvKQ8cq/wnqWFMC5k7yrvgzeAB3GC0m2SjRNTTb2JDB7BgovJ0
aJwW2DzK2CIvcymsR5izu2XpzlKAry4RHUMJoKFpO0/0WCIjeeTeTG36bMnkxsf6+up+41Jbdm5E
Rx0tUe/9OVUhN2KJOGFWdMmWuvpeQPOGOW6hUVF/asT9mhrg3xq3F+oFkYvrjjuNTJSbqNYRL6sS
MjAbppaozLGMvWcaPO2RFnoFutDUV+TQA8QZgtnKzbV7fVelipkZ/dcADQNIFLioMQE2tkERcSTL
1z0Xj7FjFu5X/OApMIpOp52rFthMjcRtN3iBBb8H1c6HeDWBgk8+weKGnkaIOa/Fudib/JmfQcOs
kOTua5A25L0N5dkE4gpYA23Bac0Pv3i0iCjiQFQAVfGbFz3Gs39iS39s/fnPRNoAeaUnjBVqgDwD
rD111Oh1RV9ol2k63Cyy0MsuW8HOSRwx+TcFFYskLrC5TScY0f+bM2436i5N9yhI57z7k8sd3ej7
gR95zlSVvWeJBC0KmbrpPRUW0nvtJoaG/0Xld9c6rV4FCL+nFAESJ4dwhRJT0GCTx5Fh8tf2RYoV
gssCPUb6+ZQS0nqRGpT6YzB2m8uMTRZ9MdvBhSiUrPw1TE3Y8GWRK+fxDzqba7exuD01r5bj+OIg
QwGVL4DpQpp1teXAgBonkS0BFlkDjIg03MtLdJ4ipGzfRiwQJiFmoQZZq9/syS8o4Qi3xBxx/WWJ
74HQCvl6cED6qWStrDZfEgrOF9trrcApcYhge/amCFbRqfACcL4yyxj2UHpx1e0H1S2QI7jBaqqO
nYTKDl9h+g7jWnTjuaabTmYD7UNSfBwHAw+5OIfuKaZ+qzd1b+dnUVd2lsfzXlkWswc/c47vu6/C
M8lZbEI/J1OeVuWoRaFEtAcf88Bh/fFqNUvJqsE5Z64UuXZfMZCbXBCvjkj4x93mtKz6JwWIWzg+
CZ1AkPd2YBVMMmC+lHYsCiHBzpPOAcpO6LjKzsjs7MEBwhwrp3vhclcrBLvVx4tEA4XXdKr2WM0b
30L2Pyix8fJdqPsUFXf2dzlaH2yeLhLcTRmp0iLVITCgU6EwvXgovQlibxP1z4cfgFN4QbiJijIM
yxwoqytys+Fx9tenbBCoQpNPpZtQVL7GUUJDUeAjRf0gcVrCVueRxleJB7sTJevVgyLWHB3CkNeJ
OtoGBguzRCY/LgW19cfFnJgtAc4y/WuZcBMQnW+I2WYhtMct/WRuoK+/bZXcl+9P3Kwek+1RCSLC
2MM9H14wtL2mooybwox8wbSNvaj9z6+YaW5RxTtVqerqX2hatlLmAWkRIfcNpjKXkZU1OA/Pjl6K
2vi2VklEbvkbUYxYePTyf95PwpSP/AOyNkW6SQiUsFPmDbTO68y7ZZVCpbgh5Jhj1l+W1YK+7HfS
N0vGX1DD3Xh90SZnlffTcRRahiAHTGKMezCMJG6DnJVmpbRxH/x4moc0amAJp1Zht2PRsl43FxQU
O3FpgVLMGUowmtH4Qkcz1CDslojewUjP/ZKr63z0nLrOC6cBGX8PAAYNq+/ROdFyn4HWZGhwM1TO
2r1LgULiuyoVyN/Cqj+tqNcpzsflZUqyInPrM6wKdBD9u6Xa9rcbxCoM0ZyaoEcXaysGCjZ6c0ZC
cYEoQO7al3Ik3AhM+2V8EI5soUNp3saMK+IjrKvFXqjQg00/eKSo3PnzbsnRgkZZ7dHiyO0cNfGS
nszIFQIXiZoFpjuUVRm76KwTyrlsAty7auEthXS0GSJgleK2suinW7cIvnsCYvqSRp9Y8QK/PR3o
FS42HUZM55jgsX3r6I6V76OEmkRkGeSXcDUyIAd0M2KkCF0KaRNynvByhlid+OOMH0raV0rH6dw+
ojYYrX3uYmlHaLlXYRRJ3mmWyLwwHp3VrRt+YEQG53wxCvcTdPB5FiVjuLuPJ7QLloWGz2U21JFd
yDMkDlLdm8dWqE+OvbJqyoh2ZV+L3ki+C5xgFXV5YLVYdEEMyqwcShdSxAkHWOWiTIhjowB42kaN
1ER4HADtc5AEpmgcWaJRgrWKZSaD3YpwEp0JU/TmbZTzHBPHM4FtzFzKMwfmK9BdHBkCr+8PqFt3
Q6tg3z2ji0IrZirWWtFwBOMLMwYjKkfyI4v6qwXoAaPuScEynE0M/ZKIFJxoOtgKlntMPQSkepvv
aFx6IOZGsV980QbgqbWwIvOa4jaVP+hdT9Jb7i8BR4Yc/0ex5eUkPuoa9yLteRMzC42Cc1WkaDJR
bIc8U8FLOCr/1jbQyAHg69H4ycJWJRlDkhDxMxw2E79yRJN1kiqBQorE0URv47ppknAuUTJomRuw
N6vuR76h2QrvIt7RZJFbzlmiPLzyp31YqyqY7Rc0ijIWiXu8xwrPB85nclpZ93DXy6YHcGPsGxs/
k8rnY9KOIJlq691+BDcjQc3oMwl0wJ+ZYBhsXEQsa3Cp1ZMV+uNDxWPCV5qnwOTPoG4D/rFyQ0ag
dTJOiB4zhjOzubY4PQSL+1SfjLxp81zLAnToVr2t8wrhMM/mASwTgoxgLioISIPSL6UBG1i4FPN3
5Xnd5TpsrtzMEqb8vBd7FOAYo6WeO+KRa9xXLxmn7oOWNJUBm9oCzYt62Lz0VrQ+5O8/RkWIcC6I
aMi1rh8G0jD9cVqlOLTfgVA53Mwiax3xEhyj2Y0oPxkVk7kLyiPVsk+u8+hbf4CmnE7HCT1DMO61
JZ3k2id2tZuGoGavujHPbgEVwD7IWumxpO9X8Wvxys6YqGZZzQAgpOg7N6TKZuqaAXW7sTz04/jG
3aN5pqxrJzp9ZjXaLtRBqC54D5wIj8nCmN8vnVl/eTqSX88b2+isbDhBh4Ibu8UCamDWAEQlQUpI
3hdW2KOMVoz25ZsYz7YxvzDpMZQHq6LFgcKDAyeA9lU0En9s827lYMMwKYXM9nn2y3TiC27INZam
VQbLS1ogeKtgFQSikIsh95yftAyWdT5JXxW8BdhvAFwT9Xnqh0ZOjPDLF04bKC+CzdZsTdfja4Ft
9Aski39sDZhbHTJg8WmqGvojPqOihZx9UKg9taR5GsDVv65n5QeRcS3X7/T8qR4YT2eCmgVQBaxG
ksXGGQEbnvZst4J74woVpw9pVWJ7YQeuT7vtRuZgkkYgwMD/nymK6jubb3ALldsJf25zM/6Ivpcp
N85lvgrdXDEVvniZPol+UtvNqph+PqT5Wxpo1jv5zgumWVlaWj6EakG0y8Rjx3FpMvLb1NXcaFuP
TXJDF01N7yRo3ky92aZHIkjpQbapjUiWcj6mAz+WSLjlw1e6yjr20SX/E8XRaMjDtTKaPmXIlF4L
Ce4wjsayNy1kgVh3+GAZjtuSyksJZr2drUINgH8qS8OV6GIIiT3uUBgAztkiSxM4vW2HM0nUIw8t
V4WNFTF0XRC1E92bZK7JS1CCAMUma9wXl2iINA3pYY43wTrpptZutcU5pry3plxnBmDlxUQD5xmj
9DIprGHvTeyRztUIxt7cQGSPpwByoCqaKj+kJB3ofV7VvaVxYicIUWM3Y6ebCHXeUyOEtXjlHwYg
OPON73nLOzllWwuYTneFjERp/wf/UgZfCTdtnthIhouT8yP+F1bivIOQaEBD3KtvkAWB6r9hYeI6
7ADlk1XLJdU76gcfyKcLRl1KC9dVDhvYM2M59DiE4o+AyRnWKAN0hvkCafmp25d1VcbYx5X2QZ88
fjqq2/hoSa/cbcK57Twg/6rC9di1OzD+7I97g743rVHYllJLPsDKB9V33LqjhvVimCd4LZvyGt/4
PnRYtxcH9ZnplL2UpfVAv3p4X33juCyXjZRw2LKIQ2n3LQqHCiuMZ0GoCwjFtv6w0j9EYv29tPnK
fHQ8qUfBRTRppouAURDfWpu19+ZcNAtHrbWuurKvxE5/2jhVVWzQnb8MM76m0xr5l6xe4AUSOPvt
NihI5z/hqsoP9UsalAG8U6p020L2H73Q1bX7p5hVE3+rLaBtMaGWDtzzS4PIrplVnIqcK7WOCDRG
aiqOeINitbFAuFMiFzuQOPG9uweEahSK29dzXLhb5iHZMmOxYMj3292m2Jfseu93Ol4bZKfSNnsZ
oq+7ErZUxKtsUUxTb6vcvAzwjI+XIE1v0/TwY/hTP53l13ybbN6Xjm7mI93/+RAYh1wvA4pg74Y3
IYaJFS1Og8zQC7PZYmy6Z41V62nl1HZoIp/zCTzPavF4AbHb8ymM+Lw+AUB+xsnCcRu78nfvUBHX
fcA8lgibegjYyNU6mNUBRT27OQ8z+vrzT4yncRPWiEoGTq/EPxnrGdW329XgJDDCibgMTR9MbpF2
Y3iNTku2yo1odrISv+8712Js2J1gGwPmoddJNZzCvnzKWYQGTHk0Bp1qD7Y3WoHwtncRvAPaYs7P
yV9KVFOcl2XXBsNMceF9p4Oeb7b+vNJhfQWR872cAaCytCGhDP4FU/2iljpgtJzYz9ZDL9pYAC64
RJNxMWDJQaFLBDDEhU7zqdqWgAxYP8KM3s59BL2AcuPI5/rRoxs/DQN1+icWb7VZnKmn6PyUnBc+
Qhy7b0YCYUoAAKKkF+1PB/6HxJf4okgmYM9hOm/XGUIwh4Hsn3eIC4Wzkf8UwtdedA3146QDg5my
lZUPSK6DFmUGOMcpHS+GJ8WU2ycXuCx0BsDt62okm1G7Zjv5DhyrH4vgkDSbB/NPEKylyK+3Tp/W
SUxXE253jHqQWnpctLpMsJ20oy3j5CigR3VRStsBBJ9wxo9N6/EC6tQWgkllCDp7wkblSBPig8sJ
h5Y5TWXxqpGB6aPwiaWNUDdesYWc3KqJtgrjnLp3Qcqx7lDvhWOIe3wWrbNOonKGuSsdaUZT4wvj
lcTAS1v1zecFAdzusAEnJV+CpPAlMAmDWJ/yT3yqByvwgnF1F6gd7DGbEKPM6NXx7R0lVM4YjMVb
7sL+Gv7MPboRJEhNh8zhqkENTnpKqhou34ku7YNVsrSQjIvn0eDYl71mk0Vvfs9hSMaaI0hctFV4
dij+oOdmDlW9HRh4BGA53AN3SnFKBRWPJWUwSdMEOvQwy4XOUs6ZY3+dwioZZPYN3i4f3AG96egz
Nv8zmjMc5RHTST+aIuPwLkExddc70JptxHyLU0VgqVD/jyAT3zwHRiNYT7yNTCw9ak7HmBSb4WHX
qDjOucqD8fqVWsPn0pxHaJ7Mm5xCjon32088/nIEEdR2uKL42X0OoyUPOhdQ8QzZTFzFLn18nE+V
45lgQ8xWAEsL2GEGYZvnntV40KisnbTxBzsiWhbo3R7+NHjIEL93puGzoCMP46qiXBS5NUGGjzP7
Oel7ImIqYA5KkKQP+6Ce+xb17OjkdDIKexkQ7LSzNhMwzayZhLjOsv+bGjF8K9X4nJvH8zyYWANy
JIKfp4q5EHj6weTFEc/3jevGqFC65OEFqpuz+UeGn8idJuOKxL7AXt6i5clXA2sQT+rUuSdpH2IO
WLNKu5Y8Nj2phRKI6kv/wD0/EU3jJOiiC9go7NtOT4hGq1sngfcS39tA5Fi7gAwAUhoOo+CKlhI4
9EKHVRJvr8wriTAwdA3Gt6TxJrAXeH1tsvUYaQvWANdmJmu2SOy6aUPThaZySrHrCqdeTFzn0nKH
MFtZqHPHdjILkPTNBQtcfgT12QX0uVWWp1mWcXFWfBIrowdgU8DPDfK1nSvTHgkqHo2BET7RlBti
DvugPSLfbeOzp2cGIpGP1uMqaUqTrzV+4s79EgYLN+siflralHUvnFdIVuONOpq4YcXFyNiGD1Xu
AOuNbn31CEXY79T/xT6Eb4s35zhChhjSEs4LTrI6J2b2Eizo91I0xqEhhJC9nS2vF4jr5mp4z9nf
+c1c7vN6thxdcuWjQm2yfUfiza7xyCn2hloK+gzJy3CUqVqVH7FQDDs7NPFSm5n59Efq0t+R2bdF
KQUheUAJJtyK/JxWKO7VZQ95EkCidXwsdsZ5cih1A5b3VQx+C6nGpsgjST/NvlsYmVgONW4R3wtR
eh3dx4AimwwGANJB9SiSS1WjkonNj1i3iJ567zGTVa3ktJjGUEC1jeGpZDggMh6xh/qZgB6UZT+f
dqKS/3u9GDvSbfM80m3YLkoZTn/9j2fbH5+GZiQizY5fM/ZbqgjzEoECix4mJVDgkQ/9Gijs7k0l
caHX+hgr76zw6PErI/ftbOR/OfB4osPXPhOZpUqOwJzKxjzJEPFdjbPramg/q9BgummP0umsDYur
9OLq3Fvk2qmHGm1cEruepB289zG67UVz3PNF/RGrpQpN067AuPTMHbML9ibkn0i0RMKdbngltm7m
eie+iE+3PQe0ii7dNZfjARSsyKQm1wEiSM8j6/F+RkHylt7CkAPMk4vQguHGFiTHtlnN6BvBR81E
NePWKhzfn+IyWg+Pl8mTzA8sim1F0Od+uen/V9ZAx2n6mzj8CBQu/bAI7xMkG3UBWfDvWquXSnuI
VwmBbd+skhywRdJAfd1pnO2WDF/42HjKDZg3LJSZ7dGATM4KtAsOEE/GnyeGTlFemXcA5dYvkARi
t6YJrd+h9Z0OYoDlzbCN0EVVOoCB/J92yc9N/BNilU0WzD+a8n3NymA5vgRry2cp358hHn4aGFPs
aI/JIIsEhgm4SVkksT/VjTqvHi2NxDroBNGj8SbCLUSR+7xFm1gYeYgjIKlV9sWOdFMi/r6U6q1w
Nms/MJKz1c6qRh/ChODu4aOa4mzQxCB6mWve6pyt4+qFw170ofctDSfuBCZkNWFkJnDS0yFol1P6
8fWcQ3TDnlpPOM1J+XEgNYemgYb9AfIJeGmbh7pggDp/wzd4gtKuLpl/w/383Iex/jUTzetxEBr5
8SuBSoGDEY5VHZ5PUQVaoVDutexbvI6+fjXLPbqFuZONb7BrzHRhHzx1zKMEqvn4Bl0iI7ciA4ar
i6PnNKkyY0F5xhj8c9xIV4qNHrvGKKcIpn5Bv9w1gvIm9+edD32CdwGjB23R+vl9LWP0/I4PxV+z
/10n6fg0HR/AF8nxr/jlcnVD7b1/6NNcpQNte8nMnSmI2padtRRnoq9dUe1UGyxarpsoi2pVNTcw
T8DDCkyRybXnCGiSsQ9RgKqLhYSnrBr9cadbAgqoeu9KQht+2Jtti08lfee4hIkdMcm2ltdKug1/
ax1VnK/f2y2EPbTucbZOMZ2hwwkxXpJgM1klBlubV+dQeWvs6y9R8vjUt5eTu3oxUAlDwe5PJCga
kHcrRrMxdj+lX/Mlshxjzo61S3aVcPM8kPMBHXKe57x98TzIsIaD7VFpzJEkxfi10pp1yOBPJBnU
F5jnTAOpbDCM8c5H/f3EYKb4GbZOC0NFE0d1Yfu8KogcMjEsGOBriA2bvlmFdmEkBG9FpegDq6ue
HuPjeDXl7tXyKtPZ99tDARWPOpv3zccLlrqLUxzGQQgTCxnx3uTOi0OyR+R6eeLKTHH2DDmE9CzC
PKdvJMEidhqPCXsDfZBLvAF1FY9lL0x+qxapepCUv/jmGR3PRrBnVwWkhppWdq8jkz8L7eeSXXIv
eep8w0a2pi03hCbnSoVP06ssJZTP1OWVyGyqT//gQq+1M2GouhjCmdj4SPJqAOVtYIlLhMClV/iB
ledrHtWfpEX/clTOoM4QsUvsHpCyH/JO14CZ+pLd4B82bMDuuQekY/z1mSrie64OXp6nu8X2tSwg
EUuQ29Kq279/9FpgGrmbc5PSwoy+9YuDZwBPwEPVGBApfcg8EoeiJ11a725Hw4t/k7O81jyu3ixc
0QpFGWtZqionx41Vr9QwoAWZbIaSM2ncY5gZY2iFKx34zYHL6nkubXAk+QF/65yr6HTl9c4WiKHO
j9I9OVREacRsQrc/f5gVDGMSJHQ/z1gpNqFUADayyIhTXvcX9pMaHEJkY0k1HHpdHaUTXlK0QhO/
XZ3kzDq+/7HFLKSH54noqjSEP28mOKMyo1CT3u7WImve2QfJd9ptASycwwovK02bUfIt7vWf35qN
pOvW9u8AldANXpbH40b2O2CtGdaf5ICEnXcpNGmP+ABRIRquG7oFd68/f2lb8rIiyyNn6JMcMyix
KYxCbmXl8D4oo0gPzTNccdI95GZ7v4M4hovXZGVgb51ITcJoCVtmLIw/khXQiW5rbERVz4J9jv0a
2blcVKHeWiGOpbR/ibO16AWHeYu/UcWKprr0vGeh5vM/3/1mHRVxjMlcIn/jt14UK6IRh9JREiyW
mWtaKO/RnndQv8+QIt4FgFxEBgWto8Su6tmeP0mbAm49AylgEyTLXMk2V1gNPMs+/kU8pFhzcL1g
5tLRYBVLAPWrn97mjBAhPOXl36keC1nWizgpjZikW2/atjMFNmPdRBdymjv8LgiYAt0zGgvHPxi9
vlkBUERblhwR1nhGFViQrxr4LqvYuGJrQGIDDETqSUakdyXIqp1K1jKCJHU64HeY8qafN8vypBFL
OssC98eF73hOC9yKOwcSULpJhkEHEAK0mq10XGfDZgLQOO3txM2rLlpsaeGzLTaKp+RcFj25YBn7
8vqElejiNlTnY9O2YaPGFw6Ei+Hz8OeJIbBcLolqWKGLw7o1yuNbVjzAc3CLqCJV/owtMVi6EWRZ
lhNrwUJSGjN57UT9dak8T46a+PlKmjdqPEcWCIwCKWAHsILzD92s+SOOekBhnTJT7nQWcSVDis4c
7WblZSmASczDpcZFgFRozpJQd/hoDoX3chg2QUGx3lSSJL7bi3OqKi54GjPAQEWm/Rsa2kxl92IH
oQABIh0Xzd7ijeQ567ZHSL6NoTofcxzhQMDfx8ayGxaJnk2JwKSOiCutp3ApA1u+QgADBLFN6YdP
ghDTt3JQ79fSnViaMENO6JE0ORYl0cygsnX7PCcKNXPg1xJqZGUj1bsQjDeqqMZn1vUQAQoyGN1B
9wBRtcYJkdYi5nNAyzgyc6AWlyjK+Hl2uSB7Z3p7a/CdYWU01bOxEBbYQR5lDUm1T4OERrvnaZiE
M77Ni4/0W9IrnxBJyfGT7CJZCgMP0HgqA8CjFg8kS6B2A/LMFFcx0yT+lsE1y4ZInvkskWcK0ZE7
bGZ4k+gNcSCWoVrUbLxxgxItF6cPTaUjpCIia0FI2fLP7QnkkKIoRm5ZLet9OgqUQwRa5ftRaBPb
c0U0JZw8N5RElFV5WjEln2cNTfLnrdmS0OVI9Lspd+avppBJ/MEvTiI3MGEN104v5jQBaH06vhBj
ydbfPmkJnj60+cPjdW6nOdLcoKEHjJKc/qkO8GRfEJ2Ddew9xQPh+W3BbMP1rGtFd+GfJxrECjUp
7c1tcrShJ4U51wtpW1vILdcUneqzYZ+CKd9zwBp9YCWJP8qWFn225KXa2tIxAh/HxCB8JZPflYvD
2d4IjCQaij+BlXB+kv8ZF7oRGC4bzH9b8yaJmeVN/leUoxc9Iq5SUGpdvnDl68nl9E5snHr29Af2
0ybk9d/u4H9ltvQj6UxI2MveQTUH8FYHPJys4RJDiSGmVow4P+6rhXOER9Ibs5L3dtNS1FCq+2pH
ezn3nTLgapdscpnenmaPeASzx9ejbCH4j+wNoqn6mUlnLmbpHI+rIPTurmPsov08GQxL95vvBDeY
i7ovzOklissBqIXokDp1ARY7QoeKUFFppPvsEc4bTBpLtId/DmXKZEdiS0EpZxoRZCNeRWA7vUAw
7LZfFw0NijYHMNccQ239zumlUxd5XnyV3YQRNeXwpfQ1bB8Fr741XCEZXvKuzxXl68QuhPV9Cq5m
R8n/oW92JSwtx790Rj9Pxn9VSUOwDW0jsLMcT4zmUv0020czUOn1BBov/PPnd3ejlbeno+TP08r8
glYgHpLv7EyJ2WNQK6t31QIKTO2vtMK21FG/9jtJUbdQy2HQAaNH7ASTzVeGzETeoTdU1CDKJUMn
+zFnH8MqhLtPx755lQ4m/1D8HCpEhTDSupZ2QWki3Q6P6gogXzrhOrDfKP+vHS90K/SxJJ6iKar3
4iP4ibZr5Huzwdw+ryBUfXHG9IVdjU5DQL9PiK62zeTez390BvN6P2Vtz/L6KKPxYUvA5e3rbJJ1
nKX3tvF1m0nzjEq98I8sjedTPo3JrxCj/92vXhNK8VdZN9m53pGCpe18b93AElhPpCxooX2EPl4g
dfRC2VP5lUgVX1/0oRL1jpEKRvt/NsiHx9ARLFC9LgPM44OG7fEZzGWliNhJ6Es6EQxVeInUd2NV
dOo7kjjZsH3PrNgEj/QMJso0Ctw6a00b1FFOzQlq3K2X6Jlh6oxf8t34Oso5pxad9Mt2NHzyjWMo
uUA4wo7mxxgAuhRykektzfTZu8tYJ0il0OUm5FG0JMu4PlqfwTxpveqB5iOcW/71z7mmP7BWECGl
wFETtVfhGZ8eXJ7NZzoi2hTo29dncqVl0PVCFLVU/yiLqvX5PAwl8B2L2cEXXGD4FStbRLGkqejc
GdraFMFWLOP0iZEHRQIAIKiwRCXrO0OC7kPyIXju+pCsAm3wOkszTflvzWg7C1gDG97Ifi84I51D
GS1u584xeGMfZBKCPXcsmnkVtOR1pksj6C3CbInwlYkQAVB0EVCQSgQYf+kD/ZjuH4TZyrVNVCEg
3oLgUBfF+viPHzWHsn7UlsH5gFV5VoMwC2xUgzx89UUNA7+1FO//3ptltZoGGnJtpMzAyV5ok6ah
IMFrePsOxcLM/RyR3r3ttIBIIyj8B5n+/knkZvCTpmPBZsimutn8UiiGNmpPlmUxxhYguVOB/JPx
ZrGEVvY4V29VdjAm0r83VmbqeAnLOhZ9Ve+kIamYPM6w701Wo8LJgWr9rxt/9KcPaCx/HqcZFHjX
X+9esiwNv4g/CNPCsnA8sPrpXfh4Kwiv2YtxBW6x87kr36Yg22JA8F50Y8f28B35qXVO55tOE8oW
uAOKYGI217uaNVbnNXXk//pZAbKEY7fBn9aBYj1g0BLi54VmTEaO7GHUfLbxAi6VzwZ1eGOHm9w6
ZAI8Iq5+Ef9AQ0N95dKQNAJsij7pY9/SS3HFQ5KdZpaRr1wWhVl7/R4klrYDkIYiICIla9wGAbOj
kd+fsZ49LQMG05nrDWytJ4/7zoaVey2m4oB74bsE8vSjsJljMBr0Ae5OlWv5muIUycKQqS8bDPCJ
TUFvb/ntTXpx336fPSR3+xQ+V1VCw5GNNTjRYN+rKg2AqncmEvwkC6Ybhl30xfA7Bwb1VFVDNUVw
ORBj0cTo4pAueOteEQkupqWFHX7nNFOpFT1ZO+SbiBruEvPL2Ahd0RZ5C2KsHarkPdYQ2cqvGm58
/v/546foxlk2Xn7RFnTJFK2WE5NTr0nKg2qr8qJuPeRQgG6VjEgSTBKziKj4lCwdZnJxMl70tZO1
DaIuGkEgo6FS7L+osqIFvwhV+LnW6wj9bh8dGr81MtYKWv/1TOlWIMwNA4UH3ooCBACNOiRgJeRA
YwipZJuw3q5aQ+viZJt6FRKkZSLPN2H63C/8NuhqYU8P4tbnP1PO/cB3LJ/QaCzx1/RRAUkVnuzb
NHZ5nn4Tk8rejDcA6H49Jfc1jzyiSdc4hMkPiznib/fJQW8tv31XWhAwcN8IXv369sAbrCxZs874
bvTQdK212U4Aoo33T0XZijJ0XPbX+erbZ5y1dVYXXBdptmxEW4BrKT43sEQS7cojc0qJsRIpkPkQ
C5JkVNbO4kqFUI3ymawEP6QuBU6HPYWjU/WyrIGl1UEJvtFFKZs6+v94KCuLjH2gBQdnGWXLCVr7
DUj2UL7a9LMpwD7HsmfWmw4hVZw1b6VF1okxUjt1qoKkHa6yVWUiKozwiHHrCV2ZcFl2a4ncImT0
dQvRrkZjNXQnJPW5IAfFtFYLn9R3jyT/PmrPHU+H8/VFDwI87NZhyoWzvrbT1xVxNl9wXfbAvIMQ
XlzCaUjsKdMXDQfS6QkeJYHkl3IlYr/LnevILXW7C41L8oiwzojEsyd5SPSlx7Dzjhv/ANHbw6Tw
ruDj90RaeG3xLB2qSMCKtWcSR2Qw5CxznEO5IlcOrySaoE5iKqFbZps0UGyHOiIzTgO4l81uNtFW
Yy/7XUlxptnK5mHVI6iPYT0a/2bUHKwuh1rPj79I/QzRpdFcgiyeUVOu/qLdCxs3d+Qca7fRV2Qh
7q7iCwgEhmt2/ZPCCjmwZxom8NoYXnxWZpe9NffzdK3lQWZpH6hJOmg/6BpeVn2iooxPMMoHsqvU
38n9DVWbH3/mnbfXwIotxaYVJMmZhVDH3koLHPUGgRZIUuJUxFRtjRuLJ3DUoRapFkBZMdNBmKL2
Gt/eVSMqdrv7Kq2mBee1vfw1rScUKhv8Afgb8rFglWffvwITwYuigxuEgg0NawwunisCRp5e+PC9
QEtebQM02UDcWolwpnjC77OlsJEGMh32yhIakpEKJ0Lqt477myZ4v/uu/jqPfjdDb4sGopGbBsTh
iklXOiDLAy6rE4jjA1vRcw16H1QwoahZaz6PSOdGMeIgHc56n2ASY2r3bHMvVMkb8HWAtsIAR1iY
37IAbuohJ2J4sLZk21GDL+C8HcfwxtMtfRzWyqrlZx5e9n7TaDXS+BcwVIH7g5oWmMc87vX3F6nW
L1k5LFW/HaDNaX/bjzmH9S5EZiX/pCuiK/YKkzWu964RgardBqRCYahIUavoUEkeGo4sKIBo7YEU
OUfyvOi1hfKBxyoxAGr8c35MQgI3mxh8fFhBL2fUrJBpQXoZWD5Z7oRWi3X7K1SXvKoCpX0H2uaB
s07wAtgWt/NSoCP9fKJn7H6NZ1wqrGqRFkM76nkaPqxCWTTp9ctlPyV90gi9JOePRVWwvYdhN1Mf
kB3IleeJx/hTnDnV8Se9RTkgUbY4+sKVSiERxePXYYN7Pi3s2hLyhv+uEJUxKyue2QPfHQO3s9R+
FZz0YNrsTTKkBJS1VhM3M72FEfZMX/kfGR0poYI1w/reogRN2vMUTlJxqHEEEmXS9dBWdBTa7YkJ
a7FLFh2uBLHYFit671NAj6LJvaizFRM7oBqdW4R2Za0pyoD6bOMt+Jz3yN9WiTKnFz+ytgn47H1R
W/t/7n5VsHPtpECLYjeY0simH82h4xuaxL98qa6ElD9h/0NynnCX+r9KaOKLxAS9DIWsVXzbxwcw
5lLeu9XX/nWxned9hnwyHju44T2xZi/jNS1+E+CPFbpgCoNjYLh+7hppsxc9G2F8POUUsL6/W+Um
4lUkMyj0bEG/4Wwo+i7EBu2gekwnr2Lws104pXP1quYF0NJ3BkpU55yxLYEN/qwmLfIcNVX1ObAA
6ewy9/+t0PV9EPN/KSXRVKfpLpjr8W9Ezp0OvyF98O228/DwAjQBUJMwptXlMGVVkSgqDxZXb69D
B3QFdGe7LLkJ4uRU/Sx6Imb02w4uaU9IT0TCPxLIUWYl1VsYIoOln19qsXBxMw93vBkFwvNZBqju
1QP7YuWy+727iI2VLCRP0Y3k7pSU9qb6Kj/iUwcp0QX+dfX2aGweeRV2XYi8OL3C8ZnkJLrf5w12
6JIdy8YUfyx7cZXopbj7nGSZDRdpLJ2lgHjonI4CnX0H7+BvLQ6qUd8DGANpjwDKuce6ItanoWp7
2sMT0H3BJJxt+wKFr2cPS24cqoc0HnrLCiaTtAclSgNLhymMVZrKEf+oih06H8o6LOZxokVvQkqm
Q807/c9DGy6AJBHQlFNK8EnP2LWLw7yKvNSw7T/yjQHFYtUPRHteSw0nHveq3JZONoYtsHON8mr0
veK9M4WGF66/yaznfJsaQ9njvc/NsuPWEHshneNRzJH19Wq6gLuvzI33rQWCpmBHkWytayj57lAB
gn9i92ftbDi/YN9NKxOIuxETcoQBaQ6pR4toikbt4VWU6Vtg9vjFhnhGnY9e36/tC9/lzMz5latG
MeyIrw+12U098K6vOvTKALDj3xnM4C/NGkuoF43n3W2tfXXovp5EpnDq2vIlOt9V7v1dbJ6RP1Ye
fBU1vNsOcxogr53s8hrFzqKk0ZYbXzYFyx10EPUkFVlDBsz6NvFO18580vrHfjUhDfNtNbzULyDT
KvdgoDXd8z80h7nXITAyejibOznsXnGhvTTskv0tl3Som/tHPTJMoMwJcH9I5qHGUun+46+Kmpm3
eX2YNgryHVNqkGoyyA5FU2wGqOrK7c+5UlX9gcTgIYb3LS1+tJRSEW5Yf65z6gSE0RKUdPpz8S8w
DIcUyJjfGPpz3Rgx3KaOTangQwMw7aPudYxiDuS4cvs8SdURmiZHd96iDcsZI1bZL8qGWBWaTwt7
quo0/k0dfIjNTygVOrwp/JEtHyB1R+eVmzKS/z8gUiYu72JF0cOqh18DbtE0mJ/pXC6wGBDvBwaB
J/DqWxk/EF888QsjD2e2SmyP+vXkivNOV6uo1AHIsHjk/odYOfDWkuHYNDPuUpgMreqz2D8iDcQ2
D65rg2eWeKhm44vQM+3k8HbbXtHTgsIC3OltQ0v1IZ8ec05AjPyiKCPAZt4eN0WbOC9WmVYxgchY
KYP2J3GItVf5Px4yCLMDOl+gTV+m/xie6LTSf+xpxfDAk24+U2JLOGcjhOnTSS5z/eT2Tx+CvETv
D0n0ZAhi5PhGsSfc53C9yJodrRn03wJnp6Z8O9DDuH/xUs6Y0n6YAqKN9ZiTpDnXR5n77Jpmb9YT
acCDV94QuQpgsoqvYrxTCVqw11SgM55PF/c4N5wF3QgicRSAlkYXBwj4rJLGx59WC9hRmID8tqV+
XAoHegJCDCxkhwhuzDwLujJacnCf/C43kzmev1Evyy777GSepDF26hrVQ93Jf/xM1AQFND/sIPD4
Np+l5pmI5l7kJTOONNGa4S+namxwZNqvd+Dmpiy7wuhGoBGSLEPRy1wqqDeClJTqxxkANKgx8YDu
giqiefQt29r7gPPbxnb6folCmqAernbvRE5Nhu9aXX2HjogRD5NdjqLdtygVfdaS6EPK1y9gUydS
rFueSf0FpnZ8Vpynaf/wdgzf3x5+Qb619YAfD08JCb1Y/Q0l9fTn46flT+N7B04D/UeO9T8J6LLD
Ppal4QS/28Sp8s3FNI6/xZ1a5fwDInXvjVW5DNZNGeomsmwFdHeOWU1t7D2jM6LnXJnULaIH4pnP
Huog+Vy/NCalw69jQDDTx1XmqmidXl5pvjstWYm1XlZngMaYwtXtAXCaEXhquSplZU/MRqItZWr3
YjoZWqZm1Rf/qkPItgXjjR/AWkeKnj8lzX/nt35emIrDd+ogBHzPOWRwwI5pJbM1GEhohzNA8p96
5pDHWJdeY2Tkr1xNeX69qc/6Vl2gZRX0VwalVXAEOAfSArxNerDFz5w3CLdKAfROquCwxnuTp/ZB
3PHFMTT2DknqaMprngqxFO6obFgapyCEYwGmNlHiJgQarmv0qHpAhrGKNw/kQBY/Dt6pCLoTxKCL
1SJWawyvtJ3HWGVSAZFmhzC78jpQrlUeYanRnZpTRIZCsUNMYBJob8CQOi7HiOxQTOqVZAsmazzk
eFjiZO0VQzNmsbtMqTgzFcIX3MTsLBKF0TMHZH5l1v3/xbsGoka43Xmr2P6OgeQXtwKcWwHzAUnb
JHVRL/PmK8ocKT7FJU2Kjwtk+M+0N0cy/REPib5Fc0wLq69Avg7zH6kn347ny1KCgCZFMJ9Wrd9z
qlFDOm4hO1H3wofEe4Hl0ztf8lCVykT59K/MgdC/nhp/n5aNnIreTgybJK4W+ZhAsDkFDqNQrIc6
nkDDzbo6TWrEn6Z6KKlKlYAZd/tTHJhIYhsTdYFyUU1HU8mTwP+UIWH18mmGscrPCXJP+lxhc/KK
7eUNY64a2xQhqIZV/x1czZNR/3Zj6+oPhQwOY69mF27gEjtGtmydYdDgwtZtgeTguwTBO15H6Iwy
w3r+hJbuQaN4LP7a/FuET7xLdisbFEP94KjfyGEKrTy4f7pTB0ISid8kVcK08jXVzh7W/EHgkpjU
Pke2XmPDMVsdU/rknlsVdFBfHzK3h7XaOEBZWTMD9UBm49TzqlhyYj635sx6WnGpz258bIxw2b6e
r1lKg2Rz7C0hlJdDn55/VviAi3BQ8GBFJ3hV9guEuM+TnIIxk3VOhwcQKSLSJ5JRBctnet6j5MKq
nHCxabXrpM/N7rEsB+yd28A4B3ox7O/OSp8VFBXD84xu4ZK5OCOGjBuf8Tcq2PhdIy4/MZBbAQir
39Oq/sxnMW/vqkEP3dpl6I2KMH0hiY5ElQOB3Wl9bqbcmvj2OAZPGii6+KswWs4M8FhiQDYboLhP
mGwk0DGv9u7ki97a1kwIVRYxunvz3rSH4Yau0zJkB9xcdkvFsVQ3dISCldDsypKxUicegDNMZe65
HnPE+o0sohO5PMZg7tyxHx90eJSfWT5o1K33BAyPDa1Vv+gfpIZanIgDSWmihvzylNz9qZXBbknK
ccpaKsN7321ZTl7ltZZEYZCT1HHi5HHCQxHp6mNvPYE0+gQ/4rnOH1Frp+cYegYzPYKwAh365vnR
iWKF0HULtkoYaWbDforWf6LlmN/dIVBaGSLEJHK1YGJbAp3ugYv25S54Msa8uq9b9iSPV8ZNFeWO
HUW7l+EMiiYAJ095F0XJ5j3OcZCweImx9Afha7068pH4maE+//yKF3caP72JmUbW+OhFeodpYOgq
ffg79TQD6UjVwa9/tJX7W+Zp8VxDwmEXFZ490lY7m6CwZt7hJfWHOfmup983XTPnqaI6mndRxjvd
owih23p7rRe21YV9pn4eQWIG5EMmKgnYoPY29twDeWR4AuM2u4DHzqXiNvPJkBIJ4itz/+xHsm1H
2slQ10NjQWQ1JE7b2hmnEcynIQWAicNQgqTJREhWBm1nvkHBeonzyxazTZfK/XOVXgcuYQoYc/oS
+x9JQPHu8R0kpNrWTW04Zv7YLbdVI2HXFL33LGohqidMCLH5Wxa5vAUmQfiXc70hS3QhdoVfT1jW
UoxhNljDiap2QFrT522FB2mNtAPoIWF/OJSEjn/Dv65RDKiH4zHPLdlxAqegbEwX2s9pWPRCM0TY
NyNtWUBMCchUaYUGRgzDbxrY+uAJp1mCBXMaJJsF7S02c0HSuYFCQw0ZxoQJtJDgQvPsdfDEFp14
OMAZPSbR0UGV4/0DZ+xbJP1n5b9QBQGqe/xa6hPBm+zKI18x2LaoT+z0idRqppVrCbVAOQocVXkG
1SUCzBIqGy3+uQWMqQbkinrwyrc9Pd14zsWitn76fCPRWxSwSayRsk40npmS+C03+oMnM1ZxMjKT
7FYpsJNFhO/cPU30TFotAdM+M880rF0toTx8ZohcNyGGLYs74GgiX7rXI2WQyf66ocUrAEbC+vbZ
kyprp88mPxc82DVuUKtPor/WXklN0ibwg4dtYzVu1SsSPLhI9Os+ptGX6ut2LndGLta251LxlhiM
noAd2Tgsi0Wh3Y9YevJ8jYt3paF5/cG1QNK+7ySAQpSda585+u61o/k6S6/H0w09spRn72lDWGDX
L1GCQ7skOJykFFcPmVIXg5ZV6j/v7XaMZHfL9sjHs8qhSOL6JwVn9P/jtFfEEwVeS95oqF/XUpGW
pV23Ve0UNLb2GFa2Ryv/Xuw3DjBw5mu5XRqkRRx0UVzrCrRfuqTTjCIB8Jse8XB4Wi3Id6vv2T1Y
4eIb85zWyfqp0idJde20d49dCQDa29VLomQ8luvTwjI6S9Qpjx61QR8cD8NG96XZC9NZSqKB7SIO
9tVFyMqs/0syQ3gxVzW1dOrlmrTF0e5XfDDLkFAxf3HhKJehlCAhvos5zpSG5mT+RfV2VS+0AYSm
+EAZ70Szq2uX5vxU+PNPYZHZHEl2FM6wZIGi2VpCf9NFAWGQzomcoxEAEqW3nd4nA0GDB3EgRJUg
juCZxr2LhFTC+PvhTJwH/DhxLzvSqwBWMJVfcUrD3gQeIrlbY0BV7OhVJe92IjVJ1rYqbo64rTle
CBMcFSZYfz51wJ5U2hS07IbRpvn/ELeuZlfKnbRcbgqZnWb5UqriSDceP3Tx4P6pM7Zo7Naz9fPI
fko18wfC+8VI8Kvifu5pF6D8nM6VjTRhd3HOyEGwOIhiWnfAA7tdJYblzjB6NH7aqrHBBdDsyxKX
k8TIhfHaMeCkbt174I8x3mQWkW/bhqIGe3OmzX7LT98eJlJ5KeRZgYVMb2KbnT2Fd2R18HLU8mmu
E45DRKSMcenjdXmkl7d6zHW9yciD84Qkvd8ZMZUb3Cx4Vw8Knniua9O2XsuDRrgK+lcjpF/dqXRu
xNFfUsfy+D4mxHJYCjF1tRI8eYUHT5VOd53wE99qbbqmG5e+m6d/aXlHDWpPjGi2FhTSbo+EDq1u
+zlepcCk4s0Sh42pczaphGq7WE7m6IAwW4FIjuiB+ILt6wOLdk75UnU01yq1cb1KBzCmGA9w6eyr
O41FSISusvA2JXPLjfi8XWidfemD1PNhKMQ1n/JtH86gBTe2uZvmkyXv9REvySYmxla6K5Nx+QtO
kwusvQbIh6yk0FubsfGnKTdORGf+X/PgE9k+OTDysMKAoAltbXCFcwzuxWJqE9EKAO7HL5IjYH9o
0+wjUzt/dk8sn6FRvj6lrqlBsOzcTX4BdMK6GPU10nZI/Ct4SxGsfAPve8kJi1qwTAuC5RIEp3+m
uue+hiAAYMgf3fo8CfLfT9PRACmWQWZHbXoY2w6Q+yA4owUF22QGNMOU0GAMrqz8u08rVrSTVoTw
0htDcMu8FpuUkP0ycAlXue483W8v8dvkcFrAX4WA7bHPQJ1nF7Pqcg6Y7TQp2sdoe5J0W/34WC2U
ttxGJpPHClE5NG86ZPfyxHk7/xFHTBESfxer6M+ymHbrnAqEjkJpmJ/V26D1NUW5oamSfXvOnNtB
ubmXbYMehXkD/+7UUoYFSADgH5ml2mloZ9YxKQRVt4RkASBozJP6y7UrsbZh5CVBSIVLrp1+9hb0
ilg/XSkg3ZQvIRQNlOWu/NGe6GI2is0s2wdtlA9NFt7+51Qij/uN64iaU8dgX9xHWs0UdQR945o/
0JkQ2aKK7awIzF08gx2LLflvOKtRDOv5ULGimpItMF0dR83CkIen6MhiLCsrYKPVKuncK75xj20a
+GhmRy7ipKPRRCfKUzVOJrxBmwzuJzN96iZPny5goHmgK5WLz0HEssDf/hMHNEsbnp9xgN9LCaD0
mt8wDpm+ta43Pf0/oxk9B8QIVk8KSiolhqDaYp0o2YV4RZJcT88nOc0TQ/cEjDUUNZ1rTFd5ORz4
XmmO6FmEzWsxMEuxgClM6K0m1kbPxjpq83zQ6Bcb4e6hKEUIegXugmGPCsd0naw4ogwKQwVWdNzH
Hj1l8J4/axrfuJ9gQDbKozi4/LCe3DpqVtwWuYwFu9QIyY4s3/BSfTQLHw7TEDyOWo5qgeVdYzj1
sBSsWD44d6uT8RWSK+RxB1NBGKIIweb+3POlaqUCgpVN2ITs+ZSUbb/tfSV7COOCHqhWW7ngb6Hx
krVhvDE6HA3i5+6jT4yEa0I4drkJ+XCO2c/K9GQYLwZVjc7+EoRyWRk/ba8GRouyyrVocYzX1/MZ
dZcyGdmtQmNo7BZdG+9dz/jUWdxEhLRSot6k9Xkd6TW/6SpQk26loCbTJK+s1H8/E7XUnMgtcndV
hno8u2LtQ98HuPAF4cWfivXys4OzudB1elhJu+7wTktRIO4FTO1FZ7Lqor7tq22XdLhFdpJJJhS3
KcHwdKjfFkR4n+68C1rn91QhRoLpqC30JfkWCK9S5tedfq/bxpvXhFU+F8o4q4i07yNBRdXBTkMW
pCNeFcPiNt89Vp0KMBIGXGYlC0JQeIkgyrMd9w7ufLV5q4T39h9QVm841T8fJBUxMUsuaQi1H3yl
hTY0MFlz8nKAL6p2sJaElpFJYR4kzpzq4Qmam5OXylwDbLntugUGXCTuzGN+3+xTXCtAOgPviDJC
YPNtZAJJXsXqCWjlfrS0cWh4vMnO/iXL6qIh71m+rffmXUsp8s79RCeFATL6mi6OP92gzOxdO1sz
+XNKVMT9mUUjBY8PjyDuuwKFxrepcIiQg7FOwdPXoP0NDNUszvCXKELp9akGN1R7pRglbyQolLOf
0KW0oqkYviVIgL+gpv5gZBMWMI5NUb6fK2Ar6QbT+AfjR8TWf4RgbQyOLBEla9M47MKtStiVyaLL
mo4KvCTOD/A65JqxtTqAGTZxtCPVrcRnV6sEd/7vqa40TgW7chSvhuAY7FvoZ8YHL5PpF0PJasEO
+Tp6MIh5zKVjgq+S5Ehcqf8tnQoA2e2vj1ICuMdbnVYsFY5gek/c3j8gjTSl6ndgoT1Ps3fW/3+k
6cq4pQDkTOq2h1OH85Gzuj4W+u0FYh+nrWlMP9jn4Gb5vaBjU7JaZhqoEVH/lLuxghshN5gzJATl
xFcTegZWMhF/LwEEMdg9xlg8kuOQUIjKq7+udc3htvz+0XLYVviMwllzje2F/ch4CvXtE3+YsQ/U
g0phxLgqqSdhO62u8TvKVzbdmdU3fl8ga0CjdP7nl62y1xyOBhhq85Ml+7oz7C1dhLyxHFPJVPQI
JerkSqiqxFfzGP+xReRCMcTG1ZOVbmkuCaaeV1z8ddJnxsaN8iQgh0iVs3nyL90G2cT9dYR4/fWN
P77ZJ/S8Z0c8kQC0a8AMcZJ5jdAk1/JcycL/LlhM4/1KIxsJpEXGCnHSG0FgRNMgl2QOfvnS/X6h
UcLmMet7/5DLlzLFhdW3KZSg+tzIwdQH26pWenJkUgekOOqZZ5pvUiWpo9BurwTJm1griuEwI13L
s8SvdvV0yejZhINp4N1hUJhplNQ51RGBpr1Mldd0Tz0pcDWi29fA1WD9lC5d0gRCrSJPvZxXwNNW
MtHFRe76oULi0g9pZwfmFAOqmujEabq3A3553u+xUjQ+L+XwG3Ie33hvUzYeRqvOIzSrqNdcKvMI
9qVYaJKdFJU57L/+UztTY5j+4lTUy+knoUzSq8fH81n5JtbnTXWlwTOB8evbvsMml8rehWEXvvwR
WQUDxzgJ+qKD2WIoZq63ndIRH2UhXOKMe/p8uWsrsNez7sBgw+uz/85s4WIl6bgYfvOMwUIeCboV
HJmjmPM2NmAj00Dtt+xyxxNWsVIPZ3pyMryOOUSZtbmoSdUGrEPaMqZf+eA3hqHfDTqwhLRpbydS
4RC9GmrlnRzePgghIlzZRKq793IbwpK9mawt9VaJ3ZfHTTFG73YnzRPlBBLVfc3ipBGPXMmGLgWN
uPFeAhMc5So+ea7mXNb9cV4yIdU9HWve0bKtFP1BR6dKvoM+PN/+UHRXfBYQaVHFFUOIr55uAcrH
O3rjMrkdi/Yum28Ofpye72q4FErY0w/Qgh3FNh/v6vygZhuM2Xh549AI/8nn9EmDyAG1spJtE7Oh
+sYKD3uGfTAuXuKUF1DKPhVpv+8JsGbIidKCCwALwkSt/k+agdEQQMOJGD6CHtNLtyFcFTm9FA7R
zo97+ifyaj+fTinHZwpPtBqTkpX6cC3VDbWA0wKUX4soWZBmI5vCwXb6oKc5346t+b7gXSWqrbAc
MVJbuZHemqrDQxO1V1dL4LlWVu0/0KjPPxmHNmLCOO8u0kJ5bLKw5LaIRVJINuWLKA79ezoOi94u
nElAehD+92RWixfDh5hJAif1+IG8nKKDyFaJZjDPE/nUYsMa8RfzPBwV+zsACdfIvcHtX9Sff36P
0fYvpAO8e0J7d1QbKNEOMGnNneK+D/HlRz+hxblFKbI9xZEb/Im/pePOcmuse87Xbyl3EUsYXOO2
a2hsiysgeq2Fw5RlybGXGxYWDusvW5O6Rv1CeOzrxC7EoGEQvZ48XjELWwOagZh/Wv6fPx0kc9E1
h51HS6By4NglE7It0sT1Y+6orc6Y3aqdDAphDqAgYbWM9R92e/dmlEfwK2FRoguSfDD/7PCrabeV
iztmxEKLCVVmEEnagLlLNwr7iWt6DCf0P4bQwjCsHNqAwIDuTT7xd8eU+xP5Y4qQzHNoCWZ4cL6y
V6WnaaqVNRqlailgSepT30NMvOECkxgAfIR59Fkt9WgjyjshI3pjEomlC1LHBWmS7KdzI5jLE7ir
uqCOxz+8y67B5+arqFltQ3ld2T9JY8fQbTSGXhaQNIaMNkhS9jPdlaeIrPmQTQSrLLH0GXEM9tSR
imbpqSlb7cxNLSyCAQJNeGubyYwboZQqPdI1n0e1lqMjLyyBInAnUYlkxPkml3wfAUoEuFuZNDIR
EByjhu/ILodgRkeL1G0iVDA8VL9ck2UcpwQ9bajID0jI9YZJ17ypVO1HWom8lBhLtXcuDGZHeHOh
RGJSshsIlNXUYAQ3DkclVYuMTOHE3hNp2IGf3UWvgF9Rdown9ZF0Gxw8QRQYPDdCMDm4lfBf67dv
jjVOEtko9WDfEU66zBKXXfpGCoauYIX1+NLklIoLXgyRIlF8Z9Upw7abAqsOG0/tf1rSIRbGggUB
wAkfAcaiRlH6qxb+9j8nbUY+gWGVpcnSlm8osrZc2Sz+CPBVW/ymNj+wNnTbpJK173F2gMqghwAU
oLziKk5LW8F3cgA6jbfrtFg1ymqFMI4miTdWttaflSV40fJfrjHEVx+KItmcrPxeF3YpBjbYDVjk
7IkFzfXsEea5ucPoiLzsPNHVUROleo8Y8UQ+6edPf/C0JMCi0T/NoPscB742+1AVRUMyCNZkGvPc
wd++An+ZG2/rmObBKoFx51PtgpObzev3ivMKZrCdM0gwmPoLRQqjTuh/NStFUGSjIxJ9VM9xzlw7
pnJbJr10YBi9mDdhkZGRVF1Koh5ciHctQRIAhj3g3uS0I/QW9ZTYCND6Nq9auWCf4YkRF3bGy22i
xO9HYvkB21Y00pqA8ikf/qODFBq4mxXRKdiPjN5Cq9YcVPvys89+O46OUKVj8O8DuhLImRR/CJQ8
hFlFmhnabdaQu1hjPM7AGGmX1AwBx08P8kBHGYWhNSN+MvAhiW48YzYR/WxvBydN+RiDx2y6X+vg
0FGhS9MtKgI1A5dCyRRStMxofZePFIvxxExTiGcVcVgNbBlzXDhqp3+xycwUsD6oImmHx8neG/lH
CHaCFRRRsHR+BELbZpP/MNMzSaQFjn/QcnU6M8ko77ENpjvlu/Nleb50FFlPh15N1FSbPjHGBWWY
C/Jk0DoGLEXlp4ksWscXBn/f0A3xL82THOLl55O2s6s28jk+RV5e2ZXR+1RUZwAxOTjIqev0J7mn
5jNu+PzXJVHR/i9nglTUlsT4qjpbkKNIDnVWv9Tev///b7mUSXMBWp5+oBX49M789Oyhek9XnZfr
Fdi2qTcxpWxAql6gLbpuwH0AYZry0rCvepgwTbz3JI0kfztAyyBudShWd120fmrf9XjKYGpZNcN9
oxMPzEQAlStiQ7jeKxmBkcYrPKsWJ0M17na3cC7tqFDJqZHeJ+MIV+vdZ2I8RkIZtRq6bAlQpKRG
rMoLiNwYh1v0BC9Ehx49biKJ0tjMwzgzxALTxMTJs7M4oVkNPLRmE/YX+kVlhXO66hFivex76mDq
8wmSO+FOhV96AxzuhBGae3pruxwYWhoXMItXyWctxD4oD1WshJsOWEOaEqaHu7nxCyMa5aAiVWXQ
gstcqhTNDEJVWN/hLlUUrR2XGET2dFt+XKI2IpgIzEjEbPx+paD6N7TitCmwC69iNBosI/TfkeCz
ggf7bSImHUaeS1LFkkZiS5jmhuvQXg47zI3pCDVcoFuegmVSmv81CeZXJrlnduxbF0Xxh4fqk6aD
268gUl/vdm/4TDP3K61xim5bG0w+Ut6M+4NxrU99gyefnbDhad/Tmdtm/6sz6dZcQ29yJxRDuMKE
mBQgk8u7aAfOjXslrCKowBKJbZw2rkzI3uQP5KrAfl71c2e5CMkqIPnBX47d2KqKVntpWznacz9G
wslTxk1Fc6Asg2LnjMOLAOIFCwXVAAyYJROG3uNWHtU6rPevRs3zrs1ioUudPBgRdWxxKlqMtckx
lTdMBPgk5qJqnYer1JQ+l0Jqd3jv8ysG8jHXEzfm9y/bax34wzHrLGZunOrec1p9OLmjwhpctyvX
JKhJgtWpbpNSUFXVoL+DcH5TN2zXRPoRieWkV4idftrXE0w0wM1AjYoU3w7DsxykVsPgUidnIfY9
I4FDdmNehfSf5yG+afrzLfDRwAMASgvJdvA87hso47xns+pH/zqIdCMZ7WvGwVWpWtupYsSR/rKR
V4NMjfM2wC0kpQQUips83AvoNRaDNigZZSXRM4t19W65bvRN6RhLBECa1A6cEhfyAxfieGuK7huv
2fODPUEe5/Au/Gzo8HEZTflR6IVqOpeBFsehxKjHpDmdU0UOUsDZeQK+Z2j/IfEe0FRTYLXnMuyH
Kv+8RMwprw/I0XIkIXo8h9CJvGq33kMDAMpX3n9Vjx41qtEoY0/Gcta7g9Z8zDnnDeZwI4MRcKWG
c8TnEVn79VWQxlZpa2cU3luuzO9ZW35GWgvwyv4STlvkqFMxJ6DwNx9heSGOVlaUlx5levs5UksW
i21oqxWSFk3I/kmiKGqmAYFRPQt2YopAGsreboiLTUQX2Y9tt0Sa6/YaLqB159S25HHStCd2V+Nl
14L9PR1BHGQpvJ6wbi7lI8JMOifUSIcWoGxT9DZGNTBN07fl6Gg1FruJHZjvkZPkq3Nqh3XCxUfs
TbnN6zaMyFitHFS1EuY4Xc2B0RXN8JoqXJ3UQ6uzbDSoSL4Jeh1KQCAgpzlEt4a6zmryp2iM/+Bq
VcxLJw9p4P7T4NbwbO4JCdJjzfUL7kassWa7ce1Hs1HEL6nF6MbExph6Ic2natDqzUeTU5+e/UvZ
zCuCszp5bMYLop+6B3dFY4tSGCFfaGg0x5edCY2t/ZUKMZ2L9Frmwwgb7VvofZyzgcW76f4KCRdr
eAb3Cagw4mt4VWS6VWGgB5TwqNkiwccjLYaV9aJ2mNCcGuvaabXbwxOvz4YygzPAHF1KyLFU8Yba
1dSNl7g6Nb8EkDjQjPf710Sbsxrs7sVQMtRC1coOH/HeWh3Yg+c7oEAdd3G4ux390UFXLtJJnV1+
7WkOZ8mUZg966B3U+pvTC6Fs/wXFXmqumY7o+WFvdTKBV9ZaXGNPZHTJHsCYQ9kJaZwTF0IlZoqY
JjpONTdGmdEkebg/fhR1fm/F7+pRn/B2xdy2EXzV0lk0Gx+yaiYsMp5C+iH4pcTkxrUjPuxrh1X7
jIGRnAb1l+0abe83m/fd0HjYZrpa4+uX6UsHQsDevlTiKTcZQQXBUz+yAjuUiWTeCqs+TejI0Wdy
CcH2OOf/EQUJfE3ov5+W8d7qwEpJYNZQ3NbkY5OYAk3B92mSvrJMr0pFuKyjUWj/y9a6iB+Ct1Ba
gnj7SEi7KeTgAVlzHYQA43CT5LmW9xf0IbkXO4EZDrLITjLE3qscPNVXRr8vK9zGc/w62ZnQ2e7Z
gFYEdcbTpCIhg0TQT3ha8Vf4hOijqFvUkV4fbGGomaJEoks2pdgNhYPGjuGaiZmeuWZAt4X/XGiA
SDDP8moZpU7P2SJuKKkZWtLZ4V6EdS0aEuSaiqrJrLGNhubWA2jHg+0CFyn6WnkK3qgzon7bhp/N
zEkIIjDu9f/YJ1I/TDBNeXqhy85EzsQAc2HHy3t2JZDsQSXtQ4DQXXL2XktJLW0hjkINerWFY6wc
YEmDhKX5Q5ReR5u4QTn5wqiIaMBd5mWZOgNWqB4Eu/pvf7gnHBGFn7+wBnj9/kbCwdmtRH2SFxaH
s+1G+/kJIHYkqIelAkwCBfr9hf+Zj905vjcT4CC9euAxeOv0QIT22Bb/4Qrbh/lmZvBgvW4fZt4b
c8JESEn7kyxlYOmQjkHPdwMc8OZBtkcVQBV9VGZaOEYNiVAfAQ5HxeeADgXf4KlY0atNMTGDYL8E
vABNr7p65Hi0LF99VvlJEPTVUQbim0XKJLSiG67kglHRZpCh+FeJb431CkkZriD5G2k2tUMYfgL9
XJlP6ZYE/iRnT7O48adTruaCk99H2N6AnZbfxyq6cv65cTcC6TjzMbwCPtRLr/RETMAcgJfoYZOE
qoTU26FjboE36cmk06H9B4dOI4ZB1BUunePzA2v/iXiH5jX1XGFSYrwUrllim6fZRPdBi8H802hE
CDlXI8k4bSgPqQNZ4vSE7wnF2HZkA2AvNYz0S9sQrn+/3g/nZ2QffOqDtuBYxY8yo1E3h9njaCxd
IPZcze8lwQdGAeMYY9PFuSklpeHuNjSaikInyN+sD1YLJrbWXbMB3Zw3w6CrL3tI++MS0VSnlx9N
Im/nKlKLEfYs0wQFejBu9u+WyGcnpyBk8S9EGojzxlyAuBJRklfTGuQgDIZb5au9MriOYMjgw5dN
tQXYfs0IbteBt9GdFLw47bK+O3phIUg11kWrH0vroNjhQhyOiIW1fVSli6NH5Du9cW76r0roMyuo
qOsq6lzPZOL6eF9Ew3oDSVbwQP7esoDytZCQK9NK1hazYH75pT584dQk9m3jE4Yz4xi5Mc2s1egk
sfKHU4wXDpRKg7NtZIdgWm6jXs6rWT4MJO+A//xGDTpQdH9sjGpA2cNALwSHnI9gzF/UF5/h8WPL
LzLwn2MZww+354Rbd0SGDCPFimg3VfSlizYq5SyCbIsiq2LZ371+/ivZfAwTEfLnhi1hl9fXpxom
umPHzyf3qqpYcB0pqG5w+w41TZasAM74NIZdZyQ5p4JFKG0zuX0Z3BrCmAepCJFeAmsq9wI6DBtc
iaNviZRK2mK1IN+G2iN/wI6Et5P6kO/UYEA5mQDnLQS3n4vUGOV5SqedlYiY0Cqk+ciOltoES/0F
d4etGsMdwv3+Rpv6iNV49tTc1nxJVPebjFwIaUTcDDQJejVaXHg+GFznbuDeBUlj3mcoaiih9BDu
J6KRT+xh3zwAVsGDJiO7MOkF+3GLjL3NMr1Mt3NUvB+gZ06hh8KS2BuBRTzqMQaNGDzRJCsiY4Mz
zSus6NlPNFuhcs+Ee+Ty8jmUGEciuz6UZw5JGVov3FKyQHD8y9R15NtfW87Nfq6VDyqFAW6YI/JT
e0vb0/xHt+gcwS/Y0FSZDAvde0Xag3Q/f9UctIn2VRapVy0+y2kdr2bReXOWAv+hIisgmlb7EoYO
BHm5JqZKgQg/kPmwqjCAbbe27TGLitUwVfkHrNmohLCPfqQZLzSn9L2kW4yAmsCULGSdBP7MKHOv
/5fbNQ4W7QBraxaAmRFcaFTbUQH0v3nL3Ldpa+56kJV+x+O7GRuWOhKHi1Rqy+IgLDckPf37v1QT
1uNE8d0GgVxH+GpfsZTCNrMC/bIYDHHln1lT71cuta8Nbt/jNJR5abCvLOnpR58DdbcRdu5AS9t9
vsUreKgJ+i50YwRX5XsGomgJTMcPT1qDmU4Q8UCVFvpNpbO/jjq16WiFad934++vmY1BY7/RDkSv
YvaPI50L2gLrXgZu442RERwAghxUBJDjMIjD1z0i+Kyp50CgQGMyjQUG6hRSS9CqFMqcrWGmQQOE
1b9ik+FToBXXIVrRhODKtKPblZm/683635mAhs/ONfF/1jFP7XSKhtQ4iX26Jf52PGsV+NNq7Mtk
lf8A3dJhcsy7s3k+4i0k4CUC+PInoPoHnrMaJvWhoD6a7cnrL2C6fFqn9Y19OWiLLYp38iU5+czU
/pOFgYrgf9+xtYQ5Zztt/6MQHILvBwt1nMGGroT3JTFzZfrnrjA20Z4CjVNh4jnRJpZhgJOMDTt0
BJ82z79CIFVlOiyO3AZdUQ9c6HmX9nmhVeYsLkwOGuNizJ3aaD9gG6BdLXQZuE1fGpXJ+PXdgLrX
nSFKBad324LCdi7RhbtM9+Y5qRnsPfY4HANttUth3kbkkTJMYAy9T0FaEimltr3wqU4snS9h5JKH
rVMgWpj0rJMveIzKA0AhWfW4tRjjbXzjtINBxbjyWy8C9IwlXAW1zSgFv5vqGzsp6+5rsMUiBgwr
fnQOZaSVAmIaqShiIgIwJ19B0fDc1lXEK8e4wmJaWtb/wmG223DHGmPy+DZSnev5ovsxaOQpwawx
MOk62Gsi3JbqmOSvr0pM+cg+6VRo95zzu4Mxcmnyre0BGQ5bWMgxcLNQw8UUzshjUV+YiH6lmM5i
x4sDIUuA0MU/kHdVX1pfAjUSFV3E1Yo3u/Fw+F3PfcDNb2vCJgsZPyv/q653pV34E8lBfa++oBt+
Et/YiOU+eHHTE/NqzXGS3OKtErwMBQ/Pz4l2iw/Nv/ipFoJyA3+3RgWBYp1jBexOJU5rwjO9RlN3
ufT+P7xTqDi/16WVsBbYqgA+EFgzwiyIodCh80F0PvQgjgkHH81MnxPR0PzGHBdDXWj7C3W+U25e
IMSbZzOsvA/oejaNLtvlveSWPXVNgIFEnWXpKhRJa8sMM+Qgo+QkZxh6+N7oxlz7w/lo869SbZRO
AMNnfMOywY/iT/FKdkJmmPtJLx9DVaz0RsQGjdiFJ2RVFgpXNnUyIkZZ3Hy2reSJ5ozqUPD4rTy3
nEmb6F/MkkfCEilYIlaOF/kaulvCKEsq3owdei1pQh8BZ6s2oCpPTZGTvz/R+noinE3Qw7g1wMUi
tCXUWZwtEhQAvJk1X34k9LXSGIoRbufaZB9oKZPdyt5D9RFfJeNjjM9G9NiK7+j4kUgPvCkZ90Li
mVCPKkpyRfXRDCo8EvWIzAHkAowIzu6l0P4hv5QZ7QjrXIIa4JtQUx22+YvzVAEN07PjjMuu5S2e
plDuIvruxNbawdpl6MkzQsTtwiUM4i6t6H+XDuOs1VAsMDpIcFk0SvtnDRK6te4zeMjLXCM88rXl
JmqBKLI0h60VZ+sJMtllDbVGNyP5k3HZYjpXQb+VgVhPKzx0bPA8DF/Hbf4hV8Q8jXipp50RvEHj
u4a6WVpT7MlWVTpdS1mR1FDwlhUfoqIA+pADboU1G+wQZ2JXCXu8kOrJ9KRx47A6/IC4emxjfS8O
/hhrNKCp2zmu1IGV5YAdEPdnP4cECGPCjdPlhwhDbhkHrj2VPtNEdzGIkv8lv/OKeTobJdZU+8el
y4zrXn81fEKjExelwpSz/31h2JUdWBp1Dec9QFPZZI4wPpRLGYkUQPq3GyI+3ggBYlHDEtSdVD/U
f7bwsymL1rh7GgmNPDsIFfFWZrh1U+9e6qJFr97q4Xb+fi6EM6SAtIDSNDchOihbiIp6U80zqxWs
BHbfsZHzoFHYMuomYUwVwg17rcOaHykkwj0mP/vJwHsZW/vWg5bj+vdRNJj2DF/ft137SPplhfuH
ex/WCHQwdV1FqSvh7Q4PjJ1ebCK1aON5AEfoyrSP0qjwXWH61hPRaa5LBMFBPm1t4w3OXOK21QUV
06HxofuBsaKmpW5AEIFUVbNC59SW2AV4e4AC8jzvWP/oYSfg1vMAFQxAL+wdU7ExmEI1p4ftMceB
HopVVvhaIQb7FXrD3c9dEbS60Nfot1rpqAgp2e6IwVr6LcIhQGuVN4Crd1Vi1t0Syxkup3q7iRuM
8gWIolXWs8ej14kIfXMkgSrY98pOV7QOYUXt5sjr1GWDtEMpHAZBVt6lteSCPtgLzJlEGsBZW0O6
x5hdYtyxuoKu15Iv+IlqjQIuM0USYPRiE1Timuk20EQ6u00pS+oyydNGUonAxUjg5epFBolfRAMH
KlBYb4liOffFD5AdTQyoNuh85aLUrG2uCPle6613rprA7QzMmFJVbud/hKUriXk2+BIVea587O+k
9a4VJG0wAz42Blvk0bB7T/xgQltfqYE8NthOlxhuiVGjuPMSx4kL+i7Nx6nr2gQID5HQ0A5RcxUA
8x5lURAJ1+iLyn220iaF6MbrjMqI2E5VQg40UJ0oDLGza0wgQGshFcRAdiCyY02NdcYo1gRmxk32
1UCuF20BZdYHYvRfnZ0L1Ek4e2d0RQIIJfMSpGt+A4Msz/5z6Dg2FXiPiR5SWtzn4WPWed0A0oCD
kdt//CCXItxeXnMxjzopmM/L9C5R/RkhE7PlPSD58yvyBab0ijh1AHnGz2LJqYiFZwpw1L5c8Tfg
+iIsYF1K8etVT4+Q6h3J5o8MeNNBwgKo9qaPDarSbpJ0Q0Lk0VBRyFSm1A1Tdpl+6O/LWiadLtDs
7PQlLRpOF130HDzSLQY82PKY+mnHPIQUrIuFv3SsJ7v9O5yMP/i+yhH+tG1MwBRwER0KVPtlGSxj
vYS24PInylQ/keJcpOQkEzkRmsobJ5pAGDjXHSRciIuAQVNtNsNXni/eAdoena4dwbLBn/Dt2nzP
naFbKp7K0cW3F4Mv4SnSfOwjlMBccJ8FSDx8P18O1G0DcFiFP8hcZlTXZZXuQ/wtpHaYrOBwLzLO
9eeSEBOBT8fOhb9ZlmI65kk/pFH2fAPnnlYF+bwEzTgv29S4JbfwCnow7h2nOP15kwKXAjD1/KZR
7H0ezuupLHEy8+u8yMYVhxnrUGYfEYrEAfghgxLe9SucrYFUU22wzpEUQn+sajWTQ671kC9SB18Y
qNIDUDnkLkTAFJE1wPapHk0TJPxdgMm26y6UFpP1zamxHK9GdSy1Zl1MQjKHX49mki0EYBZtQnp0
YgNdOyNNu7l8RHrHpCRm+fo2iNIG5RQ8Kx8ih1zzUkpdSXbOZ1/XWmhcYGx5yDpLOD2k/fkkM9vF
YdV4hfV9/AX5Ciw9aDJQRqZksLHRdhOgtuEPWPAykuFcTSHI76QlR8Lqd1jXmjRBjHb/IK1tT7sJ
atfJgAuqlGYq9cOX+nX+3QAgKo65ICDCcMaw1eLrdBnbHHkMH4HW/TeG4d5fj2VOJX2YH7836qRN
RJnEmsDvlSJYbbr50RdkEzslhWS7DYi/cX9YfS1Q1dZi5A8+FsnOalK1xGHE6hKPfFYkeEdbTyZt
Kqw4dUAfwUVMQGdW5yVDVQfoJ32pAUT0Tl8ycyWL6aWex9WAvxnYvMeqmZouxbMvfFhPwHHVRBgt
yb+N5xjYkEESddoTkTQ3E9H/Vz7V+dRqWxzHtSici2u7Xwwfdn/D6ZVFZaqZMGko4ecO+cIKWiPR
oXMBEhsmkmdmrgIfIEW07oSKmKeimxZz7bgs9p/p/AsRgwKDURFg0m+woXaICAHCATdPIUDaaOUR
kscz81yzA4YsU/MFBauemQnL5PBgBS+Q1Gbv3wPmH98/yJE1QwJwct43zsYFDGfsZAWTXQjK36yi
JUKGq6BwpSXHI1j67J+weEVrOe7vbMcwnr7G444ZjT10/cQbdF5wEW8HZDCyQvKpqgQTAv013zM2
bYAJCDAZYO+2Eg29NADW0+Tgq3F878SvHwe3fnHiLW+wDedyfX/F7mOZw+KVBgtKPFJmKw5pRFpl
ZRhzQDlnRqz7e1TMz8n9mMUqqCg75+wV8HRalDAsLtmQdnODWEH4TMphEY92ksFc8v2tI8x0wDr8
Qw1dnNjjKN7JL2RmOyRbwaD3ZK3bItZ2jkLdGuBuEDzjj4sg+Tlf8UZE9ITlw12GtnuvkOeKRt0g
MWwAWuWltDeoV0zr/XD4qnEkOGxJcqGL2fazZ3rQCnli4vjDy8dFhTRba9tMxkQPJalXb7NwqWkB
lVNr886JF5nlKhGoE7QvLCPYBSZtWc09Kqvql7Y201ogDeNlqrwMFPc34hbBAlsYd6/FP9r26gxw
DEaVAsNI78nR91RW9U+GnRLIvauCvzQtj+5Z/usr4uEfOv2B0X+q+ozv942DsYg7YyJdng9ehLWW
SVm+sD/+eJsJX5IODjMa1rJblUNPQyOG2z1dWIwYMHbA9+ynnG8swU9dgMdojS2uR3HA7PVo9cdB
04P/uW3dC15y/2PVQcds+MqTGzB4ufXJyhzkL9VIDDvoHz83d8LwQwvi9ktOJOX3hcATjy4wcq6B
QHRp2s2QSJmpQ0IUya2h6ewoFRmrZe6E6H/n8v4iUSoCv6R6QNEDlTBg2e1/vdgNdTABdT8zzJJd
zw0X5hsh0K9w0RP0fkR5QgbTa2eM/qvqGoR+gcTdn4w60cap44+Z/dQNTjGLnpE18CKK2SOCtMcz
HQ1NB7DcDB1xxF8P87s4qRjy3qOO7idiH6hNDJS+A1JhcPhi33iCkKYv1QPGeFnjPR+Q3S2p5zbU
F1cbuDRlzPUQskEwVg1CVUBl264f7xPCanYtUOcQamSydXt1z77naEwed9t15Hkq4++bOQUFZuA9
MPrCyvFc4KFQ+kCAPrKYGqOzwRlTKRSP/SkcJwhwip0FyBxXz+2EX2BNLA4nqjjwWXpxanmlaaQA
u/dxAgSAgsfpPMkZwn9o+a4DMBbBUVt+ccEAFZLJNWB4R2YePvk2wFTKKON5iB5ikSwV1owAGT+b
RFjPkjhz3ybsQ2iQVrJEkvtMcMMp4gvGr07EKGqm6qhRHG/Zz/MqoTsX4FEq2eCB5b8L+/kYNZJu
zObxEKyGWN9od1umZet3ToV8+seR70hfQLkBu4biKZgKY7b7TK4LJe6x7T1q4e31OsPUopSnpfDu
ERwChwoxR37x92uh6SLLXTETrQA/KGtQCXQh7wFmmC+P36DgKKoToI9qT0Ct1TlrIexqYZ6LBi1Q
LP26D0TSFI9fOgOk7zLdC/OchHWXKfhu6pAbfiV+ODA8d3Y+tSTC0UcahnTpVS06EaUyJ15jkk2l
PdMQbtCz+T9lvB+TmTSqR2bH/iZ+L7eSxTsx00OmV99qo2OXJBkBcD5z0vO7gAWurfhGyUesGY8K
yTfy2IMObomAYuPm+0gCoyotldVfApVCtseKeSF0VnUCrIuarsg7Sg9mEOOzUykrkvPTd5RlFW0C
5PqlqulY7/2398/5ZHqcv7M0Ug5sypV9oSd+VodwvLo/OUL7LBeKqkm52/4g0pP9WP0Gl+MRzrRo
CBWfpw7lUWJ+vDwAcm02pqcuK72tdrpHj5Cq4yS9d5DzftXOMa87FNaeSuEbreI02Ps3gRtntO2U
F2X1Y70HLStSXBzfOzRRD7EMGxLfmwd1yLNnu+vaBflzjuLUKGL5hdKYwzuaHN2DSJ+5FkKDOm9I
BirGwzNeyptLTVAgUo8ADWvd10it2xOvA1+F5Qrl+awwi1v6Zc3ZruUP34SVohBWZfmKt1p1INqj
njdu53jWjEN9SZaHTmEAcPIb4Gi2tWdr1ogKaSENvyONjwBcfK7a9jgJbyb034XMnDAzHcw6G0LI
lXV6tg6XQEmB/5L0u0JcqL3lupM9Hy2G3daxqbZC0R0koigQQVkOIfP2+5u2n/j9btTXsgV59+ET
5H7IhcregJN5/gQ7u/1xwhDISRkuvE9Ka5EqpZgmcchmjp5tQ2aiVw9HK8bHrFl/VWuMbpK7+ZcX
Td8NIqla5XW+tsrcPyj2drL74Ameaysx1GkKq9IW3xomfG1wN+zsSpRmRerH+JYLOAzthkoOwteL
LB0u/M7+OZvzL0xSk4RI4CgbXQXHC6UTzttzGWGC/MqW4aZ03t5Ml+JdAHM+ly8tXYPQP+QrWyx6
+kE1sYvV5GcT8uHzJI2q7c7lAjiEVUd+eKrt4hnVaUq8IBNHaZ+59YKE4ndu8aPDD307gzcrbjeQ
86QLPAobgWA1hniM3w+hmfkusJYtfY/f+jVi6dXVLxe+iIU+8xAo6RmHXbSKpf7I9+b+mm0HAf0m
hVPdef8Zw65LiMxr3N+Y9j3ztWRCYkqpga0W8k3jtNa5Rm//glFonxB3++PSLyn3tcYeHbybZlnf
wmJEFNEF0GKrIWAvE2Sc/dFpEuJzbsIs/+5LY5c1KxDGwPssclyBmW/rztdgZI6UhZr6G/58qm5i
zjAvgwVEPohj/b6aLaUm0jeYR5klTq1vU7aw0ESOJwI/ZMQfR/hcY3RTsrGNeofuHG5qRZb55TR+
mA9Mc4PDEq0vMrozoaDOP6U4Ap3K0xO4KHJYxRvSjVoRovMF34/kZleSdei8zPHdtFe8cNkgQNnJ
ahGQ9e0QqZBCkECCJx6CDRQAujWGm6vC6l4l82i4pDdBQG1En273mmm/x3KJjjhMSEYs5j9Lqwzt
3pmiyY72xj1fdtDf81i5fqQed0e/3segnUuft09uK3NB/akOrERJBKD4RZDYd3dFnTQA9VWdxR4v
HmtcMdN6e5qsZaBirirUorDhWHzYzvSMOfNZ8mssVL+2LrEWZnkdMyDj9XuzwEQ5vRs0vgFaIpfW
WenYVUq1hRnwaVsGbLW5/70RkN8hznYKbGDsjkg8sNgG6UguQFHfbKicTNGuK5lhwuorRoDlrnad
GqGcJ4Nen+U2TnFf3Oj8Wg37aumxILxzW/u/t3fT8rxbYeBhzkT8d0Q/2r3Pi2t1GwJ45z9KNPjl
wdQMhp0Fm1hXLiM2LBy2IC83YBzhvENulOdFmi6lvSbl9UsIk1FoCJn9XBm7wyYeXy5CJ3oR0WVx
aVA6ifkEAIBK8/+PGdbZKAvoYLLT+hYRfd7bzN6h44BIPusJJOeapZgC+PG3ScGsnArJ7fZcsc3m
3n3zUeBFYBbVo/sQsG6Xhh+7E/dJhZ8yGBEzFCq+n+mzdFXloB810pOIMp8WjAWegRQMQzdWMlYU
nyx3P2q+HehYPxMmDuCHJxhSmycleGLEFMQe7ybbfW3rGZ8tlDBFPzmc0PQg0cq5a/TOt1xA3eBH
4s18BezlX+KxvJteu33EDH9mrGWl+m5GfPnETTNUNj677atMTmwmbCcCKuNJdvs3Xr2kkpslqW/w
m5nAcKHQCS89107p3RxbHlWGab4ag19Iuu41SU9SofJzCnFbkzd7MxvkEsdjkRzesYPtAYr1cKUS
WEY9uujmZ0xHxn52caQ2u8jmc7UEexkiTNY4/Di8JsbmO8MutJpEzgt6hjq3Rx/dr7McxvR8fy9C
1Xghpll6EWxD+qGYlRzs/v6dzQV2d3DkeU/VVFkEen7XcjiopoL+T/nbG7EvZN6b+f445fkIhjQE
za9kgS9WUdwwc83taz3s25+cGpq6V3lTHuNhfLGRpqJSeApiFqeb9iHD2FTp2l79DbZishtolCuE
KLhwgSpUBE9DimCc1JaR0scaG+iWNJ700/63qZPr3vUO/F9OBzGi/qLEMY8PQ/QW2ELrmnZDKosF
O8J3/TQ/7FlFDJ0IK/uqP1Z8RNPnx+Yn9i9Q59MPuyilZLKHo4QIvdpWidEyXZ/RT1T7tlLKIngz
z756hMYmmBLxjKT//Z6FLCQyh8B8cSSETeiqMp1q/OupUTRANiuizula5sJTYTED+v7sgxLtInHt
vtrh4mglfWffs8ZbFB3OQX0zBFyz3+R8MmSXeAoxvnVVde5U0KHLG2fKbUHR7Unsjiu08jSow04T
m4CnhECJ1UrEp0VOx9AAmCu1cuNWGnhP2KCYmDIQ3heFtaIi0ahzMpjm9L5jDMB7Djh1LI3t27dd
TQx6EZ2mpUAu4dUmsgW5NyEP4sijecOn2sxKtbzSxqU+BOjCUhYQY2b7HKccYp1FdRO6InT+JaK8
08P0GijkBMbsjKfO8R3L0h+TtnjJG3132fNghetTt9iiwcgTQrLDHgBgJzkIEX+4ojhq5PIm72v6
5hlidK3JgsZ8f9jwmlF5a0Pyqj5T67CuICRrPw95DgWWoxx8XtzzSpAYq4O2KoiAXdtD8sjqxMAC
QrlK9Ecl3jsEtopXpOprsIib4zmMivV20FV6AyrvPUzhscmJcWaSI0uG+JQchUHloIhvVUVd5HN/
HLApTAEbaCvn7W0rme7OnlPA2EeQb6JAvGcKBLv8eFX3VPG/9NU21A27QCC8kbluk3/Br9sc6RRt
XKNilVdWTRk2NwpKbCMBhXqGD175I/Sic8j9God1TqaEGQLmnZjFzJY9ef1i5izKSzCGRMXjtz+x
bfNgcK8vP817rVwvo6Q4AmFbjTezWjsV88J+C12CL39aasSfYhmTi2NHK87wQ2Xiat3zyIt3POOT
7phEZV4FpsozzFN9I0TsRs6lnqBCa7Y8+SJrqMW0qC2kQShuku/Vf0jOIOhy2JYrqllUsIa/v2cH
EwxltxhtdNJDfxXUiPs3BYQ/6pmu5wV5tpRWSyGaoRVKtESm3jSF9wfDkszdzhtanXtz+41RjB63
5pUMjxYrpOxtgJU6u0LKLYd/7KN/9LKO/ji+tHzw9+RzOSvTMY7+lBZsh8ISTqr9SZ6BjD7YEUyW
J7SMi94B9TfYRpiIFoQsxpbGbD7CqMwP0y+XYjmGccWMmcy+IFV49praSpBBAtAFFgl3GrX3Dysz
zR+GQMUkCOtRdV0+Q49g+ZlnRCUOYM2E0+7lL+aBKKvn5QLFOcmrs4s4E6YeWI8eapL3RzoHojSA
tJU+6nFdHg6IVdWsMsTdpE0dfkFd6FWCdN+3I5KFlHxr4BKdJN27qc0ewrrUH+Vg8dgVrklbioMU
L++m0VR0zrIp4cddmMS7jqY2M3vkQWwbJ2tbqPUMR51aQHPfVPxS/eNByT62Fon13i5uaMzXEQTu
3Kk8tX67Ygi5VO3Q55+9Mfs2N3Esg4UaDN9GrEYUZhNIlGjJIq5ZOVVn2Uc2LJmN771GTmTGBzaB
1zELP4P8p6AOq6LSjZuUBWARMC1SC7KFXolLw09HbksxtoatoYzoim3T5tP1RCdPb5o5scWRzqBy
kvsMDpnHCIiKYNqjuCSI04KaAqaFfW48mqbOwuquPebs4sr8QId+CNcW9AgQzCE0FD8zso44aH/p
Mi3d6S8A4xST1/YVgCDGMJnP5MWJbYZISijhDdxBgPr3Mqd1gCk36JlkfWdWUEwcPtbAJw48unoy
uXvPdeQzX5LRv38/gPVXxpVpb7BgFqjCak37Qc0NSKL0jw/YePZrtmfNBU2Nt4UBLGPUzvFCv7rB
6gzfjLa6LDUUYtQkvzbBZYtvimYjAVmUCD6rsG5W/zns9ZX7Dy/ZNFkl9ODqDwidmfUJ7cCupe99
WwGDBAJDBA8nlOKH3cIhKK8h4A0Rmm7SBuFKh7/aPK62lhGfZCsrKzv/ei27ppgZu+ocqk2/8txf
PN0+H/xoVsvmju5X9B46x37bIPS8wNTvGuPe8KYRLkKaivLLdpybPifcT9i5fzA6x2IROL6t6muk
VikVnTlr7ft93DLX6XkcMd8G1oI/q5IaaqlKwJl0++XG2lnDUbyT4Gy1ae/pjG7NCta6j58IXvnh
NyZj7OJxC23yT6CmCR8cqCX3mnp8pZKwk55wSIr+KVMtPH3z5Z1Wk0XNLu5qWflWO7Uu5grB6L+B
obSn5zfqj01VFWtYDNK0vFbHehniTfjf0ONXIrqJ/vL0f89X5+AkDhetfcGtrtOfpOMxW78qW3wP
XkAiAFmhGl1KvRpgjGtJ0NIfiCrT6CdjrCm5ZmhfNvx46oMHHzkgcmdQ3C0umaeUtg5j9G6L4RwM
so9LtHRe0uspr12jcE3WZL1/BxC2r2qazAA0ZwfCWQiOPb1NzGMH/krNIwm+YznHoCwvQ6D/JvgF
TsGTnbeuLmevloUgYiD0nXRf3TBTwEesdJEW+KGcACLDOIOa1VqGv4UnSMdhqxlviPpGfpy1PKGx
MuAD/4yn5EMelkihH9MNpNFCcuiuu5bu9o+BxQC4nJb9lsKy1n07xs9GzMQLqogdGNMhCU1YV+iL
8xKK1tJ7Ih8gy64nnw2wW5/kZUFf2tlDfDoBgGZkU+Gou8Ajw3woJ9lEYq3IdOIhgkTreyGLCWe0
P/PBrKFAtnvN+sQ1UdOlfOg7Lg6Mxe3c7ICQqmPYQOIMImc2uQoD2WzqiiF0wdn34Y0sgDQJrTnm
SU0FHREB6f643YMuSshMSzZZOuYOYF1nq/yoSMEy0X9HXsGcBp6OWRmd9EaUeUNyynniI+STzNsu
4nouoTF29UpN9U8Hv/2/Va8KQ+I665oyXvn2+8kNHIPMSDYFdG8Lvv5Dkiun+waF2F58Gz4FYbjr
Sy43ziWrysmGRyd4aWquPj19TTPPT0aNqNwOP8Hu5irY+GLO8ClQkv8oWUSi5dn77nNz9FSZfSpT
K3Q66gcV13Mmk4UKo1L1fmlcB85+chEsP5n8ArJszFNz3O1/pBoYSbiF5IWcH4LC/7K/ygHeasrF
/PWtUZA5uFHK4aMyOcsk+Wkve+Mvc1siuwV3lM94gI2qodjxscoo1rfDwLI6N6/lcj2ybjvZqzRf
iXOoym+1jCByUS1A938pjAhKxwSs1mBs+K25RMuujZPyo+LbpBwV0um17QvgweNHJ+h2jZztIAeY
VLwX3Zwz8empN3r2hu7JSx0boXXL5ayBBl7GFqf4OquWc3JCs5TlCgkjVQkdHDqrt79Z2hCfG5KA
tObAlhVTm23LNjcgOUQUZwcJTTI5V/FqkD3sXx8qSzLynwnzBTZIC7yMYg+yvVwarWi7PGC31zpw
n3gn2mv2JLct1QslCAyf4mjm6KPBMNOZYhW9shTUNm9QcllHTSwbu5JjtmJfOOmsEM2o/KW4xvzC
QJCgQaJkkoNOCbQ2iCK3ZIxUgZ8m54KJ76YT1L2iPZ94rfUKaS93307RxlO2IP1Gmk6KNxH2zLzw
fJVmESevbcd5VuTh2A901pwDG+eQjm7LeYQbHLTV8O4Wzile3YcfEjfQSwmnZmFi+8hHFpnfGJpu
sg9qqKnPK4JfLjrEb0aqJB3gy7EoVgtHL0BO9Mi/A0YdUPAePa0pgku46I9yG07pMTVBXOgxR+bw
Y7lkiItV0c7mKh2HkIqfs4kpW+/BYP7Ky/EiwwC1gZ7pUHB1n2rVPHeMO096vTCXvro4w4ohZv6O
Naa8qjxCB6ec/kT8MI1zNikpv5EA7z7/Ve1joxaorfMfDEFc9tK8DWBpEeNETYh5UQfWG6dqM99y
97IAmhS51Olh3h2fLvnKLVB/YMpQLWit0Mn70m8ZHU7m+YJPFjbeIjluiJq5aVjcivq4hXYARQgv
LyT3jbBSeFnMnyMnvQAiawIt6P5BSMH/x9VG5VCU+sZTmuUR0g8yO0e2ZfJ9ekh1yNhynQWY7O4Y
oB6P0X4cQPujDDUysWHm+SRaB8w+JTvOvcfdcqikj8is31RWCNe/Kj/qvHCzZ/S1z+kebabEWGnm
MFvvQIPnm/zE6++T+jiKpfNAPFErKh2j5XEzBcgXPdzzsPdvQLRZII0h6Yamoj+ukgnyE17LtDn0
repHHH6dIZBhhjvqA2t9kCVETFf9TSM7HHsOurtbu+W+3egFl/rHssmV3fb4UYNyePVPAeA2oUQO
2xX7vh0B2YlUl3R7VU+0qQ61utU+ibNSS2m/sKSs5EjAydXR8qbMLFAw1/kjKm8kge2elOM+Y/av
igO2HYX7A7OuVdjwfJCeuF8ZoWcJX7QHkjahUCUfKlAevR9pvMTRMIwI+0hp0CTAbHiFnvpF8ZEt
wDVk7/j9ILTv65kJLaO4yvKx4ykZdE5sPxMLaY+by14vvLDUuHFS1+lJ7tCX5RXy/+UxF28jrVHl
7fzqwHyyeuOGUoD9AGZdCY9aCRBvVkGUwSrTZUQNaDqWChygEBWwIflM7pi5UeQngPgsx+gFkfZ3
nP36MRNymxbW7jZYx1C9QkOxYP4Q752zmLGKys4+zNEWhD/JY3KvbxiA9Zx6ldtF0fimQ1X+HJB6
WyJHWHwuKsNMVoZSgjfKcqug50HvNhhw3zju+89ujKUiaEc7Sol2Lm0HoBvbB9NJ2d4OS2T1Nu4H
63wvEKsY5b1HHRoHbNUr8oFjFdLphksTnl+KDsXL3NiGNRPdx+lkB5WA+DKvpKFMzCE7ku32ODgI
nJKDQp5ELgTIIv3YBqWZyxiVk0HUJnZhCNZVujpSGKNUTOOQh5Fr0zjJvYAVmmzHVm6okhPEwquc
GLn6LeaUQinyXx2EBbh/P/Qf7sxwKHzcKNgxOtXR2Kcpgt9CEoXJRXSYjAq2K/CSO0wD+zG4k3U0
zOlsdBkzRNQJNzK1qZeLXxYWBki7A7uceFMWUQZX26ak8Ed8x10l/tAHa5oekDXxeVVptBzju2l6
tR56DOvDZ26RDsvvdpNawjbNYQbiqk87bsocKcH3pr5kzIwM/Tvh0E9N+7VThHWm5d87gfgfUaYw
KFmQ4uzm47SNz/7Fp7AAdPTyTL3MMNOAYNNbmN6SArWR2EuIqWk/Lf1ZPSFHR+SsjISfW4d7o/UF
NPPQ7TvpC8spwNJHzoq+bwa7Qwr1sQ0Ly007pTBdFvy8Js9K5LUPTBE3pCn5wVhBXlycjL/zUnGB
ArFumGKciXw7gt/v5e7y1w5ilCnCIU2+ui//KqmCJQztOvPnjZFWWySzk9dfHKgRugZb8r5qbeFf
xR303tQM8JuiFDyiG+ylAJvApjAraKRrlDRanaDdet83fNDwWxSU4yZK/dTNxgoZyb6f4/dTvmU+
n8H5IrzBoHOg+A0YUkvc8ne7sqLS8JgXl2moByloIkiv3WCQIwrNkh4X8wMOrLD9TIPo1tVx+O4E
3BJDua2AyYpWp0G+7NTMOoSBPARibv/1Mxlmo8iIyYRbUY693N7JZjlEOPczAbPoUFYEEl9ZrPn1
c/RDmHGGFtkQPnqPotKqcN3WuZRGdabWP4PQR2x8lutzs+yTf0UlU36Msoahr+4WsGagY8CUpsrO
YwsZTKPg06Z7hJTCM+75biAFPWiWfGxAc7ltR7ptW4iVHV/YzxlwnHMjbNXL2uugY81nOVktC9CO
OPWhLUECIg26ifMUIQkcED+S9mbPgYi9qR0jK3pvo+67NgkRD762/Mi7bSx9xmGRAxmvMfjfEzpz
Uuc2H/hS6UYt5JZYxRNa7rv5t96hxC+NfjgYSdrwd2j+mFVDQmn1MHNgGF9AVTTSs/RgiRCqPc4X
Tk9B2PZKwhGYmlGhGHhpgCJkEtK+7uuWvmaEtMADlfEHgZhaH00CT9w8TOpg8wddTPcw+IYqZykK
/6Bkn19YSi9hbhq7IMbl3ngOR66lUxmsi8rq6z+tbD9Uop2RbCVg+qn5jISqyiE/lyb6GN7aUp8Z
uOqOfgZQx5sOzzAq34k0h2YTY0kmsNdN1RBWM32PUhEj+cPJ8rZanVtl8zqQhCaYhJrHMD6wzzOy
dd05Je440d0ysrXlYCA3O4ciglVhfYEPo+3l48d7qtGpdTLuyhdTKPLYdW3Gsw4wIUh7A8mEsbTK
pavFYxyhGcHwzheU3tbpxxDQ18dxrnV6vFn8NMyEMgSlgVtLSUGxmsGGbY5LtyBMthECkHjvJp5T
GstnOZc1sSifpbYHVM2cjUgFV9i/uQphNgweZYwRFzCOCjQQUUakvnmCHg0oYFf0CmAWZCXCmdnT
QVeQ4+M52i5zeZ/x+FIvUukSp9FXH4gFE7PO0mg3RAwPwIaXz4WaUm5DWWIuR4HnqkndSrT/Un7R
bJArnRqtdKLW9bZ7nFewoai2xjCQTRDACUY5kPPgdONhCvcLiE2le3zV2Pg0UGcPohHuwFeHAYUR
9oeYz+FPS/NFH2ckpWZR5/a3pyupNEm0HZciWXWXg4Pcm11HFKzEaZrN0hHM+rEo7EVEJUh1WyTi
DaATL9nvvzxzGiLyJBT9SpOcNEXYsElMdchwaExGxdXfnqhNJ01+cF20+1nzCyA5nxI6EaKEMwIZ
iOky45Jp089ngr6EDQODG1XWAqKlljg4kyeVdDJVdXqiqTlp0SB+gxjBxBuTW8femJp+l/o3w0PN
ebjBXVF1ce3oZM4ii1MviP6HDbPD+PdjQ5dZBeWMa0QNsYdBdBEbdN4lQFLZRreL+qcoLqqSu8Bd
6foemzPl4IWbwQxlOUQSCFn716ZkdsgJAUjdQg6jPvowy+qjdMP62gMuRhQlGqk2Bem/eVIO/anA
OzmLx9cj1W9uzOA7KtGT4umx4K0PqdBOJmA6B9QW8x4MPrptAAKR3YaVk/zDqvqMbG3Z/3tzBSu6
6tnBWjRThaM0maYVpClvFT+M9n/1UW/ciARipBVVNiS1rQVXYWMvQ1wT9m9bpBJQ/FwEfD9G7pW8
E5CEWa3mNborKdF11IfgBaJZUrxtXaPSjK38Fb73alGVtV4F32EBAmpyXaGy+ffk4bezG0N1dBaw
5oeZSbxEoJhGbjojxeieYjUnY4ANz5dEOHLSr9EXbk4vI1UL0Ify0Sap4WHuBM0BDRhJLRXB9VIe
Z07iH+256hiaGtFy5dqLrgmWAAmwh3uDVl23XVwam/zOv1KMG4CZ14b8unxWikmaka1Vqqciz+Qe
76iuNuJYGmj0VcOu8kQgH/MZu2B2U//OJi/gEOCi5stqEOGT1Oi1FWEkzFKNSubSKIBBaOmoCX/I
+oSQvjRtA+EhJW/pDQmRzRK987YousUhBTBFKWxZgTfhxRA4mONdOwYDcPXuWDNLvyuqERZJuEI8
3sc4hfCcC5dWzFkkq6eU0c5IdibQq/vuIqgjifBrOM1ddpAV+yiYhaCve0pX0bdLJ60F94ABhfts
DcliMCxe9/wFGu7IK+8ENKGxBd1rAqzboUNlwf4UWVtohMFTdDILOk5cYhB14+jS68MN8PexfntB
GVyyQrZ9A0/4PHgElaN7b4kkzC97Igj9fgBYX88IBrQZhdPF7eRwy4l4WdXOe3j/gyrP+LbAvzh8
FLyROyrFne9pEMDNZ3HCn/VfTqqv5UaWDNW3cot5wfwjgF5qVdxZARWwRzRAg0h+HjoGQ5Ffz389
elxGmu54+HS+Pviawvp6OriMEBli5z/am+OA9BaGHnwL0Ir6+nOxyCPMn9SUyvNtj0kcIY5l8d1J
Q0WuLgE8pmbepQqQRt9pUdW0nYoaFurO7FY5GPdn2pS6LMmT4HhvAnwLpzlIBmS2rwaCgLAEXOhS
YeQyBbf3tLZ8qBG43wsKyeMIV4OAztYp5R+s0LKIkUOaA8T0vUZ7VjfIHBof+xSgBrkgnV0Vvs2+
j/layVPMm7Q4PjAMJ6jF1R1mKEFYoX+CNxlhD6FWnfPjk5zZpEtONjBnyQxLDN0voehdp20LTFg2
5C6KbvUOxPbv+/iGHkTj7frxc7GdEic7yDTVmH5k/GB4Rnm0h8M4JdsCccdSuexJIx+KoF0/oEze
P0mm4WAB+yHL/pGpRRM5M4qtJZlCfJt7NXjZCRUEoW9oou9YCX55KxI3+EjS8kBXDViNTx4F7841
BH4PVznHB6WnUcXW3ucz/2JF3Fj79jvxie0dtN9GwqfEeJVZU1iC+2ltGPvdIRVlG39BIeQZfuS0
7yu5SWqPA4vD0JK0Q6/ii/ZW5LaEtyFcaNXfXWJ2Iw9G7C3C7Z5IYVuTAZJlAuAoZPSuP7aCNVBa
CFf52EgiWZEaEG+uNxqQCkeepPQdCEwocYQ1i3CIdIdEHeCu9aIS8NryyKLhDnZ7PK8Sa5qn79MY
drW23ZcTHDXZ1MVixR3O983Kp1UZMPbpqOLO79TgrVuU2jH1+H5XXqE9CeVtL6zcCGJ5aY+HIHGJ
LYPBgzdSPi95SW0iax0wcKhcupQSXZHKKwI43YRuyUbXBKkAFbbmsJzU2OCgDL6jPSTwp2PFfCS5
ZS5xwEXDN0V36ULYoAUgFjGBZ75uStkpUyOzPOM5aSffLkGWDqbxJNDYLJt5kty3MEkWciwHs7f8
a1PkF8cm/+p6VeNRv1znNvUMfyAYV6SfsqppkETdyJFxHSV8UZrrexLbuaT4eEl+Xkjf5hkwrwf7
5zLpaMrPO67C0+8Yj2z9kKGVZ7aPMgw2woXL5AeOEFb3lkExqJNnAv4QBhaqd9vVHlSzbkaNpUNo
uZaVDe3B7DE2BsvCkJc90JDEWPjFWEmnkncvUI9wc9QaWk4KF/s/14rlUysXA3Jwhr16fztvsqjx
BUtE1Hp5CLlkSdKcA5zO5OiUx8tkl4WNHQ8LOx2qSaFfY6rI+PuFIdtHO4jQZSOJZ5kiIMlc2qtA
ju2CDgMUFEFinBeh/lkrMTY2xna6hMw1SwRlzcHCCQDEKOnHOEtEY+YIF+manCWjKEEnDVeKQPlV
hem4pl9AOSGWptLGt+fg7lezR+niy9cAwJVplyPiGnIPIRVVDVHw9LMnChDRb/bLNa0WUECOgnMg
Cwbgbf0hKqKO9/+bezuUv1FZtWnYfeJotGSmjJnHVFC58hH8S9o00igbMIuJD7qLrr/W3wmUcgrZ
NwngcATZEqfQ+/JonCAZEi7bDJBsZbe33DRBtnGjHhp1Po1lnbxjgkeAqi90k+FHwaPGNH+65hN+
HvzitMoxZOHIz1QGkR9LLaOEFCxG9pe6X9x8BtsSiYiDZpl7Zz/XNhhQSdBZ3VwUjnoUhvr2+rsj
xu1tm9U+hDLlNviXaxUo83D3+C0OdMjIjLTsMa0vRBXfH8t7GMYMGfKj3hYOpDXRF+jQcOUVBEws
HviSS9//W+lVvy2GRIfcXykDVwHF9PbGRwuFjWtnGi+06p2cx8o9u7lKqMMXh56jP2NBZviT6pWA
av/xxuDdxKoDhM1UbFZTo6Lsrqv/VaEfjpSMLmUciHCaWdn+0i9aCSrs5xzRbelRrVjLEfkB6wN9
urOLLqJPwC76g3KhKFV2XjLZDGGzoyCi8rUPfenMxkLkhWBfxdZZG2VecV/8Ii3UHNmcKJAsYgRz
5PW+VZtjF7YJm0GN5/LowVmtrwpRnI64QHi8F94NrP9buZElRWcEbbUltDZV0OYHQX/netLflxMl
SbikJSND52/93EZQNHdlK6jrSxnqRfHMFX/gCD4iZhlkc72gsPbHSVO7KAe+JlTKuav2nwFY/hNI
oyeOS58prtQ2+RqtDgdNWLllfmRDBzQj7Q2lqYTLKOEwJvvqP9HfjpmDjdhX86GqGSQEmkP2g5hT
p+fxZI6y+KkO1RbIDfvzehrvPqh3fFdcJG6e3KHUHg1bOBTjt56IbXFTBG4K0xo0NdUMbnN0EBiE
aO51bD9OquK1ejmaPaQ03uvtAmHt/RlkvWZno3DRch0Kb/2+C2dQ2t14XJNnZ8BvfK+zDizQEPMP
YU4djphnj0hm5xcY7Aqh9+qQ5er5cfnzB/TxszeGdpxxSMt6JMBsnGYjonmCc43OzBHPRnMKb7ld
S1MLceGF09lxm/M2ro+NAd3oCrKKoNH+XHEslafocLtBa2jEbKhh3kXk4durAMcjBES0QGhvuizz
V6GBgL5GPGRKSP2N5ohaedNH0BbCTXFhIJeEM2sbNR2FeHF62nExr3Qesl0S8q6WR7q1uhD6KoqA
6ddl18LHvXrcJ6lTEXQWubTUXHwH9olqB3OA3WWNmzrH3ndh7nfQlnPpD734xtPBZgFPC9DDDb19
+CjefMk3IFsCnXB8pAzclpxIwGas7sT6M4fn0gw09MPD/FsgrcXIObsz7wOG8lbNdvZfGofH8TzZ
+mg/iukhDUugFjt5NSYM1i8QOAk8hihTbDk6mGInVVTN7jkijSxIlIjDDwc0W4Fc+Vus8b0KngsP
HXiLBsysp6NvY8pb5EKng18XZDdj/QcPi4LhU4Ta7ZQfHOX5erKiFxOz2VwT9MX0XgJlde1DrwOy
GUD1wrp9a3sbuipUQQ4o6PKdvQrUkS1Yn4yAoAClQCH5RSDMRUmS8X3wF29ZAMWXNO5RI4+8ukpM
eDCjskk1AcvB4Fl/xmLgzD8dctHhIFyGe0kmGaXobaAf2K5IazCXAEpKd/ggY+oBauPRV7TaBJF7
Gxba6trO1uZlP00EDQ+cGITgHIjLINXpUi8QKz7MA7zI8sMw2xaEN3AEXXIMgyXH0DMtpn1EpRyN
ZAJQlDVjP12EzPiMd9ooSDYBaa2xWx0FsJ7WqahHoR9ASZg8SQzPZIVkwXPBtwhXqXhR8wG5cqow
P8VjTczvXSer69gVZdUTO7o4nHPHqA/ZCWqpxzVZOwCr71M+6bUEH4tmnt3ZPpPxAej8ZLBKGYrR
QR17wLx11420SMAxfiPVEGaX36CHzuFsqZjGOEOtK5tz8UaKcfgrZ+ONSaSZGIaYOTTBHdsj1Sdz
jKfg2wZXhmETvk0C5ESowPfDqoBcWT/hpVpMFMTe3+6644UVoXvgiQQxB2GSspBzHZ6DelfR+7SW
hBRAL9s6/7HjKxcGgG+WV6h3JFZdO0V92yLPxe+D/O2CECstoGHRIMwMjpRJz19x513/T+2ShVkA
jPFWofHI8ImuAIeZ/bsCHDMUH2rVpCkLIzaG+L+ToaocCdtGH00hgss82cZ2vaUICXFFIQq3chdj
pc4q8RNDjRjUH0LhMA4mYbdhx5Ad8YEKc+VzJRhdaOU7n42POhjerkcgTAT9o+XhviEoJKeJ/5Jo
JVe87+al0HVXlXip2JEUpbryAmtxtLkW9Txc0HjbBHM2zHYW5HLNztgh+PBc+rOB7cjCER9RH5VG
K5Pswo20MOexz4j3OvwBvdxJYTMa7umaF/xyZsgQf4qKcD5/En0w2X54p/CJYJ4vJl+vZbiQj3MW
HaL2apnqcvPLuE4CnmAGMyI9VnYhG3c6fKp5QmvoIhSa2NBBJjFaIpPoGwmxbl9HN0npsE5wPbk3
BKlZ/wINnN6Z1cY9dUll7ebqmHQZVgy+OwQwQIJbyWwZ1iEHTfiX8Af7rnTTj/GnX6iCDGatg29Y
Soip4wdyjjLdE6zRRWmNBFzJLtHQnOm/lV8CwY2v6/6vxF0gBr7oNFDbnSeB3ePzqOXgP5peSSKi
300VlP1lkcwbbEpWwvzoMnXowDk6Ac0ITKCsMjGJI4aw73l9H0cVELKjvPxnA4FjEjmQhvRSgEUz
dXD+kqL3sx22Ydxv+57zLMCrXhV/9jhEQq66WH9rVcFFxQSmYTQWyBeTYPVzIFRTnIfNQdMpIIvC
ruIusWzX8zgDz9RBuhacqvaayeN7pXAEqUvLMfg1KTQbF5lyIoSxeQWvB07b5Y098A3gxm88Fp1X
DqfLKD/4fAGgxWbx2YM2+iH3ULkF9UqZNHYlluazHuC8nlZz2wcJMoMBu2RLdWjT9upUHgxdItsm
NDI+gZhoKpUnmZjlM2AgrS3XSDYkeWhSzB08OKeDUhgL2ZgV1kOWM4DQNY/HxQVdjlJ2AeisdYsG
v11VgwwwPdwIxsneFdQqDsIGpiJtPjXhDEh4HeKQFmUJsqksywWij9tleM7TKe4rohvXs3+DwauS
3S4Ktn2X0pztT42DzgU/tVxWT5FEEfslBMF2yIf6qz2REpbsmLM3q1mUdAghlcjcovJvmq6w/ajB
IweP8NBTVOf2LIwmghM1z+fXIwT1HXXbO48zOIp0Lo+UWgTrO8QJTV8Xe8EsCTqlooF4C3NePI24
1dkxvTr9k+TMJ22P+9G85G294XBqpIiCREf8QkvP6aa2SkEjuez/o7GHR7vuGwGOLsP7alX6qmxK
YTmLD4OFNdc8A5dE9kdQ9HgaOuEx7y640auKPEDohFJ9Ed+Zs4/BrdEs1YzGEwftlPdRgyth1qVw
8sQUgBMMIxCaZ309uUSIBoxCjU8n3sTQersywLbywtfD7icLlVCZPBPwTvUT865o8Jvm/OQlx6LZ
qXDGiVpXXCs7M5laAelFohCTIwZTIfWkSQZWDFX8Gc3o9+qRSPWECrCc5Q5fGafm0dBaVjo/4psc
hjYej1RsN2NDUw3JawhhBbvGaWy1QQH75gI4xu5wn3XxZoHBL2X/QiecuFHp/pBjaltBL8KHUi7B
qHfv0PwBBPiZl1wolllIH4p2Ud7cFQwdIMs0vhD/DWX1gwL2jx2iBQ2iLn3l1aFmHw/fkl08OgQr
VGmHgyzbk033/ajipDdUeNmBxlFOubM3cPBInxl+z9Kr1r5RCpgtuajAS4VIuAb6NK9LeR6zOrVt
lH5KRGhqGOK216yndQOYf2mUC8hr7oGI/me2Kd7L8l4BUsDS5/eKCLm2xcv9CW0GglWwKpPbGvoD
FWxzVSvqrr0RZgscCQvMypXpthSSvjp0up1Uq2RZwgieo/ctFQ8lmPBJ1M8UuvZcG8GtpBh3J/2O
J6n7hA3xB1gm6oW5cptg/mqXAAExuCWMkXWlFeC5RRG0R07Y+GfjAi0YfGSSVmw8qd06dXNXZa5V
fixblS2rOQ5R4YXhDHwq0jDUWb0q8ZHJWGixivJ+ofkPumWHe1B7rPm9g0nEDA0/YBTCPsQmAvgX
X7KBwNqgWjoqnoAugSWbzxt9ZZi4oxxpdz+nCdryQx9bjYOETfMcaJvL5NMac1ZVutMug5pcOxxt
zaax0I+Ki/nSuiYq/of62afKzjjWNmrsaVOfvXWJfg/H8qcBcSQrd7AS8mdr5UxRR0Q3tnxR0B34
Q9bNB+3cEE+6sWhg12+fOjoP/XVa/pqssiGxBV9+4RBl24BOVMRcV3DKPCH+UuvgvsMHEjU24GVX
TK/2cuE4bRj61DX5ATxK4bzQgxxHbsTb4XKy2Z2tzjGIjgT38Z4JxzT9M1BLPvsFP9YK2JHuVL6P
Cg74jfjs8DpUZWTsezj8a1YPRSkHI+AOr8CWYtpuF/QwpXwJml7qb66rrDa/kvXrJyNqBvZ9Aea5
zth6ZhpDwYL/gJlUxAilb6h6NHxn04EdS0nT+2TQXjp6I64uE+o+I+y4y+Bor8yP0Ecp8JC1PCcx
zww7drYmAnt4N9/HxU6u8VeJrAUEO6cfWW7L+gtCLCFTKZSlmiTwLvs9YQeawoM3OfKdleqVxbBX
HkqEhDJI3fDqBLIHjGCa6D/O8FWgsywO1kVtZlRjkURr9RCSOD6fgOcn8dnZod6JGLimN8CyZnLD
ErgbxXoKmq3C0ektAh2EpuDHOTNN0gUr+IYBJJW5bOOn5jiO4bxl/l+i0WMIyIJTtZV/ws+EMUkt
qTOHsB/rtDWuU52fYR9/5fvuA+rBKftp482bZ4MnNVqG46cxnlxXk5gHO+cCPXH6VStwOGDgP8Np
gXO5JIqrXpC6xUvAc7w2qFqpUrEMff+EKzjko7fPtK4EsPrte/GrItkBa21GozcnVtP+AyEUEs03
hr5PfKwS5rCFZn+OgHsVVFTZXtA+MnWlydMGE/lnzWQaTGy1EoGQt15K+UDKr7hCrrjqsSAp5IOQ
81RGFMBLcj1aBLFfFNV2XOEGe92ZaWirRHMeIYr3aGC4nSOEWgQdYH5dYPT06H86hWM7cMiEiD5V
EZXUEyINPU0IlePnCaJHYf+7NVWx4t4WDhScqIFSe/2DdknZm1KGd7ZxPwMCl17ZAmny5JfZPBQr
hsit5iiE16CL8kYvJ0UdZfYyusx4alOWknPGcqPe000WbEfr11yTOQqdXU519gHhV+xaIC6inmVL
Wv8RbwIdp6xAtDsWlXJGAhlyMJIVIfcfUdICPvsN2pnvWlQnj67RV3V1/WJHU5e/s0d2/Gwxnl7Y
unmIH1dNwx2oSKfXEJZtHikBJ3fKYYiUTpm8EsrpKFkOQRBrrY5EFd9vieOHDcisbD8he/oJCWOi
NtPUvLY3caeyA2Ku3N5UnXcDbe0mz6mQAkogEekA3XOo0K+Sj4ZE9FkHFP+HJJX93r/hoMc8H0bf
HWMOFzktr3ZUDtc7vtnni1/k0WBhSg8zI6RHV7azhLebdOT9kyFN25D2EqJ+tgjYinVkYYzxe+Dd
OwDy1h8B369okTpysBPs7dGNmzTEbqUcTyLxqNpVeykgE4C9NyLmA9odLugR/sLbyU/LlxbuCLNL
wkI7hsbHEFPRV8nt43s4BELPlJUw53nF3tkShaW3TWDTNf0Fy5H51QMUCDEij8WYrwPGFi1GPVhA
jepjvHgKLCYaKH+igRlZTP5SGg3no1EVLxgWZtVrb1G9Pu51fMjN2/1hJX1iuvNaJgCm+H1kzJr7
ccZgPi2bxBC39/GXgaYa3RX2A7iEFd/QHwh5K4ZDjLKG7Q7oZp4OIqpwpVYT1299+xhrn9urlxqZ
btyZbImCtEusY/NXa8DG6RxAjzC7hdgMnVUyfujL6/lkS4cLjF8woJ1smQsLu6CKXfmASM9r5P+v
1MDS9zOJRt5CqDLaxYZ4wrJHlIauTwkTPOYNB5SRI0Bl/Mg1f2DL9+LrB7i8bdHqs6ar0fTB8upj
IpcDtht9dX1htGlxSq0XvhsB30XDQR0uiV9P3Ov+89fmVuIVvRhIDtQhE40JmtdKA2LW8K2fmE+i
05JmYnQTdstTFB/uaIn/4X4+FACMNS5xm/k74jSc4H/2UuFolCmQMEWGdS2yD3Mm1cUFJWb9QnCK
D1xnhgEEknV4UB1y9cuvlbO9rIkt4a6ejz5p39yNGc0sgB1ksxsm/7uRw4mFvA87EvIENWweZl8I
OBMGfA/RCzwygkET0Q+zjvZM+63L20sPpB1Ztga7t5ufSbLzyMhWYACqVK1/fEV63UNj3lONOCRv
SXtFPbCoxcyD6Mk/jltFYJegb/cNfh5oKr8K/CSwBby2MDCxbL5DWzrPIb6wbsLM03X7hzFVv8ws
1Gu13drLJXCAvrxqeHGZOquJppk5CEPvWInb3gSfSNsWYo5YgVva1Ie8C1giUaGWLXlGyyANpJS2
7iD7Z9BhiWV0DEOfQlMhQ+t/s0p7kQg2Q4wFRGcBTxHpzaTda5otUmCQWXzODH3eIUXaf7t0hoCC
9PiiLerP6WrnVEHQ6/1P8e8DVKyYqdGpTBhc25gAgYsEQbJaa7Yeu5FnMYyLvZyE1+Rl69y5skhh
xn/ezgeIBkOS4n6GzBrnmBH7f1q3aE2XePasvAKnJY2WC7hOa5n3hLtn61ThhnZCtsqwz90LnprG
jXgMCAFUP0rHUgIlFRI7T0CTVOI3lIlFgXqnQMsXb9NLvQ8tJquFs0fW81oCov5ESPAkx93KEXvl
MBuey6Jamy2U+rvd8wBq+5NB/669q4H6g1Cc1RhEDFpFLf2gBm7YkAX4qUbyfgIE84PgYsFyV/oN
1nIQAvXjY9euUypMu62s5/+EZWh1dZwrDbpwcryuV3hEVDzjgcQreEPSMZq1/u2WC7G58ygyeanw
xqyjTcYSCpNXTeR3gQixGKiAhANV51W30YnGU4olBfenso2oeBWvXCF+Ja5bL5QD/EuMtTzP0Mcx
zpSRFa3ZxtuDNDJk9Hudo3kFT/N+gxgot/erVHC5+6Uc2uqHaMDqgFILzVC775RueHyLH+LE20vB
xoF0gMO645xMdqn9O+n8UGhGUWR+S7jqPVz3PPidKEBLb2zjEWXEsnTAgulK3ybKTVrk0uc3MegD
m8lMJXxnaumAz6ayc2NWfHgjwOPypr5dLuNG8m94CAzDzTT+AGkjLUc1AGhO0k04ToUZzUxs4TX6
t+x2upuHw2f9CScVkMYAgaDjTbBzKWpuGX+EFFmu4Whx26Yrm9hZ2lylyZf7SjB5dtTETF/yrH31
oqNA6imd9gku+lCGZg/vjXeFsWlVjU51lQypOGRzcoWHYQIb30RjYTy8dsRuwTiA8Vo7Z0cUQVrB
dcEJG2aozoQvcVNz1pB0HMIVveafA4ZDmF6lCHYEzKUZ5JpWmqdcCf7J4CZM8IpBK8TvXMwNyGRv
1El6KHLLDFBQEiGfynO8B37yEyt5emsZrFP2LK7puBW6E+bo3f13ZC7W84LFNJ5PsDGHQrnFZA9a
+Y/uQh39jATvb5TgLwRrINT2dQENAbBnXAuC6yS4emO88HNbC/Dpj94j6fH9hPX7VG5Nq7jog0DD
ftI5okIfUYcHt58im1yOQKg/ZJp6ESdrtiNR4fBE+A1mbmaoAwoG6q06RvsOTENNnGknSZ1q7bdB
f7GHNwPWhQ1NGlvh0/8VbQBL/SwP8e3ITn5AWZoRu/pC9sWD+h3gcNGXKqLGQYgV3nONpLZyfTQk
vLqSdpSoNrE0NHDqiVLTccZ/gQ1qhMDoGV1eigEFyTWGrJJ/R2O1qDk5VnYpUBInQauCQuRrakFq
eG3AAcDMmV7whIOLK51ALMCdqixQf3d2pnAkLG7nnI8Efx2UlM+Dcbp8Q/9h27sbERod8P7oNdqu
TFQV5VxyN+VqBizwjddr22n8OkdxguYNZgfZtBpZX1UIR/Y+Yc0B5ByabUqyef8EVnfM6Hv7wsz5
iF91rpgkzmDePrOO+QSrdTGahPn4uk4CJXsiJADabi3FmhixoUgaaBWFmJ6qSqBqBSrXzYdQcZWt
y8TFkk70e2BTILdPSKuqPaUrJfi6Pu5QXec/aawSbdl8rPLWwwZqCEAhQSZgE80+9/u9DFkmNmGm
DK6PYAIsZHArvFLhYhI2i9Biebg2dtEnAqhMadUyyFuKquDG66iItPFukEB6AIvhxaZFaaL+Y4D7
EQTijMWaImQcJF3gmhvSuXkW3QId6B2lx3CMcUU2+kSvavz9B1q5lpyeVluLGsiu1+ZWAfy29rwb
wTkcGJPBeELCNgkfp5oYAHwi+VXq2B9BndDUpxEunsarl5Hw0tsD7e8btNawYMWwLflxS4262ZT2
mAoaQupKSQiUwmXXMfe2P39asTayldtR1I2e54L8kusqLOXIAFvcdL5X5US3Coiw+6J7EFCO804H
1t0jp6q6d5CBCn4RmrviSxV2i5ALnwKs9e7sEVgPaLcO2/J+DjAwTR5qRC+5t7nkga/BMOUZrMgt
hbPVF4fEy/kgtbTA74C6iCibewnhQ24SDKkMe4VY3weuZ2wvodmmjsCLWc5CwRo1lsvHhewDx8WO
5hoqy0hcLKCrXCjlmqcOTsxBa/ZmDeDnuOjdDzW4xKxZPahOAhWRJud5Q9cSnoq6YWlGyrVjQWg/
K1rJNcFNijPb+Xm8Ym4pLnnwTmKW0GivCjhwtcl4zj6uNOvleWmxnmrRNTszGHDQGgAXo+HBLA3C
yj65YKGyhYJLSpWTXYJhg7o/SxLm6eUjp6HifWvNV5chCMVD6kesXMJ3QCOwQu1xsllPctnFB+46
4nBT5QpSnG/9CW5NYdFksbZR43jZEVqQb9owcdAwonsBZ5ALhYzgI+IqO68DKKDqTqnKfd/U8ciQ
4O/VdMUZdmv0ECIaBI/5ab/0dq3Vh1qXPR0IDQ8sRHoeWvKQVAlNrbN6/xCxRq8chHjbxRj11lH3
o+4UBTnP2vPlohoNMaCdyfi+U1Ol1OLswwE4PNpQlOcB6b5Y9pzkzcSX22WUW5C5lfw6vOhaF6py
CRrG0Q82XbcxjzkfVyZrGeNn0Xmt7/OtRt9ooINgH+uThomeVQGzGz46s9E1Sd3KCK5tLMRzfnMU
Z2tSrwflN4IF6TJsV0Frs9iip7vYzDdLqiTEPqUxdDK8bh5SPXqEG0StrcmaySkeTkrubCsRzu1v
uzbnqSRIvZVfwyVbjo+kioIU3p1Yw/e2UnyK0Aqc/0LgRyyvgK3njiEGDcTRrrBz9xGU8BNjZ/x6
tdQrcSA2CO72GgoTCYutXnSGYpYM0YOQX2bRoLVPtN06W+qgt+DnkqzOb8x/C15PpwQnUokDVFG0
AYB9gaKklglaOLd6Mvj8EF4zBnklacO6IpXfb1qluMxGwiC9Aw293UFRAF8qoD7oPemsXD7HIZWp
qrohNX/MEhgF4dB2k+IT4sa1aie1+zABomipfcvHPZYEf8rxa+V1Um7cNTiJaS1WRKl3YRVmYSYE
a/jYzcvzJAvnF72OaUoaAEoEzM/VapCdoAGwKutJiOsnz3n1EynZ7h90YkDSSCNQ7YUinYR4o7r5
l1f/vtKdfGhGm91w91MpxMtQGqajWmuFQMddPqf4F/k76kQ2/tyLEH58GgpS+K3XoHloP/o7yi4R
Npyi5eqTBjM/4s7m+I8daG/87+n+ZwOYNwzEY5gVKCV8lre5jgDWn35w+P324yijn95X1tulBKNW
UbaCY6iPGTic42uqkj+BP38rupwUQZmCUUSdEOlF561sv6JbyhTpzjZbY6t69sZj1KwHaQ3uMUeV
r9+OxXB3Rh+D0XVL87AYxGOJzxftPaX8EjEOTQ5gGYwexQsc4YnWMLTyW0MF5uNW9WYz/jVfep0S
2FA6EEAoSPeFhSK6CN3I2xQZXAYQl4xbWXkrZCARCuxhS3mgSLaY+UYCs2hveXDySB3THc2tCkpR
18fXC8cj8X+oIQaXZa+n4xCGR66KGAauWB/Pf62cq2cnzgNL4cSKIcBIhw/+Ozppl1T/p3AitfeZ
X8NlkQmjxWmUVXNVXCPkaD05pa232loCLv5Fh4vHFzpus8G9AlOkJnS0U3wXiBZbDi/qfB0kSZAT
YhAVAum7Utk5i0RkFYwbJC8f7MP+qzBuDfe48iWl+rCHeb7fNKUjJz+jy2ArQRx9m1pquHymt0fA
TtLEpwVNb56SZafqCMeGm4eotnXLLgjhqOJj5qCyqPzjX1oEDqA62OWTQ/OShvWKs3cMPgkLWPbt
cOWyQIaHfJhi4wrSTAKW0UcBf2g1XmSO4lKCqrGlAazx/EzfmIiFU0T+HMyg2H28mZJp1bhAGin+
hjDb5z5cmLPyQCNRYmFlV+yeSzy3ZFslxF1tclkOU//rVWj5rgOQQqo63uKqb+W1mBesKXq8lr+Z
ym1GbctfZd3eaD7pI0xwKe2rMiVkQi5a7dvhvGLhUSkkEMf9Yw9e40/8WYGvSnwBT+7Wr1RTpDLI
ignG0eMfuvEh+UaWt41y1Zfa3jZ3UDF5oi+GumMY8vHMwJI3DHCHNCvs4p9vQHalW/f7PJw27iiX
2rDstD5IK7qrwQKcmiejQdAv1O1NEMGPWKW6w4rvje356BsfMQOvhQEDuuXcUaWdZbpqJQDCfyDM
7+sUaLPWTKvflGmY2EOIZKvlV7XTwF/MgXOzAuZPR6TOMzzfgLi80d4B1ns2aTe50+GdQqaZfE+i
mleqDdjQeWuDSXkti4N8D2TscB6KH0L8Z3m2pa9Q4NN9ZAzMKWFIQIc/cz2Bzc8YEfpsX2EYNc5/
JVJAbkml7beAVbwm8ZCNMGN7PJBkenEkR+webjCBM0KkYv4BDmkCsp5FPmjDrIfB/y1yRKJfQKON
WwKjdVZCXtmLi3TYwNPm6Q9XTaosqEsKyGOnKdQ2PYPhOdRcpQJdRlJfnpjVimJU9vPBfJtD51ZF
Vo/jztn9Dj8vdfLK7/dxt6kePIqxsPiOoXDyxtenHj7pnqZUoYeGTSPpSwaXo2moxqMAtm2Pgqxz
UkzSWFV23zUwAupM8wzpxTGxosf5QHe5vvwAQE3k7cD+RCt0tFClAakuyXaH/pxwB6GApcccH0CJ
GKgBHCkH67mhQUgjhCF+LNq27TRGVbQl7aJ7fIowURxC2nWH6SdF3pm6lMca4uMmrhaxfOqhPhGv
b/Fn81h1NJk9Jz4b6A6QEAubLHkN0KzHvuB/ql7kaqMh2WqXCrlr0Djr2olqvbYXsrrF4W/F24MG
rKLsSzuCVb21DCX06MyBEIxPnoZBX9WA5oZWMS8h2ONblGua8X2F+uft3tqVA83tajGo5fZ8LiPk
RCzT108QQI8YbLyMCTOEoY7yIQL0OpQrxCoRI64tUrrV46VlR90WVCVZepCe2Y7dqAJiO+ty2y/j
DBJHVnG267xvWd5bGNhK3o1gyhOCItBLOwJxrv7QPTxU9lywKQBzJzhC2NL3QukF0lC3ax1CKv/2
ANmb9Js5VEhTZA0hLkdFLM/cajBJgA29bb7Y+gD4k0iU8sGySeEIgx7Rp80tvn22Cfbmw6x0gMRh
T8fIEkc0udp5KrYWtABOyIeY6+eDGp/VY36bJotjMBI2+7hoGBzIu8paGCPcUWFGBj0Ssolv1dIZ
D7tdeOzl7FOJjv22DKAJSujI2IcN+wROicxTGz0C2L1r8DTE4Y+SWCQYAeOb3xjVLCGf+BwaQXiB
DNNi+2FcDbPBYd83rj/6pRD4/HRXLrv/7WmlvL9mzQB6S2mwIHLzrfHqjHq13MrroWXPGP6JJHDk
j+XXJHSYy2FtL+tYzmUK1Nj9+zIHWybJxsjMdJNnCXBnYqlFaM5zZUJMVv8W/JAJLZQ+nv2rVwus
q3jeNspHSeyHiqJZuMe23iymvu4uWDRwyIreeBZEQGjwD5HO+tcl8AAbnGr+ZpTGjQ5FNBdAtY5C
60pd1t39IZ0AERoRVvrLUpWFUm9ORQfjYLfL/0eXKHJNVOv8s60sfm4NBCFdIDrRpnkIyi+sFXzu
/DlaUQ+clSzbgcxWrM3vEDEIKlx96ShSsmWvyEyZiNFEDw8MiY5gWy3zdXkUyPG3I3eGIZrmFrjL
f5t0hRR8nJ6NiwSaqAbiDnMvBjPE4xn5FfcR1ysidiqDkPsJCbDs05yPl88uwu6K5SvpXTwVr/RE
+MN6fzjovSbQ6nvAaxKfWysvvU7hyCgRBJmaVn0m5A8y70apflv/2mSvnMgPhxGt+fsk4VSzYBn3
xsylyOshYQ57yxu9NsLiWAPOZwjl9GeE4AwRR8Hn3pXTO5aSwwTV6EO3e8ZZKVdooavBse0vYawK
TpPDhI/kuP2Oe2rWdHvh8XW6YiwGYOie4m52xYGAUxhwYB8Q7z0TC/Z9dw3z4RyqVBAQwfrG8ey0
+NE3Qxlu00fc0zwafLW8QNomchas9adaojgXl/ry5jbh2AkaFNgWzkC9LIen10vXRDchcvNOJyHo
pYBPUVpgLQu3uHH4q4PiTKFg3GQNXqjArDlYhiIkDXVVYL2VRAjtlX09yKcV/M4wqVNt70a96ncd
B9kqPVdVToBG5IXOg2OHe+WPxDswD2I9xcuz/HHBtMJ/n80NS4+zpwBWiaBBTY+ClQp6h1l+sIo4
h2RviE7KZI8tZjSs24oJRxf2w3Hk/GTuPKnsd6+Me1+Cmfz23IgznDGleHvONQyV8l0VhJBecPqW
fxiFMUDp4VeRAoAcIAFpphoz/40pNA40tdm+HapT6fLlXxU5Nk/eVApeTZcI8m2s7nkRl6ZwOaaf
gTyfWJmaDAgCIYZ6AdU3sZ2Z+evFyq9mjGCftjMbloxzT1gunR776dr+GHKV0p3Kege+SInpBGgB
0PL+sNp/S17r4cVypfSiC+xC4Zj+qV/tnnVbShiF4cyAhIiiBVyaMYoUuu4n3Y8DfDf1E22Xtlh0
00pUqUl/kfF7Apf3CzLgy+bJoS+0zU17w5s7sB/2n+rRHsZurm1fnrGfRalh1CaiNVCNKWbdZ5IY
RxRLZ3/FeWEm9/Egpj9LDc/HjkOX3FkDo06Bh0Tm5sxZo096/6EwNLHffQodsaNJg48Lzt42xWjB
11wxNAv9ks1aRqDtAIg9bc1sr4Zg+c052BoBzDKek/hu4DTKPDB3FpU4y5oiE29RBZ9ypOnOpG0z
+0cDxrGh2p49RBDWnDUiIQ4JmSXrMgxX/YfLJsvtwfAmjzhTwfqrqN74mBmDD/YDi8+tPBMSIsY4
eVVzzo3ECtiPgWVuohP3QMd4fBbPZJI/YnrSNuiC+k5EPmH4EtzQ416Hqd/ffedwTTvBVkday/nV
QHlnWytFBmaKV6CXvf67STs6vM9ESBvpM369mrClrUPSQHw8Kgt6A049KR5TTPe8VtRyeK21tUX6
oADnjF/jpcuZFns/ko5z9YJvJk1nI+MuLQ8FI5lmG8PyF+0oswp7tEH2f3OEMeFEhH7fOiFH7HGt
DNdDDYge30f0rCecg1uHIMURhfsmYHVeULGVBVskf0CLVeyObVwi6dy+fB5y3IUntPztrE5QDWDQ
vngCS2VKgZobWTXdgAt3wc8mkLTLpfjavRfhc8QZSC/m+BbHhFjehQVIZLQMaI4aiFMJEU+LKnpY
7rm0FWcJSNzdXUHJbIVfUwewnxl4XkUxs/dTBctVMFLujRy8kfQtzea0nxUKmpt+Y+/2NzrVHNSt
3l9C9mNsTyek0LauDkFxBG0mYcsHIKnTWqI5JeeahvZeAV4g9pIb5r9hl3axjWg1v9J5XeoMHTX+
tqat0xUZaUWH7fr7/4tnF13hSx0AdvhwrSa9ceGvyTTYdGLhCa1TV8v4ejjJsitDgqB5FJaAVKVy
T545ek788NsrJju+VvRQTIUC1l1gXYslFYqwcAvRVHUWAHULXzdH2OQ9sv98qPhmU37QKaYydjAW
2SyEOos6MLt0gdam+2bWetQ7+co/An5FyzqfeDCbju+xpnTmDkZxwtClBYt7bwgVoBXtpJPcLbmU
NnXvv2BINaficAhKr5kj1Qw3VhejRA+68RMNdamJsJ5qtA+ule0wGLi+uPiI3dISFv24yn1PYeAq
VyCJSvlKezLsO4KSiTgDOh1Hi9ItnPy5vusYYjc9kz9eqFtdO4TAyeBTC528M/fJt2sj7kyVUrTB
JI2qJvTx+wcNrhyrAAyjF4qPY++dBYfoQtgZkxf6wpSdyieaDkO8rBkDBi0Ij4Nofk4V38SxbvXA
+tqgKM8pR/EqaMceTP+k8tap3q6tga51/Q/3u/sE8fjZuy4KyLBDKBBOZ2RT+OEoLt8BTLS7mAnh
AswF+6Lavn/pabc27SU7Vcupvv5oLYLYuemxdwEsljUN5LQ02dj7Oz68yNeT4FEciTPEQ9zrANJU
jcSWHt/SBCqqSc/ocebieVHabRLMK7ni/hf4wjTBwRqvdPSpk10cHTLBeDdW6/M/AnmHRYhoW7bN
fKWKn4sHDS+90FIZ76yj/a5mVxuHpwyP9eomcEuwVYKDUmpqwCnfFvf1MltKu/Y9XZlfcVDfly+x
SaOdAhp+fphziJcar55ltmaioJlUdbBo+CTM+6pPdPoSQdw2yeVfqFgvxysq5mjSD7jey/q1d5fD
FYOquKaFTce87lLFePrjU8gOcAGA4s1KO2xjWEC78oC8kKVB04/1545S9P5vCLwOcndXaFklmf8W
tzJxL8ITTMsSu6mBK6GCUNJZE0duCJzVu9lZrOOdDXHFeTvE1SaYRL/COaCnNVTFbR1eZlLtN0vB
ih3t+Ha5tcnW/1v3pAyU0dkwW9dNCvhTFoBBDQwXBKY2gWO7soHxg9y6QlOcIz3qU73e/M8tF+si
CENfmBqYnyhdazfkyWusC0nwpJUc+qvkwTNWF7lfJPzy9+ER0qIW+04ALWD5K/iaqFpxkzYB3tFZ
YmSOjtqzLVshSBS6myJksIX8a7sYjv0uxK+vFAhIvJXZ8cVYKzVRDsvurExNJNrHfr4GfzfulPos
yKaDN8rPT+cooM3puVmTKToHiORR09r72qzkQuZ7fqv8f9YPHBEJ1dQooYOhIQgEnRLGFzERq88V
rIz74pAhPvi5oG6G4sOfhK1vQjyjS25afkqyxkNWQSKsTIVr322Hl5qWhkzmJsE5rAr0/8pfbXYy
27tWMgPjkCVvF8HpJK9uGkOVy2hYlVWiCZTqIs8NS7XnQDnG4PNLiop9IsMWLfOZdd3OZqfkpOAD
Ep8PfHMjIkD0za/3ulTg+WFWVG02/VGT2gasc06XZXTeOz84QVbDTNUGFEWpP2YexI+vasLWNyVE
zoIOCN+b24fFhy2W9HyE3i5n8En6JKdMaEbiwC1AZ7tsuR2LIzwXjWpdxQx8dDM8bRZoAEW0FNmd
ytWVtaRzRZW6SyNtlJ69F1lbzVH1QgsSDq/pflR2eLeQxh+R5m6JzQ9YrCgjDcitnN7b38agBU4d
6JHt22G6k7Yzh5a+Tl3Ara5IbSLDVigDeKK+i86Rr5BBhU0d6/XNzupXBzhxtq4Zmj287dRv/YYL
LluySM3UfLNepP176JO6aibLbyA0aDVV6VIaCRbGWHCBq+jzcGDH5UIotwPjtAOgc9HZFM8mtrL9
L2Wq6WEaOnK57tdwTH9slFHnKakYpabxuoAAbusGbqEoQX8drgKRdQiQoavRHjsh0958CXHxc04u
AIA5OYi+1qYaX59ROOnyIBdp5kr7kvEa7LzoM/DOKPS7KoClQJe7Cpy+BMnttnqf1SMyJKPdBbuu
bt3YKVhBOAconFnqS7N+KJLMYVa2IyWiyYJlfXDPRTr/pKvAeuxlhoIA4x5o4aHINAGOgq5KZZFI
eaxlTqbXABxlIAuMfr6GvEpRb3W97QZHsOvUsbfCmc0BIoDqoPTvruP3gNIqMbTeLl/rJvvdcnr8
vHyBe+46nTkn+dBMva7S1V8LAFuGbNIVcK2OqFBiB9yfZjdHHrAwBccyVxKJZecJs3fFNhQXRDu8
PVnM1vIOwowt0lgv9iVxhaC9/zqoXR6j5NX9pK2FoT1wfVI2eCwZkD+ZofvVJwv3MGsQ2hqbYI2Z
VzYDUaMHPQsIH+riyoG/Ag7Qvd7b2ueIS7c8mBUTk93y+X4A9ceqWNU3Y2kHDtfLAsDp5rOBdNtL
xwdl3H5f72fguDsd3eSOtdPiq7WBRv+bJeB4LAQaAsyDAFEJmRYH/iMlcKr5GAcEp7ugN94Kz8EP
k+uJROAO/9Jt1/CJ+QDXnTszV3/6dnByCN2t1MWRifJtLb3VOUuMJhcPmmyuHfE1AJYRTilIWYrl
o992F5uJOTCUM3PwA6DSjrpFBrIZSEGFvRJI1NEwgqhDJNAlaMLF1bOVKn5u5aFLhH8KWSbtwZGH
6BUTMQrayYWmdGh04AlKIEqAdckKKClHXj96lF0WOoGmWdF7KnzgQdQjSC/Vfb+FUIwWNjDSDYUs
d0L+2Ow/mnLQTPUe4h94grPIjsx2ou1NWL4gnUDNr7g99PXpB4rt/a8PaBNnGlupoJHHNdqRYXsY
4qamwo+sbNVIAi3t8BE8Nzcl496JSHZsdq+tnh2P1Sa1+2C+o6HYlT4DrQiavHmojf9H/VEfFtNj
yoKt0ASABRMpmSGZMm17NpGvMer5YnAXfcFPqNHYetTuum2KTgXrQkHedSRHVBjYAsTTs4SKq8Cq
dhTHvZ1hGZA/fI7IkZtEyhmd8IKXQ7wpCZkWWIm1mOgguf0UStY4UfmrEFUqPkaSaczyafTjZ6Bg
itNXITcANzfO+kneZAggb//gsZ6lZi0LtgKbY5yivjIWBvDnto4Zs0I22Jjhi+GDV4Gr4Zrlj9YF
tie0sGRMfC7tLdHS5RAfYI9y9gTBAez8JWD9gafMlrSUxSG9XjdAYtXbroxJbCgGEQ3XuAQ6vdAP
mmI2eQhfj2dbYB/zRkDGo+GusnGaoMOL/HwdKcUl2+g49/Kjn33/5qsFGLuXuDrCIbiGNZ+LXcXV
2cGhsbHgoYKn4BZRvB7Vrm20xrW++Q/Y9HcFgOE/SDuxybdfmvMpT+nI3eT/QdK1A7jWFlfrJ2FW
Mevt4kZyUhQUf9NAM6PrDNPrs5lze4Hxnswnr4aerD8c6hZAxEe0K5lc9nsRUwCWKPd/UI8r+uq0
wLdTLVC2ZJQQYC9EZoqA4NzfPSedMvVgXrWvo/7zsB+j9VLeB6Bx8it7M4nCPc1Nvp02RrVkAJ/+
PDFQEuO7DGV0sXVUM+AtJhwajKymzF9D8g5sCOyXQncUj51+TWmqY+n+/9T2hLusm0hxIoMnUQbp
yId/1/hKb/xgVHswxcY+4YajsaeUWjmD6c06ePu78GWmhAF7uLl0WCmkTD+3pKR67IKCX4qlJqin
7aJMLFdNbVeoCE91Qi7IpK2TLD90G/TD2UD5Vz2QXyfEWph1vIqTXNc8ZpoIZiOpBZMvTCadoiWz
AIztg2bgjhlyZmSbu7YkUxecOAGknqE7ZMdaeU7kXqUkalsl05kBxB+gWY+ZPNfqvvabTLYHV3An
dQ4B8QmHhKuMaHiCB6nY/pe3Rm5hv+GuJoBGQxammYVvGxF2+PGi17HuPwEHV6HGY/ctUVPokTSg
xNwQkm7keuUiOakvBxPpg5a96iNfiWKxD8LVatsT3TdcASebpJhz0Ci6n0Cx3uwN7H1rYPStMKZZ
vHnxelwMp/m5I5qlU27YkwxkrjDKbS0HccsiQ0jwdBI4Na2bQuCPIt7q8bxU67S/oxn4eFDJcOFu
jPK1X24nEZc6UVzVGK+2ararzGJeWtLPxZ7ziNRsaF1oQo/iYjUDga34mHt5iCVYyZsuS4utchn4
GvSV5cnQUV5QQfKxQ6x/S/KUOWcU7t296zno9v4iTj3PgaGWm3InW/Q7gCiqOfvtAPOMiQl0gVX2
VIWA2Hp5kXie7Mh4ecdEpb+YnzUY+rv0jtVA6jcC0bc3GupviH3A3Ujt1MkYa/JRFCklblPoQQAl
ge27VQql9HWTeaDvveUJ4kNB84b2n/BffKP489EEDKyJRe2RD4AD+r6yY0mDlF2F2EkUnZkAvUyK
pRdB6Gx4FSrEolKksG4pTg55rvwJi1ELcB0PdVOVHvvK51rJIbJMvfe5a5aT7foB5GJl6zjizVFI
0K1sUbpWJCnRItBZDpCiu3bhSxiadST+56fFKj84Qwh7vKob151+wBbb7VCMiFFVB41JrRgjo6pX
TcqokzOD4pI18GJ9UCuE3t4N8tjwbfj1tPVAMfNQGPQhIu6XT9qF2xJ2BIqY5dmgq+lmNKlViHgX
RSx//CkPm3GWMXPUyy1H7XvnGHpNY5wYTRfkGRzzrkEw93aS17tJaHrks/9l6hOPL5xTWDNX99cx
4rtbKGUq3eChcB1E2sMIwCjQ6BCg9DTTddTIAVe/VrqwPxkKgTm9JZFp9BTrEnc2EYGDygrzVuFC
+iCi8YXQs16PFDKkekqTh16YUq4BKqKxLQnabFhF+x7LUbNcoVghlLx5/GgVPZbscqQfVc2DTKuE
M3aZLK6Mgex6HcYMkkNHM7jMaE2pw5PFdALKCGpT3aLCUOw2iwrSrps93l7ztIacZHzBbT/pbfVs
VCU7A86bbMtuejrUwVxpjPk8MOyC2GyRY3HGhKL9QRg/6wgaDcZnFj2UoOgE2YkBp2FWvYZhoAo2
Y9UWexYOeiytY1Zqm1YiUrEAFueDzyEjSiRZkThlxDO3DTBTt4d/SCotpM6mRxum0yNTe6S5gh8g
ajHrQ7Ma6nFYKN4S7ozOS+AvmzAVYk4aISEdc9EqTbVyWNlYPlBmT6/q+cLSicjeCVw9pOi/KEL+
LlTBKZXPiV6o6e/0VvbYncrDM5WfnAk6xJ9QtEcyHIbYRkhZkuMsf2Nwcg0ioc6KNDZh3wopz+6l
ZiKLA7mmnVrF4aSKUhrrIX50MoIqFmHPgDeoYWgCNMJDIKxMK5NNGeCd82Qr/cx1BPLoDY1pswG1
6iVu/h72veRLbg5yGRZuqxsYqgZvlBr0+44vDlHqlRJiug00uge0ZFyzFjXSWkiSPbIjeiEnjOsi
O453hLUqSSb1+t1kIxXhS0g6aH3RXY9C7L1Xt7Rw1vj4I1wMsdKK+NsapGIHO38H7iHjyT9Hy07A
aiZ89lF2Z+w04IWJGG7Dgxv7MJLBsVHtnP6SrYaCHP4lq0BrHBZKMBJz6AfuofYK3UrWhie9Ohla
Ie0WofD7gAmCAt+k60OKBoOhfV4djFOEiyYB0d4OZrKa/Z1YWsXIoKMMUr9u/R4ZVUZWXSDi7gnR
NREybRZv0Q1ja05YTB2/MWQVK20y59syu8VsuyOV9vfMnpaY+ZpQwt/1VzMhGUK8pBR0V5A6nAto
bROCe2sGIG4iPbzu3L5p8vl9F1qqN3FCktRUWqQM6YqpmZL2dm6kOIvJ0qVLMWMJmNdJQIXVy2l5
x4OjnMqj0poIT6M5XD4YV82u0LkaIf+ag1XYVt+2nLAkRtrZhaoalcXqGyqjwmkXFQYplAZkaJXJ
8FcIMtzo0fcKx8xaP65UWfN2xEMiuj9N8OK06zczftf2Wv7xr3yo/MFEuFLOhT4aQOw8RmuWKQj3
iUaj/6ACwfUsgNhWwYGT+H785EyajIAT8llFdWsHqP6LIJh2MGdEBAJbUt8oqFn/mNLyxflmlW20
+BT+jFmDk5k1nD5HzucFr91SIXHXphoe9iloI8XTQlu0RI1iNJgny5DHzv1IIOi+2SNpREbxKpZF
0PGNaO5Vac0kIsWBODfUiUN0HD3j4/Z0Xi3y11PPo/kZlxeQrnn0nikN2QZ7MYFv9qMXzN2vS+Kr
WrU4SNU5b79ageoaT+PWdjrxqXZW2bECYgUknpOdVq4FgyRldDQs/WnmJi6uLLoeAvZyhGwibCsU
gxMtm4Smbi/Mu5vLFi33LEyrZfJpTDi/yFgaRlN5YZwlRaWj30o9VTcPt3gOoCx5gdX4IQuZK29Z
j0D5r6o2ZOHquXiKLwosCm60NPYxE2WDNGxEqWdmRP4wg+G4mLORJ97wnIapNrSNX1uHleRLVLpb
qLFhrcB9b5mk6G1sfZTQu4HJq0qkcLusBVqE+r+5UbkDwLjIbn4ViMOt8nSOGnibLAoGy8UTSIYS
MognRiNLzlKyxf8EWeYdJYiTs3ItLLgd5RFbtkQbcV4vs0RkVPNCFBSrTVIP3C5yKFSaNuBYE/wT
9XLtHBLdmPzOFwLhQ4zl7weJ+mpQengjZUKX9DaNdi0TSfFI9zjLBDjYf7Ls8oAcokiLL/AR7l+O
GLX9tz1iTRIgfBtW4GLftJcx4Q1mw75wSBtYjYAKJLbTnHUoN+dJxfX6srU2a2ifEv7lWbPEUbbG
4ocppEOZ0opz6KLBku2BximJD5t3uJh8na5ODoav4HCwtblFzlpXhuclLYALXw9JpmMpFG7U/8ew
5nUllK7B97D3+Y+ha2lqhUbVz8rxXNcj1dKBQ+WU+kUOHP5iFq/jpuv5N3UhdAKsw2A93bt//OsL
RqrLmCwAa5aSUtTeMB/XLNNB+ziPb5rNl8vo22lv+Buw+mPJo0AbiyMExIvR1SmXIx4vCw8K2GBQ
q49C0JOZldF6svLNn4c6cDmWneAsluQeBwabV5hRsitXUya7qHkcuFjgLHXlgdz/qAhUHP3xP2Py
Ls5UL6/QWz2CMiVIaYSEj8566Y0XZxy03LaL/5kf7cgr36I6jSsaw6iWFsxoFaPeKKwHrKih4mid
45gwfSOVsaAvBH0vStwP2/1D9S6O6VeCY/udkUdn4PEXlK+PzpARH4cH/vVDKAl5DA0e5LV1R0Oj
roRCFxQb6Purw4rMHmw1OT9X99J7bQSQOMkXuIcWkWSB8A0hJhOcbs/fk7XVVzi8c/ATLlqVYH0p
xOmnF17d1LeTqk2gJK6C0ESxiVOCWiMSYJGlSeVQvRdW/V/FSMYuVuXc3+wcZX1Y8FXd1oUVFyip
hWPrZuL7Hd5uzZZIrgCGALnPyOBudXsgyNY5owNaafFbw7+//YF/EXGvv/W2z/+UWvYSTba53Shm
OR1haFiqT+msc+S+l6uX5Mj9TvLmwhqQ5l7cdnNvrzQpFqAL0DvHX7YKKuv7QhwtFPQp7bLMLut+
ZxEZNW7p6ezGoKmvYNYZeZN2MlSZr6YoHSfpJBWYOfnwptOw/tFnV7WJNYSmLqXYZO07wX63UcxR
e1qZLSGhTeKebSX1TkLt2Op+qX2/udKaLDsL4COQxWQHwfZ0K1TbXO9hWMT7rL7etFTjEbxn/RHm
iXbkzUIjncVFEKn8zBrTH/6unMO8F6PBec5yAimHNQQBc0TPLHvEfUog8DRxmlQFCSz/8QTTazW6
FASwypQrF1fucVtUk/RzR6/CcpaWnIaLGvSVruuPUrLATo+ediE/2Us5NqyA6Wh50cesypUZlGgI
wyxl7Y3P8NfBuRPHNZIj9yA7cgFUAJx9H6/FKsrvDfQycEtSJ8owsAW6/nZcHzU/R718QTxn9Xbm
KQtr6iD3fQss3Z+kZMPS9JSrS7iNrhzHn5zL9OMCZpgqHTS2t/uOEtkCylCMtLbPD3wE0m9UezMA
n6Uwaxy6XixuYa6aDSQbV0fWVMD9k+4Fe7baG8s2bXCFEiJUMKU4jY997HOh2nXYOxdc4Pjq28fd
w1TBC4h184AjhrO9hESEH8cdnNZDep72nEmfnt5uVK4npsjWLaiGinhcHok7xNfQT+sH2WJ8HqGV
wGQ1yMFUWJgUVPNGo7tS0uE5j6KBrid4lC3DtwZKtmMzH4kq0RhiM0d9ms56kwi06r0XHFk1hvAK
xXcWTMmwlTxrMgjyZFUchyaLVwKrpypVRSJS/Z5bKlxoV67ssyEBF8UTszKVTYnE/6tXekrmXFnL
aFZr6RP2VRUpWr+q/VAKpdvrQOK6l4nCow53rig3QdcAmpRTXEjZEBf6tMMZ0NSawr3rCX1Juhv9
crV8lWgD5Olort++mvjJ1kekpURVmucg1i8kqzfEBZdGfyx/6r9C4esdoNMgmSnczYilYT++JCyh
hXLti+3z1LMCrIVXKu0wInnCgwNsLxf1Xm97ieX0oNBx60CXqJ7Agv2MVy0mqC0NgJrv6+wCMX27
WE8lRP6uZToE3LC+5DMN3NyniC/CApWW9bHkeeYq+kLOl5QL4qdRkRFvRXnD5WczdXdbp0SiPzQZ
e9zQMC+4CxR9OKw+iqYyxSkwL/wrWjVpZO5U5V2RgY5UN2UQT6AeAmZ/dbbK9hawX36bGVFHZT3t
2JiNl85gexD8xZBZc5FS0ZGPZdi6wUDtvlMeBKDzVaMHgacLPZkX6H/W1S60MxKDaewr848dc0AK
UBFOcTBpkzPNLHdLiWBAbQgWkae9tIrhXNSIY4Z3+MiXI292r357slj1M7xIL+S0katTz/fIPBrs
wwB5VbNjVFCOjMeS+zoKVDQGQTyjjR7YGWVqqcVWYGLGWwNzk8aziSz+Elr1kXBURVWJOM78PUTk
wRDQrrAUkyXKn2b1D+h1eRUJ7Qy17XAzK4AYQyqvSzNKmiVR0cmTOFpK7CAJrP7NJAtjcAO438eK
ieqx2hCU7+p6s9jDCcRX93Xy+RT9r0mfBNPu9GWFHZdcLqF3h6oS+QmZX/rtJUMGBfOpUf1ymCwu
pYMpIh/KPkO7t2g0BLxsnxWZBlQdePX04ehYJzYq9myrKDfapIpHe0NsycgCrSC/KVGyBalAvlua
L+oWXU0q/X0UBw2CA1hNLPXDTRTDcnSsWhz/FnOEBfR1SfeKTU/2QdgodwnYM3SBK9Rx46Bhqxvu
cDgkhph90tDSj002zTQ2NGxpvsGCMPnYTDQGXyky4q9DXvyHK0qxH6O2uZMPqkPw0hwg1S9pGojE
f+apHPQ/qb2YzFof+FHQeBfDTjNE0Q4YdMM1Dtw6M5tyLJsQjtz/Hse3hqVqlj0K1V7bohkfLtIm
JS+ddW1Unks1ez3J2WdV4aQU96m5kfiVRSZOfprINy0j6N/WGN29i4GOaqFh1rZa6kjzjR2Qe4gh
0c5TYImYUaqvmveQZ73TPYK9jpedDVttBSgbF9v72fBRvie0RddgBq/rg19UE7bee+xralg/prwR
c6sG9hhP7Lny730GIKBMd5zxwAMKHTKaSP+F4neopo5MHGyc29Zpyy6XICPrBFFkJrtTWJC2n9w0
1qCeKS3s7h8ri9oqaiLbldwVqWLP+cb4Nxqlghmw3zDwLuRpf7bmFbP5+EHwTLlWPGjmZVHrVGXV
bRP3Ip225DK4iucEG/oR2OxUTe+3rkxn1gfgg0DZ1ilx0DghaRgIsH1QrmbBc+SxHlVDnk5zaEKf
EI4V+ZyMxq32oGa4xSulXDUozp6o3jqiGlChiwp8i02QkTSDVTNOe+Zu0+qOXmMX1lxXVSMJT9u3
RX1BZckpnq203lTCK8/gAT0JGgTYUVYY/hhiAgqi7nIzLzeARHOIm9oIq9/l6Rzm3SJS6RrYwUzh
Flk2oS6TC/Hh57LZ8a7zy3WqF5xHSOEhBIZtfDeade56k0pLIG3znjz+zDyDiyNv48gDd8Gf0uks
wYbQXOPrw9UEvMZahmukyPXdE4tX9jCVKAEqvPyzVUr1ZeLD4+6ULBbeZAU0o4jaRrpJrLjxMK9h
qWiMPNi+72+QsjfI5qMkmgMqYBcdN250wbngFWw5SOP9/8CABpCjggBjpV6guZkVNhS/MvYN0eRI
z6esUkLv5fWNIQafoNN33Cl5nVk2yurYXFvyqaDFTz4EZ0i1pxN0ysawMG5e7AKKcOPiFyoBVjhk
64b0ZmHk/wkV9iWhlY29cChwDRTpe0Ma8rbskyMi5rHkO7txWBW1HVyuYrPGch7fC1HK6GgFWu//
cIZEpKsQaGOKg4Dog/Wi4vfuQAS5/FReHpGqwZsy6+bEeYi14ZJ20L3SgbIHPMyEWDsbpR0IGxoq
XJK3lHahARQGVWRBz3cdB+ZuoD5qLSOiftpyhkrNb+Vb74fPWxXrrer8ybMvsk21aeAf2smz3oY+
G3GMrVxmjpZIwtxLYNoX1/RxpxrsDeMzZD2KK3kUQfbwMpmYrMYkx52YejRCvPWntu34pJ55m1yr
5KyfSftIyXh+TjLmzJESAjJo9Tvm1VjylxXmwQUKDWhpKlOytOjQvW2BJW7gEEf32UQj4ET+UN3a
2RGbtxTFefZ98VpT39t0Yq26h5uAKTXyrr9T1KPtQbi1n7ri2aIjDQPyMKOltcPT1qfs3HGSfIQz
nHu4nKAfGGx93wpDCgU2/VDfuSwMbBgEwDC1QlCne9u8/F90NQmZcpMWOFuIWYa3Piu82PcqK5Iy
khYLltc/y7wUvKTWO9QM80xpzEQnEQwaDQ8Ar4qPiGoiF8NK45mQOWMfDnlg6FIOH2K01DmcdJp9
MI0z6akqjAAQFbpzuFESbyp4x7uMM/pF/ZOJmgLWPxeXh0U534aMcsbC7OAxqdkpLf2Bef1MrXD7
/25Gu0urng1YBzgnqBLx/1Tp401AMQnX/JcF4Hurp1Ez/wHYCmJR7L+xexAF1sJrscMPhLfA6IQ7
l5oCH0eArNIoy3PxPBQ2CeWnO2SwRvtHrju4XpJACkoL3ZieJTPC7huk/EUwm/oDzqHnbxTLnEEa
J701N2Ug0HQPNTna5+wcKEX8vUqlBBVliHyjPt41EHM6YxMugPYnoamA9QD6B6gmlvyaKkRGhj/C
D8/aZuC7Vo3k0ZaKA299dRk97kCVeYazJ7+5OGgwBcHps3rZpSxAr8AVvflPDtuiofbUUeKUgNGK
nsI3oS4uPFqHxaTWgIqy812tu8QmRFVuqI/3jQneIjuhoZy6YllRxO1psyElHIix1kGmNa6nq9zZ
qE9ZBJyUv673kezYU3hftxdxcRAhOgKmbBjGbLQWtVxIFHAGxhekOwv8K+KBn1HNUQdtnu0nBjbJ
bcsq/7h0jjzZQTj2pOZoxIKZ7WoC5rYPXZOFCv/39OjsH9/lfbYg/8yMylrAfgAi5/Q+bRAt6NKu
QtMf9stsKsOOmML/BrXZF26yEwQO0ZuTQb0984hVwkPD2SbvyHFyIy45UzV1coXHuT2bDnSOkpBi
VD8ZSp4bIWVOs1XUYtmbDy99Sl8qQDdx33rnIcdOFRE2HvkyYf/BbnB0kXPthDg1fjDZPSyK8F81
ZyUlau3QOBR/CPbsmtN7R8eZb+gJnE69UPEgc3ApbUGdULn7MEzpOdEGbiVomlropalz4mKsThql
T5BqviIsiK6dUjJYC1TYS+JlSPPPc+P4J11pAw8J2Kpoww4aoRrD41Li4JFNd1td8xPmph35CBpN
+8KR+vYLJ8aSQHi/C3GkA0iC5AKTqV0yr+cIpYSPUX9kSjf4ncRCgIcIFOsh3G3JOenaOi47sF9Y
2NqgJ0Q2/5MIWECVTm3r2Ad8or45RfUsEibkggdeSleR7XyBVm/Jebr54n8bfUhm8qlVwsQ9sCmO
io57bgzxAC7a+sNm4VDSTIhBt28+vnIUG34uHFLODHTjZI1HuQErP3Ym1HqGw5H77eToBbSD8YyL
qsLUEc2UDgvkR/9fQzYvx5pwt43ffsiO7Q9zN4vC4x5aDOdofNIX6wDkNVk8jSkTTFrjKzfY22xj
T2TGG0rp3iU9z+6lMHXyW4nF54Me84/K0rFiY0KR8tMbCIW+N4C7bMUAFSlO/HQmAUXoVd9wlBvN
+Bv7zpdfwfZiJDUqRbPAKf4C70/tdCg4AucJ5doIsNMkWs23TDtu+vK6kiKup25sHtow37voAkqZ
tEiJxha9c4bKf9U4IkHUZMtJ0eUPzhQeGH51o0W2dspnwT7XmJdwEmazaw3mLhImy9rAURvZvl7E
FzfPXnG4Kk1BLcjKXLjSBpHxkLzuBtzypUL82lSouX2bxh+QIeD8Kntx2K2rAPVe3QdNYrT2K59Y
xwuYaylP7+wY0blhcqQ/XRfmeGTWA6jilVYJ62DKjfWWdEwiN57Y6OG7YqVz1fJsxu7fzcNtIcg7
YTigTZJ06AEoKK5fgtDYk9mrtSTncgJYDQ6lKl23n60MXZqWoxSouext7OYI3r7tbqFAAf9il0QT
ayK4uqY2EOIaAl4aRAGYjrthKAOlMru+NVrH/V9IEM5tV+KKwsjINLgjn8Dlk6R0mfzi+BgZS+ub
AiMp7xGhSgEP+8k2f5rm5irDwNkKh4FDzr/7QtJLhXSwR00+kvWH//ZoVOG30XDX2F0CZjX0vznF
VHbpXZ36MEatcWVdk74Q0SHXeigg4ROMG5sf11LGFTmwgSXtMBzvA0//mQwpj7kNH62p3AdS+Ez2
EOsLX+OkJGdiRvI1wgu9ASEsQJSIoovE8prnYe7BRfG/q9NUG+AFl6CsnHSP5EG5qJpUXLda9xSQ
bKROEeQ3GkQFEfo5bh7wTXgcc+DOM/7BjFfzJeQp5r7N75X17+MEY1wH5Zr7GRDXPE5lgRJanxOV
Q4nwZKdYGxmUMtKs/1g4Jimf6YVIvF1d4LSPdc3wvvHxipxN4TPXP5eIOkb9Cr93G9uJzE+ozxX5
dZZGQTUSxqqplDHfWHWVMJMoB0AFtxk9a3wggtCojtp01ZPg0J2fObJjNWK2q+L6HA1MHdp7O5Cy
Zt3T9ZT/+Z0X+rK/UADKQpGSWZicKdahmAYl927+OhfVgq/f5LfnV6ciIcF8A64R2DFvaLJOKazK
6OSm6OFCjKuKNxu0I02sZkE4XKZeSij82RzwQn6984aDgxIzS2L07LinyJMORK4GEtQSmhMrlJmA
phHntKFBds6dS0PiKFu71W5Kbk6HIsyBlWWcxkYmHa1s0Dy4UFYs8VpqsbEq4QAdcyTuy87bP/F6
kq3zsSI13hbz2nljH5Gy4RxDl7ZJJuvWz4rLUZfcdFgigQ0fS8LGM6AYIEvoBghAbNtRkpjjQ0/9
4Ry0zIQw6q7h1OqUWlQxWqz34Rq7bY3X+U2ifR4V0n5/gn1yKRJl+lSKcpo5nw77gVjrLM/ZrzLB
KALa120WLxmQ7cXBhsidGrDwEPfg41LyaUh+hbMJwvPqhHPuIogKLGzkanVmzxwQyXLwBUcLjAyh
pCpKDeBGXG58C9vYTdoV75hHL0QOdsYHwzumEFbPkf1q1cLW7WByrsZe9xrd/yZyiMatOfu9wvSC
y6r6W0dmYYiE6qyiSLFbwdSd+wLrVplHo1If69o0sBV+r+vsMK0EuLGEZHCG9HXicP+WCa6JZrmq
S3gX7g/kwJ5f3SBrbI9z3NlUSjM+6Sqmd33ctENnopHIbxGn9x5gpJ9NGH/Ek0dXxaahUXAwJDUT
XsdpZyGFeHUBAS+JIeBrAfV7bjabYA2cIkMJ5f3DNn/aZcxUZyYWEN46Z1K+uxI1i7gya1yZo1GP
bi5hAKWCehbjoZx9HU4EMFClJ8RkfgsXXnJWAZS8Ji1AEgwxh1FCw7lqUKTV90s1dWORvk3V096j
6Ezp6vG++JHrZYSUMvvnJR5WF5Cd5anc5wcovEBa9mJi8xyeYqF/dP3BsGVu0hXykaXAyav2TJG7
5fbP8YU7gKI01pak0wvtXKnnffWNnLWiqS6l9Cd09RA0wHimCkww9kSIFGumAR0OIGzEmdQtJp5G
9Vj+62wQ3U/fgt9xm9yGTKYYJ6NZXX/W5eY6O2Aq2RzniZJLovrxeIeLjQlrx4jadH8nrmcMZMXn
hxkhAId+VJQDKvytytmIUDbLQZLWEaP1fBH60BL/RbMjtfS2k0P+OQs7O6CmGIOOupFc13lL3z4l
Ia/woLyLFCGNg9Dy8lkE9WUGxc0gMwIWBW1uX4396kcIvyp1xc+q/u28IZgQc6L2UCztVWNnA3O3
8uM/qXeQ03h0tuSrvt9XWnAKkddJNS+CKn8OXrl1OXVf8BlUIdVrk2XlUi7tJD9LGdZomvfcXkx1
0VjcshAoRmxmuKAbgA070DLGxz2GkIyqXolp0Qs+SrDJUap4MQM8uBzRTrsnR9KLb0pH3LToFu7w
d4AuheIL2F20E2PgkpzsYlW/oqjSFLHheURYA+6r7NzREL+3zkskUyIGtLvDS5ep6u53J+HULsz1
X677tlLEuTJZw4cXYjG4N1o/v8auPIGuo9yWTn0n9xwjN98v4g+NdqVb56mRgWg0jibHMNV8C2RO
2A8X3WfzdIYuljm+pFPn32OKzWE1c2kkaWYhxM1Om8okUR8gQx3btMV0mZ0FnNcsEB+b7lxRxKXJ
JcOZQKwI7cRdq9cFKmCbsVztq7190Ey6a/n8YKTGALYYe4iXAVgkAXlRgRLd+u6G7yTtQ/PizsVv
uJiuQLOHFlGJeWwhRTP9gFdbtiEIOt/0al9UcCEfngLkWYtqCJmTyUL1QgEwGfq1gQ7NLOTrxwvk
87W4MAXRW+no0BoD2I2cA2VsOtWYMAH9PIhCBzJ8CpIOxTrpn1DaU3ba3eCpAEenFu3YtvoxAsXr
AGti3n4UqcwDAuB27qK0Vq3KBljOiOQTF7pyPtGfLR9SSyRYQmTunPsWlxft2ZncZ/IoytvnxO2/
n5hqc/3X2D3cG+0LVos0ZEk7y7xFrNUHHzvRvFAfaXKnjxF7bzQcynkqyBP00hziOb1YJZ47qtCq
GHLXC59YQOXDdkhQfhKYyRg82GXu+uML/x0Gpm3i2zP1jVhV4MgEXQnIxmpn848hQklRx5LZFH30
TIA5R+GgRGvA9TcxvlTLl1ffSOSgcixNmsBc5EkXEW8OFSMWM8M6wTReIowmOGZjZxerzulksBZO
tmqFIwWmDYp7N0xiIXFFze3UluYNpiJybJQVNOyZnk4LktRngX+fjEBpRsGirHvmcn2EcUmM+CQB
Q1MNFThAhonJug4Qxj12B1lS0aETNE2ULa5M3toQN2riegKTuy25P2qzFKBUVBR1eOvvPTrSRIfY
nM0Ve1GwvqkCqSh7Vzn6on/vYrIbv/xfCQY6iEx55QwhgRfelimUnVMiIGLu5OI5n14kF+SWeCPe
OXnkdqQ9ZeXXGNYnt/xTo3+o0Ob0LYuNKCZDlvkrm3SEC9qOKcmtth1lVfkob0jMbqQDF1oi4dIM
Ij8PpXSgc2I4Hqru9Avbjk/TY2g8O5hwEuNcUCA271WNYyxy3upd0TPen6yMNNvWnkFem4geIImL
I3IeuaeTWmWvF5IqKPYAY/bpoX8rpAQ246bJmiWYfOpxcYkD1+vyb40s4JQaXHTzzTabdz7oESAS
bMCGOjE6KpsLBByoL9+pIjcJHf7gDdkbPTLFLXzgbXOm1pawUFyWH7QTcTFCzhMtBUYJPwwF3fLF
zn6dDn+mRj0JBAeMznqKLN2I5L0BqjcXyVda5DiFah79OnjKRO/pfd8kFJRrJv3D917pXL5kcsrv
Em75jzLqmMe4S1mvfxrKZlk3LJh0FuHfWD93IZ0eJI4jTEBt2WMlCU6xAD+kuKQs3f1ux756eowW
TZWg+Bxg5AnIQJp+jYvH5ga7CQhV68qxtyzEsnO50x59zLEjFWECFHPpB4kQzOyGG8890Mv5BkkM
xGUNLRc0pG00P6r1yxIIDiGE6zEEFDVGXtGIxxA/J1/isPZgE4G5kaX4Hgit7drjS69RZ6a/k1RA
6N9HY7LhueoVWRvsdZqh9OzjxLjznluSAaDduP3d+xBOmUwoFEBhIdTlLVOzuZrgqUIV+RMLxU9D
qHKrsRtyNnGgEGN4GQM3uI0jr/3J96NVB98K8fu9nigx8dZx9P9N7a3BzPjPA0JrWUrubGy2qCVQ
cWy5H8bAeMLW2WjSvUl5dLwvFVwY2ac7ElNAp6TOpMq+YVbvUJcMg2JRzWn+Iwl6toUD7s4P6taf
LV2t6cVfT0NdC/GwBk7KzQpSWGdgiPauXtVGZzVBFiWEORGGqtdQ0nVWVsQbshu4TXph5017LcP8
+2q7X3BwGmrV6Sm/VwUbj1WHwGicZmJVa0n/YaCvAF9AmrAQRTyoIKIpVVi3IwmhqOLpfyR/sDIJ
DW1MLQyhP778FjbljfhNXr+wSTNj0NBPpMZATCEJ0V2M6THkmplYZFZPJu3JBUa9mhiqYj0CC2st
4G6Zmed9HBmp6s7p5ONZ0gbv7XTNmi0RCRIAtUMC0P2ZzQA4Sj+4k9L6tZAbczOZb/QNTaKORzpm
dDX1/UURMjXYYzbL39FbYS7rY9O94AWlnBMoIfJPL2266nSKl7GNdKCQEYjTTlbnq0VvOu53mZq/
yzkkSuTqPF9xdiRrUXFSHBpIlGIXHneMapdHalLpUYSlJSmseGwtKm4uLNqJE8WDwhsBmUDQOqwx
OIXUxifIAJwXVni502T4W0m+CPnpkgLGTJXjhVfQiSy9/kXaOy5Msx9Fjhb3TT2rckznpy98VMDw
q12QP+zKQBBAHZ5Hi68BNVWOiowsRpz7NBGt6p8/eVzdtB0Wi6a8xrdfL+Y56SEkRPk0n/wleSdc
ZpmuP7o5MZQVmaGnkZlfkWHFDY17qHbSC5l3yPN3hG+s8Q+t4JtTcFVfrPfJZWZYEtQmeXVy476v
7ZUEoN9Ov5zVCM3CqJOHNsFzD285iBlLqVjyDFtpcl9aVX8G10TIQ4iGo5FcN4OIcReQRBZf31ks
YAsPqM9Wan0or5/2cpq6Ox2lSBJOPdK7D2eGh9b9hv69fWq1fUuWhWPVsXRR8d7MH/HKrF9Jcji0
gO1FA/JYd3wJ+AMJbZdlG00ejwKJjQO8f87vHjXqSQSANmfBlUhk8Z7J5Z635u0fdSt/3Z5KpTdL
TnyEpAK/W0mgMzHgorGTF7wMuvlrJBlMLuB7PbCrYw5F1bBVuv249lq6/+XPImVBwIMcQl2z3EwB
drmjWexHYOf0/xOkVmLAeM8aex0c7yn0HBwFHlf6W674LxT0KoTCAgssk6ZZuLNYM5LhIW7kS+Vt
9u/QgdyLtbxrmrKa0x4QGTeFAPJm0mS0wqUVwrNdwGfhLtojMM64iMdXcD7A8b8QHhHx40dwP2G2
I4FW7rvVw+cqHfmcwFDC4WMZru0DyRZlTWGZDve2HgC6GPwLmHVgzgtX05sdWQbPpx43zSE8tXxA
B2KOKslMiDKsnYDijKJy02fnN/LpWJ5Z1wrnAXqLshJYxbe8uLdUiKIEzV3XxUJRJeRguqTYQ3Dk
vqbtSHn/al+aRcK/D+3NcAv/iOJTbAjzT/UQUd7Vs9EBkzpZUb1I2bFrDC6ZESQIznnlE65wzuXG
Tbc0nbd3eWivo/zjMDsPAL2viMRF9LiZAT2gFEWDJ2+wKrfTMKJzHoPm/qQF6+3ZQezhokuPjm4D
cttjYUOPUVVe4FqUl8ddITPNBwor0myYSMFGf8cwjrFKW20139FUs3np4TcRjVAuVotYZCdSeBOY
2pDKIRdIWQVzjasXVr4CV2cu71TqVlBYL991PCQ2CGduNvV+rrR0yqlAbPxQl93yZa5Vkp/v2Rrt
EJoaZl3eQELeQ7R31N9KwJfIoyUP0WwybsHAP3+O6swwoVFcAZoe8CNkYPJxvL8aE0vgpfKbWhEG
k8TS93dDzmNdO0dsrGa0/yKH0CBQwamXbA4Mom2suDKtZXFb7otT7FZEuYynHaE3RMKcedKfUdXa
MLqOZUL7Ofl6IoK70IXVLzCAh2mEgLpMUoDhNCBJjy7dKgG2w7osHY6Gcyr3lKhwtgoVBzS7Wihd
OXaigvss9HbYPKsajSg42sN6dWbmZilLAGuH+0778CCjhXOMxE7idCNJX/LbaizDFiwkKKardmc5
3+1O3A4XKMV/HiqkpFr8w41cQULhGdn/apGnGPaVLdRYTsrg2gn6oMhBjll4GkWdO6TKOBsrldk7
EGEN+3jM/NnBpX8BY/FZM2YrCvj0JOftzVm5CCtvBS/n0UgrP7zdS2YwkeZMdFtPL3O/aMRr0fdd
lJnevClgZPHeCkmZvcGDSAjzvXzjTUf9KGrr48ZsFZ2xWn81Y3pdYxzc00bSxMp3nEGZhQUQk4rr
ajGWv09LKW+mNfBrBpWFMhG1VGWlmJuzcuhU7ukCNhG31PyxESZSUMeOtwkYYLN7DUxwW45WSsDO
gWO9w/SuLsv57l2Cf8Hq2utdxRo4hwNXmleu9azDvnBNQ67NMxhEbLRMPSclUrt9OJwPjO6POzjb
aUDbiJTqK27E+VRVlxb7a3NSwFXULF6yoogP/qvLXfyFB5E/Wdug2a48v+9azoOUSEZaN0CZN1lc
8qq6HbR+zui3zEQm1ygr1rjHmxALK7NILil1ZrAw8ddFWoKX60hIVlfl+PkXaQS5VMgiLLkPPtj+
cKh0PzQH9j8dp2fm75XDGn5jGDMH49dPUCmFZgaepnBYRHoQ/zQbZRgSVJ/v4LTgn6docEUr94tL
jbKLgLOtK9EB74L2/9I4aFxZsCtHMCm+VAeihhvp4+s6WFCEKTSU73HdqJ+sGk+G22iChLTNoQsb
spQeYRfxVP9bYr1GSNq5TRELRbwJjffiCTo2P37SlGYF9UkauAnhpi4GylBdeI0+yLup4AcrSDIT
Fz9Ax1aMy9t3uT7MdKRFmu7iE3ZyQQ+HUvbmE2glM++V/oyAzSH7UqlOKSY8RO4cKJluyO+lKMmJ
7o2ToLZpYim7B44LwVk/ISMEdxJ+F1aIEC9Why3/WvLYCUJKEHD4CGb+byAVvUUD+dd/OsFRpgAl
hlDGg6BzTfJ7c+qeymm0PN1Z0evf1B2OTil0xZ0dYEquzXv/P4SlYpbPwqmyOA0gCqH01CvjPlmH
YcRPm7STVYtd/k4J6Yh22mnixl+LOOFWYLh5rFVTSCkpe37dgEmxpIfQadz2klTQ0cCpfXl3tlh1
VK9XvQfaRujbbZ4rp8bBzTtVEUqD/xx5wuoeBa+aCLuPNd2ImtDKZHdC9WdqTIoMIgQFcoiynRu1
olKw7VPECTsd0qeMduoYCEuM6Tsu7BHCo7DIUv3eDjuLfPkE7wxmC4/hCYOhZTGueyZjsZqpK0kb
G51f9WTk7HBTK5b4CDGm0CS6p3UC/V+G5sWITrVl6cXKUyJx2b2BdEpS5Yl8A8GBcGwGvziPDnKO
DuAhVk05tF94OZequ6I0R42OJeZRH8GZWG0fDjkgDl5rDpxs3icQcK8OLbxeGJ4y1ZTSsUIDL+OS
vTrgRbnj5SAGkqlRA73YOtnHD0a6Q/GIjUxmXUwRgX0IrmhbHkHBc/pIQfHZwhEDve6R+cNrXOUr
+pgd/litj0HcugteQuDXujOhDT11cDkk/4LQU1ytt8Nz46XyCLnJxHpw8mfHT1kuSbG3zV1MzdAr
8r+Q4uYfT50KsB/FK1VIZX7wnArcepz9Mypb+4HJSfMnNEFEzMXLfNml5I88G/ut9kB5X+lrmDoN
baMRzhk20T5tHcRLR8NuO3Ais4b3xm3Ee+2TnKSuUlaPWLHsk8gNt//y1SpoTZVXhqiKwaMLBZwl
XV0m1t+NENOcwe/1cOrdu7oHOKV0CHJULuVq+m1SLTh0n5ORkNMo9WyMFtiBpPoGZYI4gd2hlD3L
7MPA0Fvu9GCTj5RDlotdQo7d/IJS/5+S+dUk1cycepOQ/hMl+I0nGdD5mfLMy6joSCJjMOQVNg+j
22Li4gqQYBFjhH1yMsOeKygs5z3vUv4wa0pjNZGsKhB72VLoqaIN7e7HhMUe0C4mfdgvixr42/As
3iOqi0c1oDms1hj9GZwDHEBkFRpxq+ZrYcsdWU8X2ELdKBR9tjAq3zX2j6wdvAxr+daB48dGQsRQ
4t8x8h65PCDDmTMeneCXT38B+Au16vE7my2QR4td5Gi+zKWRx3NabTbO0v5tUcmLbQc75he7n9bc
Mwtqyznw9z7QnoU7Tc66OuqIFJFGtmbnUQ3I3yYp4YhuzE+0PruwSjFjlBw2eCYyASOA6RJRVK99
mqvah3hHtw2qjuB3w37PfZzS7lA1l+xKHL/bhnd75qv2oUyJY2EFDIknoNvZsRpw0WVa8Ql2+Deq
9FBF0iG+3ISSMKm3ZRmMtjjJ3lP69wQdmqQbjs2KdnPDr/ZYyqokBo5tMv2sk1J3mmPZ63hexcIL
Zts6qRQ4uaOA2C2bEypmt3yZWhhSFXInwt/KBK2tQ5iv2F2GEZd9YxXdns71gXxS0PX+zKrHFdne
48VcaikYsiZnnDC7zjkcDu5SddfVrcr6j4UJWma4AXnkP50ZIDueDfT32H6gzEFltQF0IwS/lNgq
HHPhHDBFwgJAkiXqQaMvEJPtCwFIiL1Ioe1Ht0mIsHvimrZ4koSr8PjBbdpe/HkoZlZnjbJ1c99I
IknGwAbQ8imyxh8dOcpZQtc6CcfEXkj7qyezbqJ5wVE1cuMoJmEcRvbIxQ9gxX0WUqAgXSLynIUE
ftph5YZj994dRFENHjZsH5Jz41d2w+YyHN/Ygf+H5Ln6KQYTyguDqq4EjhZUF/lc1Z0v+hvt5UKL
r7ICtNMeRO8YK/o7rf3v19OyHVX6jJTN5fw0Eg16P5tuaLZEXGBuNiQGi4+0bH8ek9W7l39nAw1T
JMXVHV7azYfQ5+Mem9lC8mBJGLWcd8X64qLJ+NJtVJcX8R+RtBVmXsFz0nMHIk0S3B0nQBK/dADh
J83jD1vMxw1b37MvGfJxFloDuA/5dQvn6/bdixvrh1QWtDfJm/eFz1axJhCifFqqr9JLME/DuQGv
Dde9IazerzVEdPjSrgkCp8od6FBCZswhavKAKJb1wmVNv4hsvVR1htD7XihqYxuDdHjU/Skre91Q
uU2oOB45NGUPLKlU/ZqNK9Ehz9bALwvlBgSJMGcT4j6yy/iZWlIBwBnPMfObC0r8QCV3N3T+rgZk
naV09EUFdS1hSNoj9+tJUWUXFm5Feoz8+7FzflWCecKUwX3T6z2e1kPLy8ZWqh5unkZW+6vpT0mU
32YITMHtoSpG2MW4BhNXW+21yC7P9k0Qwxm6tPcbkc6s/e4WpirH43zusJaGyoIKYc8SdQacNU+N
7wrieeYwau305xII/U81UrHjaI3o4trTXdAFXiPGUJsxkyN2UoNHGiOHcaVVVExzDR7atEdXKfT0
3LC4fxKgn6+BOYyIc244KFYHm2nQc763aaGbZo3U1tZ02AvmjrcqELDx5+/iSQVx1ZdkNiCvfPIi
Dy6a+Lm+COB3MlV5CQTaWlR/f2KEHXkjr82JGT8dANkCsfnTW3++pDXko5EffLlYr+h85I+ELi+B
46G/CMDuTwj1UTEqgO0NF0oOaWmmRCeaF1bsz32duVNtkQVzl21UKBRQAyTZucNLg75jgD1rvl7m
ncFF49qQTC9+PU6vcCGsiq5JVAimmsW1TxaAYqHjpV4hL7hVasKOmrMnPE6mNKjHFrQnRe/K4ZzB
zajDDkl8Vu5mGulu2po+fyAHGbyquk2UNzTUug+T9XuqGcZ7k2o91KYqQX+G9YWT1Ys8tenVh7Pf
msKgjt720zASMdRrmfc91o8kW7KSrFkIuxMG5nBheG8KGWhYhoQVmzMaSRl4OqIgrRBui9HtLk8R
cTqWa5ZB1OUxoQOpprwwEIrLrA6ElZQtgVMFwp3Aze+F5pHI1e7tztFx5KbA+CRh+5SXVkH8hIAA
Ciyrnx9oihKEermMqc3yf8kML2yADWkfSIMJBXaLgCcnSrmi2NtcqsnxVFllo4An1j53N3EJ0HDE
B2LFV39dq5sKPlPtPEQMMSikVqjbPHLRodxO1yHhdwNqfZ+stCYHYdTT2ZXWwff+P04NqKZhBAaj
BthBlV07tCmHLRVtDDOJhYH3JzP8M6npysuMLnPAu5T9VRmxYd1/vR3JLhpXwieX7z664XfKgPOp
k82dhQYhQa15OBHPFpUmNd6uZaLOzUvdiBAtmjoYuFmzruvMJja2ZT6KVHFSywSYpiOYekFvbzqq
vjAZars/Zo9H5O8n4dIUdDeD57gRZkzFgyVGbARXOJj84uJOL1mfZFZ2fnjWRAn9+1n48rTv+hYQ
PnNiMKO6VfxjmtT/WwEhDM/VoLAY1f09XF0TEXtG31i69drPYco1hYhHf389p+T9e3PABXf6C0Ri
+LHhz67TFaE6Ed30Jg6+ygWiQOCBqEmIJ5vlH+Pg/BVug/L4WbkhiGvECHVu483+Oph+b2o/RqmT
tlBV9r/9lrAoPv/FEOX94pcYMleSWlVsTczSjskkB2GWhGbAjTJvJXedOczI38YF04PfvxxsEh0G
0/oikPVIRV4AVddC3Vdc2uOwpHRi6EwBw2ai45hvLdCGe/PNTumXqGghtc+Mc3jokIapLBO3xWRL
d6UVSkHeo+eXhD3rkWJ1KN8CISvjKQLHG3Gk3ZQN6cq5DIz7tbvrzJPGCETv9g+/qgCZDLz+v3bZ
JwYnsXIDIC8KCqd0oEj+T52WohppcWTJnNgJ/L/fACeT/sv5hHoF6TC6XrwKa7n3ex7crrKbfb25
nXZhFViOZTX8OsW4M7nlUUOlUGbS4z72JvWUuu9qVX43ych7BmbTYo+AtKQg+U8OTjBo3CmlD7/o
0XWyzbkzcvIT6W0hB87qIbM0HFe0w3UHGJ2TWhO5tUGaNo9l/pCAcTbhTT7NQCvEHFuyMpgg4KcO
Fl8XvceRMehG1+kiuwRnSDuWcfinVWDH3TvHwnKY94zw9uUoH/AtDFS1GEkJBAx3GTboTKNqyohb
dSnzSJ1nY9VA4K2SddswHfwHFtijuGcv+0tPZWWYUXHxEmbuWEgUadqRUzToYjqO1IEtecsDQiik
HqBDAhyI+tElKnr0UKtQCbMp3aWhelviKbu8/9hJW21hPrxVGFrY3YW1kRpazuvPko272y8KU2tV
lGueRwnC8zY3RQioRIXGHkW2JH4/4+qKn5aaxbzN0SDXERq1zxJsozaYDgEJyyv0/vjY33xBOnLC
pxOM4rPpMiv+iXR8xUjmOSO297kb7rIDv2wj1DMQ34qgHtmPyKeOQPr8tC+z82wmYOnUAAnqpASV
fkJsWG2F8wfHJQMWUs3dRAedy9fI2RNz+Ew+4FL81UYv1+bleJ0Bwkj9MKPAbqnoJCRN0dm5VuCG
Vxncm0ynPVloonKT5ZQl96RD5V2KbB9GEQc99jgPY5hxMTA5hj1NkWwPmw2ZLntYw0fO9nIbfuJb
ve/OLvzF8w4yhPoxtlFP0BDc+/4rweNAmE5SV0n+y9v15LsvWjUVQO4CQoBSM8sYSXRTszpn+JZL
Xe5yI/5S97mghmMPJaF1mFbAoUeCO70vwMV1nLYpf0CKu7BWM2DG5WVULmdP6f6lQVH5mtGf1mWU
zbqsN1b0AcF0P+yf6tf+tfQLUJjzVPAP3tvTH/kmMYBjZdPI/VdTgecKHSXEUjQpEa8BD35W38O9
f7v5vAs/Os27OLvTBolra9rko65ExNX4p7O0IIcdXdBKehDH0xyi2t37AosbBLBmhF/nm2qShAv7
qGBmvb6F0lzhgMKIVFxYpi9UeO0OLUOaZh4mreIMtOq6tSo2hARIrZk0fl/024Vtp8aicRyyejY/
ixP9F22Q1d2b5r9dpGZd4y8x9956H50sPP9/+/48a54/lrD+zTmV3Ji5jXM7HhjQoCF2hAsJfOX+
cYg39Qahwdq59EPrTSrEl7YjiIA+8QDn8u7DKg3L5wXtic6NfkxKxcVY9xX56AS1R3GYFdsRn8dI
qJjLyNylgyZ0LetHDy4PKhGMDIo1axPv8xES9tyGlSEW1AOnEhFhXADvayX4BYXG1a7nJVb0brUZ
20Upk5wxmWyI0b/Sxy5Na3dWQs7+4hZNQ+KkuBbvo58qKDugar1yj1+SvVSqvD6ZJ4UlMsoxQm5d
/WczThX6QB78/dD91KELEbxRR1GFcS7Bc+ywXbO3+o0buMLva6O0rrpCWi0JrN7qVmWrlfn4MoTp
NRRjIwlshcW0TxEj9dlBzBg33TKBjywpaw7JEvf2bPDUnOGMmJ+uySj+yIE4lapN+7LD5SALRRKK
GbU1EKjDpQIDo1uirN7BXf5R9wzzTk0ioQysbQZ6Z16zuLxo16oIn0i1GJrfCfyIZol4eBYExe/t
2r0K1LjThO/M/KDQ3sVS/KuP6d/L+C7g8hraI/81Hca0OWPztszrxGxX+XoVQYQRuxitAAbgM+WY
3Bk1NLF2V8WTggDBwXL+bdAyM6hBaZTh8Pe0I0VHTKEwC5RLvOFQ8PcvZvEPv2JHxc5r1CydwiPr
hEBueyYE6iD95js0ZrsTjHhxa2Q4Bpw/+2sDoJfADrBvvQqdwYZSuW/iYATCNc6otrwYVL9q/zvw
HzKJax+ZKzB3P/W7zF0SCodfgtUKDM+VWryf2KWpRGNehEuKgxaxHEEmLvuOdDzB+9fX9xKEWSgM
OnxRzl8sbrLbWR0g3bWVsykx4/03QHhhj9sy0iRja7UoEP7/dl7TS8Sbteph+OMUOM3mPNeGDrbW
+CsR7pC88VJIzEySf2+zrHXBoelscHMtJ4hFJxlq67/g+xK3tEqgi2tXHA+kfqrimO7NIL1Sf3no
BtrfdLT7pvrtWnQ1VGghlcsXcERaqbvFKgFw/RPVAqwVUpn4b8H8i/uBo1uT+UCsiv8csyPTx/Xm
K2Z/6EePal+pTA0y0rFrY6TrIgC7SwwZRuU7PhQzM/ATV4l9/XE2hvkrg8ls1/tAuy/s42VpO0RY
f8cvXfnGrcjg7+nMU6hdVL1YZV1/j9heZfR4qSZID7ZRx5PDvw8dxHFDaKOHuI/mj/k0ieUr3dJy
bFPdvsvc8Gbzb0NZCvJbPwmr+tUnWYg6H7yswtbCsuSgA8caaBaJjnbWVRC4QOhBjuELG7UNb/MT
noQdNeg0wmBp6mR3aFYHqJZtdaPLRhfgh/uyChCeP4qP/auUq+pn2djjHdZWDf1MtOOz++GBaRIC
oio3+AVcHlKmlG5LWBTyG+ipxo4ouatyyDzgT77yyn8tyn7sMpsOvh368ROmoULVXotrU6NO0mH7
Tc1SVw0Zd+EvrnHWH5AmRrSP7aQxab4HPqLJOXHmXFY6S/86NJT9pvymAw8jlYMAt2wXs49e2FiP
ZrqjodUlcAKVpdAZNHI6JtMC/BpdVbWLuccpirzHVhOh/RF5O06a9UH8q4czjVHd+UNfrud8fhAG
Ucc+3JFcEbt8v7s0CEK0okLB5OVK9TnmLB4eNXdxLZ7Cxn+r4kNnHPi7Gje0lbR9YDyepqPmXCoN
2RuI3DT4bmCFrYX/3KDGoedDMgw0zKIfVQL78uR1qYwVSbxX5pfvVZMzIXJZhvJaMSCwVCGX3iKg
xxMDkPHs5W12vWsM7eskD68ItnnV/NVtX/kAJfydCOJGga7WLDmEu1Qrdegl3dSnOnkJ5m8rnBxz
msv4Xr8Z/LpLgjGEDpxp1B4FcHrB5iFvOMjaVCDVVxKoBO1ivDR7f9o6Ea2vcdslGZxWGlaOg+lW
ZCbZ7EB5SsWzdgh/cmO2Wc8ZFVB05jZFBV8yHfKMV9Z7m9EON/Dp+6V04w+ExOr3+7mzqjP71by2
oqyrrR3KjDIKdEIeGM5UOHMn14lzmAE54Mq41dQ/KBkuG+3dy5vowuYGgCxs6r+zQMgQ/OgkCgv/
z63JxyLyeTV+KFODfsdGWZl6MSkRSsnR3Ch1++WV5PYCivl7jT5Z84M9fy6wBmEc7RJVqWb4pbhd
H6QgTX/9rSZ/2G9I25mrrCzeXGMzWFG2RuFQ2OmafztbsRo9IZ0YyW5KNhrICrdtT0Q6UkVQHJ1V
mpeTkBlKY+y1DVNdy7w6DiK00A3qBQUQeCyc1KzJ2Kk7PC1j/9UXKUlcZv1ImXP1/rzHCYydjJr8
r5U28vhHFYNt6crfb6kGYloXR/s/GAEyQd1vNIsqN9OgUNLoM3av6eyt0dvMaaJ85qEB8InXNB26
KpStOesHbB+spRIrmectnqvoe9VhFpWrTH6yxNOz8oUhsvm2b3GW9ydHBwsY0Ia0MjUlSmAEqZIC
hwnf2Us3OkUnERPDuupf272ZpmkTMWg7Y1sCYYdoKV1flf0cxSfamQMhZQsjvXzcGOhZ/FuBURsw
Fd3vJqi+DEH2zp8HP6tY5L7de4S5dmU0wxJOwZvQ1qaMqMnRUVa7Nqw1yLuNJ2SRA4JM8wE3u761
fmU43w8E1NrhFZyIcwg2cAuIYMT9t03QBt3pgGbdgODK2q6RRhVywWEkFACYTVuNzUOYKtKZdBA6
pvHeQoBTUI0I/chAl/9NuxsWdV4PmbS9keo4QDFfHYhQDjsj4a/dU6QDIperqYgUmfeIY5UQLTbS
zXbbUQ2B3H7BeuAOY3wyArLtGLjm70Kddv0ELfFTjv0RpaPqYMDDu8XEAcFAG36ZI+AE5IEEnyOI
EVppDsNcddUtgF3NseVg7SRhtTGt2PJxt4xUII6xugkIuQ+YmxUBgwD2QtUdWwm5B81lGIyJ5Lhd
Xq4e7Ndc0CTXfLkKoQTEV0L1sbtoER8EiF2QY/eWC+RqiUG3AaHvPigwryEbrs6uQ1goqNzGT2P1
BrSrM56VWUYg2MfBwXe1TGVC+hv6llREXsMOeqr00m8FW4JOGaUJg4SCgaZFWBrVh00ON215IuUy
fxVHOzSOoUEeosgbDZpkRi2KefFGTEYoPb8WbIB5kakpo0M3/VCsF0g1r7oO6NG9V5Zum3lnU9sQ
08q3v1+ZjSZO3Dj8owRj+EdoRNyLhlu/wJNFD7QhaRGKMKExqPI6+ohycr566GUVRU9tiotpJL3I
XzZskgcv59oH1+M9JIar2RPjLrGNhbkCPKB3595EGQS6LUhr0Zwh/IL5QR2qfgn2ex49Ha9xGFI2
LzKZiomHxvYveekRPCEaX8LWbN6eRpsGkZTB2PytVI2TJlsz/gwBwyprwkNj9MDo9s0kgGXxSk5w
DbudnUOdr8UNN2ww3ZLSpnqjvYO2uJAaCvFgTPWiLwddZ3KVXSBqj4vnb0NkAzVsy8m0ZAGBYMin
+npcXAIJ65vHAWdQT62o+ZXFvP4UQ6SDHfhe2hgDvqDSgrykiE/EzimVSE/QAINiq7E55JzogRLo
6Zshtyitj4Iw7DDVbSi5C1+AK6uRg8pE35gaEsIQ2K47k4D3LOjhPh9l0dVAkZqxRr0uRJngui/K
DOPbExf7UiLByIakKxNM8xzQK/LeF8l6puh6+xPqqMTatQPh5pS55cI+/r1sn8Ml4frI5Fg1ic7S
MixmJAVImVDneHAjYJ9oc6tvXGrdUKEWbgCsBepahjSkomNu5AWTdfXDR2PSonFGvtskeXIrTm+W
q19duqBpCRKaVXH7FAfSeUbEoybkgFqCrABtfT5bCZhIzUHxeYT3SAMYn6V3jdPhJ+zws5TucDLN
Emi1Z1InsQdiAOazHURUlhzoIe7kXqGemsfSFJSgsf26p0wudf+82Fcdy+VYSao17TmwsShvpuaK
2POLRKwLkb0DIP4h04e+DzLUWRGzU/UZ3LIOlaNx8LRdVVb4CxnfZ7j3ifpo3OJw32UEArzYLRny
FYowhSgbrGV14MjR1C7sXvNMO/hWNg7tWJL1wzEs1a6wozi6WicrCAHjzKiYeDumeb32uuVxevPK
m3Rp3fGX6QH90IEDaWBTUrFVWDW3pjhVNGsP+4czUBEwbYo2XN7Ny8XnkP9Q5hOPttTxmRXt4/qO
KPx6LMKMrUf57E9qTHeCw/OeNnIAqenYqx5c7shLr2VHtz9JlZjMuRrQdNy9zlNtvz8nwyVQxSW4
21ziGtYgU7o1IgJuCrTMsbkqd7LOY6ti5BegoupmWXYoxQ9LMtPPTpECcnCElCEpXqTP5SLFN800
qSAY6/E9DAOC+9RblSt4F3oMVy3JiIqX2bh1rxJJ7gQBSl/STMsF/alpLmmDqSDGo+aoYJxjhyE5
b4+P43x5IabLOg+u+1trLgn9AofRjtMycKTQmBCnSSTWu3vfOVAw+LihNOMvwuXUUL0fX+ffl5A0
M0vNr3AF/iZ9fmte9W9NTcI7usFWg+UVUAbb4LoBd72M4AtwbjkxIYn8b+Eiyr7wFT78IkR34do/
Pb1Q+mqZOlvTZfcc/W66hP/NFH/tPnONiv1ua5YfuYDOV5SFLnFPD9qgu2UiXGPiRMlT/hLghhcy
ffkL9w5xmZpxOq8jIUaPmt7STFPGNn5vFF4lmrz9IzLjLpjhEhOTvYZJW0iXwUOxcmo1pJKoxtW5
uZSozgv45ySjBDzzB/lEIw6tLPWpqc5Xmb75utnnWd72hT8ZIb1JRX5K/KM2HlJo5FIJ+qhnWLa1
dOYqvWR0EYOByNBiSwAwfs+AsJ0zMWwmRHh+GX/jlhYQjKM7+JPtkVPijW+L0O1UwL5UxKcDtRF4
rFVY1jDhK6km9Xu6Am8Q07uGJ/+/EobC05Nqc6f7EJOJlwnAPmLKEMr8518iN5i00tO7JiOQpf1Z
hJKwhFGnEMzEjPjHxEYlTWT/JhhnEIyDkcBssK/DTNCsV6BIIivY4Gk1zJn82q7oFQdB9OZkzGlv
GvPDjyrEsxSd/zzTLZgsPCuSqY0cIarPO9fTw609uCrbbjrYCQd86yD4ACAf/rrsN8D9PRzitqmx
UU9s1yUVdc/dY4elDe1WY3u7cNZTwOlCYqhadlnVb5aALXm5EpeyiEFNBgDaG0Ya5/+OqWUioE2Z
mEpyuDp8xRFarPRweCt4RCiKIO9vRw+vmhmZrK8T1tVkKF967qG3izHL2LL3Cl39BuoYNXklT0jV
Ea/v6AbzU75BY3rrkXxcuw08jiceQ+HXzG6IAniy9lc1SsywdHh6S3myu1pzUDPtkr+UmDNSTrZr
VndboIx7CzkjOLe+1fK2cvneTJl6HcXhKPMsUrUIqnLkSM2ZtS4KI+FtzzB0FnF1M+PUQgkJi0FN
C5iRaba06z1BKTc2Q7oiP579I1ZVEbMECYvzQUklAfmEB2BCxK5DQC6Q0KSJOZCOHTI1kkmkKATh
l0B934w6oFtUVlRbiAtvOmnJLW/mp3Cw55Wr69aTDycSOUH9KtM/WQrce8wyD9euTxyg1YqMU82g
FaoCCclwUhSzSx5vKJpwxOjUCNjs7X6mVhxpjhcHuVh4MYMKCekcBIcIB825Et4ebk4GQQ7R3Bvw
7W6/JwTj5efg0MAwBegHLKr4L2vsPyJSNH9o9TKUoJbHeGJFzuuaniWX6CPIaFmjnPT3xA7UkASh
gcJLcburRYcJwidYftdcrXQGG1fsniusWMdQ+JQEKcV7UcczQ06+snnFGl1VZMlWxpDAc4EWdchk
cnTiNpbsFkGnxLT6GWEiXF27N18O3k46ima0QuvmYdMNOTxvShHc3dKs55KiysNhuHz2xF3uOUjM
NiiTTByLO1pKQx3IigDJpJwTpv2qTWHxYAf6+ipm4v8dPT8ssSZeSJmRbQ3OjVCRr1O/Q+pjkdUM
sMHZNxrMJEwf3tQDzuXsS9d+UACWAAq3K7795Inqz3GqFZ/PiyP8IMG8nk1HO5xBSJSqntlgPJRU
Z/SW3UzVnB6FJOHT6b9IK4KIpHVcSbna69qPxbijxSAqaXHvGN5BFy299K8z71gom2CdT330KkmW
fuJk8TAYTo+yPiIXlVrYtLHcCJGvlqc6Q99hCz5Iq0aECC+dgsbuXy1oEFNPI2D4S3aBCj7jW3zR
HguxqftS17tRtFZPTRjj0Wp0cOIYU7jXelQkPn7S4IdQ4OXwWS+deE4eKnXtfqwx/AthMtLmR83i
AY/2qKZC/+LQE86hiuwr31jX7JmYxDpgaBLM6X+y2uQEcv9cm4DoJQFnMkBt0PbjLujBrDL/8Eg5
+653zdn3vhSNe+y1hNejeJ/MAF4GQyiO0i4Mglg2N0k73qTf2S+BUeUsc647O6EooCdhFxXNkcnz
WCI5A1JVayZQFeEy5Tr6deeiHzwHFL9B1sgdP8PWhBYN0bkqkd55bCOrIQEOYoUEG4YyWUd+De6r
8pQ23gvcY1YKCeSSaCwwVfHS3/jXdqd3Hzhr6NaJ1u1D+ItF9X6OWfutv142sR5UXhAs0E+RN47T
0lJ8lAyOvRxvl8d+RikKJkhV+U9IfA5KosV3kn4IFDKtsXoCQlfFXkX6Yz/9Y7E1GjPXMdUmdmjU
Jt2gsGHvr3lL6UfFJ5EnmoC1fZUIYZ2qabhsip813YNV9oT8n+8yR5zDWinyKbz6t6gxoLGp2bsR
6Vzr2fLnCqaW7BBZGPPh8aV53P0fVOZegd8yAmGPjY4W9fj66SB85DmewoBBnXLWA5g4aUbFQg2l
jA93etjQnuY4KK7Askfa2I4hJ41YwRX7YF0SoUS6qNYjttV8fJUPkoHqsvDCStm1xZoIGETEXlb4
spW/KkSC4T+aSqdgQ6cXqw7yRmTPnhyxU5fH5njW5kP4zK9B/QUiTHxuwMu6P4qwS4jyWMAjlUaQ
MLgf75QXeCUX7OV1BEyNI7f/KAQaup8tnMH6va838u1ync3MNXBv5YZ6BgYVqg96SQNqpIy8wZua
4LsOjF/VIp5KYygVGKg8r8z+jJzplxzMUTxvxzzpnGSXf0J/qvsbk6E5orYE1QIJO7qtY6VsnLO4
HKVLallRfqpTlRC0wPH0UNGfE30AJDbGaOZWd9ponhdUMSfN2bCUPdFBme2a/N3++jaWRVPm7IB3
XsJgG+0t5QtXGTnQS18lHZo4nFLBDoskHIFD2oAQo0TNGO5/Fah6P7uQKbrc/AleHylUy67ijykg
urRhUwyZUMuYWzX2BSUOln6jBdMB5ezpPXZw5e8qDQ2k9SMEu4x4IpMMTesCaflSvxZyKVKkuvhT
YtkGEXnLO8NN4aZy/6ESqzZTGdcse/79nPXK6E4ISJCgntshB+2Ar5mvXwphw3p6sH1fb2J+ftWt
C/zBvbbyhUq4J0xDy2zKgjzHk0rgU3GutpQycXBXC8MRySXvrXHakME5/+G1K/xmJybHNjt7LwrF
KPU7/98rAbvGPge3QsxRFQhx/0t/9nZJk/gdL0utqYS6kRd7deFJ8RYYXlCUlEq3CVv3tZ66pn3y
jh83BiKx9LNOyeT6rveftm2B0zIsMSrF+WK+Gwc7w9BcU3zCVrBNAdmBXYq3z4WcDl6312bD4WqO
gTQprCJsBiMycyCHbe0IvuGLjlXYRDeRscedgKW1c4TedCJcQeCeuZNFiqT7afKhownCKNTQ8Jb0
efyQ9V41FssrvEQyybz/IJmL46jCrq/7Y3TmTEnGTj3TVbO13hSRcR3It7DKKRYccssejc4hmMFu
MRYg9A/vmDnONNPn9q/iH86/1C24D+UWnFcCbmsKZ83I0jLqyourAw4LmGoezyPSRs6ZGKiW+7FH
5AE+USEjDQyKNJcDXwfGaly7wWTBdGsnc4o5xlEjTkkO+X/MdCobdGStz98h3k4WBj6l0NYWrO1B
J1QkQq+aJLV2QSeASLavncyrsvoCtqQ1TgJIttKr0LihpXX/cZc5hHkrOalz30o85CajqDv0CLHG
EY90NefoO4LjKG+xnC/beAiX82Zp+NmaOu7h8JAwD+hsrXH42TGB4TiV9tXvnLe+HwXwzS1OuXLL
IZ3lUckCFKC3UbMGzeq4m2Y5AN8CBCuNzFHiCh7MyticMkqRWQxHeEqEDesxOpHztaXdFHDLBKYV
JPWmz9boS3YD5NRhFIXSqVV3ejhtWn2dR7H+7fk4N3WVHgutcH2YKPJ6I1Sv7oGWRv01seMLMIWv
JY4VS72X+fmllAplf9/5rEZlFRWdmVlJS0Yet/zjB5utHozCXUwyTBqxmg95Xv0TIE2+SGwLM58l
7IkUiGPePv3gN5LjTob8GupQurePDqQS8Sob3zJuTaq4c1Y2iZvuh00VURMSsyLpKfL4e1NQeNSZ
wdzf7fpaHSRBw7cWVuKKPqsUt3pmH9Xb/BQoEanohx0WbR5W/3xxb94LizKp9ZT+lkq9lzDzhmp4
T4ltgOtXsTOjvzOHTMtLzB2ynaAVbwviP5FFFQueNHOlfUGwBIhcBRFbm/3UmPfqdva2l1fyqh2l
abCftkrbOOgebsDaK7F0e7R4nX6eT5XAxdeSJtChRiSrc9jq4FIwHt46MlWjokJBJ181pTS2Dt0q
25/u7M47qz4CgRy5TZiDmUTTQe2/4/7VyusKQpHLsACV7BCuMlCPZC8XQ+wgFntvCpFgsuk3q3tf
nw1+lydZ8IfJotEImxosHhpLxm2Y0kc4LjXxNyR8kORz1KZn6Vky+dOEn9f1pdkIbNHi+cEByGFK
ZHQ3C+s+bjdBeRGe+WRUsHhzoVoT20W/0pWs1cblC9ZNAsNhYufZOQG8G3XRnEleMF03xdX9scaL
wkp9SGktRkAOGPffkGqQZxOn0QFQnPujLVHaoKbCuIdi1sXiGAtZfP+S0ms9lXkoRfRp3Hhbj5Sm
83O/i6blWcs2LCt0MDPaxiYFV7tPeUaCYFzlnjgI4TJ3T5jUwzSiX0Vy+paXTmOOyRf4454yyt+5
Y9UqbIQH1GCPpwl6Dma8IYLJ5DnDY5AHOHmL0BixNBHmJ2b5ECAeWVODc8RASh+mM/Pyb6jTtUx+
fRKcc8tKLhkiL+jDjNvNBfoPouE65dO8e/u5QC56o3Hjn2D1eXKVBi4FFiluDmB4H70LoJL0ZOn8
jryF5hC+BHzDOLRwVklLG5yDYtXWOG+532JNjx5MGWWEPJgDRNk87IKMv+MbKkne4AahBXH6JZd1
czDtV8pqz3JSRfeX6dnSc3Hfb+Kcr5RCyga8wd8VMmC+EFVje29QAz0BWxJfr4WyqrPfdVe0jQJU
ZW0/RuW0/g7HRX1T9TfY7sSDkNO2zLswSOj7qFohrwWTz8ZEVva++LSuCGgQbwCRBtccT8FcauVY
xURDogkKWrBbEbuwBuz7tmmCdRXvwejZ2rshiP0tSJr75jvU1ORD4srJJDOfu+CHWn3H8dHpHZly
xHyTFaAREqdXb3OLbB1X0QgSDsPC3AjshyX/0FpgRKxxjUS14JzbLQs1JIA7fH09quEcTpBVd5sx
2++sZ2z4wpUHzOXhjq9Kap2d33bo+11Nmp9OlFqsZ+gvxP7BEe33uYM/hgf3IYcjPgz74eD4jyxT
/OHwZrpSGBp1owRh24KgB1PUXVa4iwtGOyBTmesqJyMEYUuzDGo/zyzBPFBXgMzf64KbAYyNOR/6
PXoYQvkiQwUPKDSN8kpisDDJy9ZR/u0WTZvuoJz9vwe+gDJgJrlThtmDNmWjwJHZRxxXbqk3uZC9
WvxPmw5KFBQnPZi3zg4AgsaN2Mkp+VXH3ctAi+tVzqPMhL+YtbN5S72nsIwH+00kv3Ux/T/hjm78
qPabLXRucBuTjy4XtodAZEOSWqre3bC8s2kynP4JgJK09ABgKXhI1+MBocKUweE+ZP66lyGS34Yt
vxYvpRm1QvY78DFYqQE+jbmbAI+wLpdKWj+usdiXDeCy5yy/085mJGSsDAtqjbs0rs3Y6irR9N4q
BoEDm0kHyKcfWG6XXHwEhk1YesiUitM+F6yA3MjRYU4kKgJB9JMViMeCT23EobsEDKaZeXd4qKV2
S29FPsMq8mnWW+th/gQRNGw+hdYJcvE+r2JoI77axMOdy3M4R08X7UP3Rk5dbdDuML8/UBJgqm0U
mw2fAJjA9QcsmTp+YJNF4gJdSdcwXgCX/mpWpnFjPz/V9Q6qjgt9JNzYMgTHTce/iNJOWI2phEoe
wabaYVkT2kaiguNrjqdHyubJwyuk7F51yCmoMayzd+ssqHU4ifQTx5G4OWu3y4e8Pbiz8/SUR95h
LK9TetA4UQCnGspmbzNSq/pVzpHo9XHMzb5HhgvkeL6eyrFuteDYHa4m+ltuOBYbrzB1Y2dWkh0R
CFM+U4HqfzFYsqRe+AhIrJwsakI705X1T1XWg8F/glqC2SYcKAAq+JCOtGL/0XYbipSfs2KVqhnv
08uGMjZDLUORvFmPEOKf56CWP3qdCNe+hZxqhgVuoAE3WmkmApTad7bq5xyNfCpGSIF8AD1Ea2xA
MNQ/CUrM0c693Xjvw4fAXvTYIpTI3/GnmBgyFJ2emQnIOv9f5QsF6t15rJcYqjDHNAE3KQuiNEP6
NiyVz77SVP7dAoi1oUPvy+SKZxXNlJ5mMsa/NHTwSv8ZOWTRG6HqZbIcWm0ND3Zy7rbIRE/RVfHX
aAXR1P09lvlXiG+WeBDBkf+8zkGa90g8GFvYNHOCGStyIPrjuD8cVCxYaJU9Lufgmwl1kUZvqU5+
luOpdv4H+41Bp9s7Vovd1u+1Pf1l6oUG7efp9TLX+Tlr59FdDXz8d49xQxiRi4qSxkd0Lq7gBJ7N
KNijERkzWpdlk2FBeuzLikqL5hujVJpJWguhwrmJuag4QPSVu7guBIsq08bvFLq1w1dXjltTsl0L
nISsE7XRnMsdmshE+MOGS8yZCuhZE0e3Om4t4Ihgo2Z50O6xeo1J47YYhz6JLcC6gLZdNKHPnqwZ
pzu7Mb0cgpWWj0AfcN9PGL0ZH4xeMgCHRIssmw0yPdjZGP8LTyWDD/0mLRWkRFFfxW2QDscs4cCb
H0HhLQfml0+JnYN8pYEb4RaWM9GEKF+Qdp4lgIZnjiMIejuaQuwsIu40LmbHvDOnAHtM4/DonjRM
Uq96VWZtmLgCNMpU+xC0t5dAeG4Wz5tNe4I4cBGr5dF3np4hvStme/aDjiUutyBSzM/rckxTER+8
ok7WsslaaJZkKuLKRDPYBBtG5x6oVO01IUWLBcSj47cQBjVpwMfWMKDDbWTVC2pdXT5Uaaoqhmbt
MZ0N2wPJmw+QV9dQd2xh+J9ttEunk/sOrfmhA89frOxZFAv/H/+oaut/FI0yGpdEAPY8txGQMwnX
D+A39hTm0rJmepiYGI4qou54EHtPaXQknIvU3tRBdms3wsWEnxoM4WCt3lt1PMJzyCyTa6l3dWTe
s+tFJFZbEgGywRMwtCc4iYfRpdyOY42t08Xc9ABK55ngGFL95A7MXdVJikWs7PPWKm477Fsdk66L
a5SVEKo6yz1yAS4EpEybFA7JUlUpHtvLxcyLFKCUgtu13MDPyPYZIFT7VH5JE5EfCg6m9h58aCPw
nlRQuuOC7ghFLK3qudMKxowqRqDHBKFctzCGVKuXjns1Pb9fCH6q+MqverEwIQoLaHxas6Ww9dRv
W6QWumTun8SXBND0Xe/qbvARuvHa2rwILXwlUWX8TjxycDdd51qFasELtcXJyi+Nyhlyjt6TIoCi
Ac/nYzNFnc8lze0jJgXzDyn4XYN3qOfWV46SIYySbuwSmtTVKen4IUdIx6h6QsGZQ4gD0752kKW6
RY/D/nFqvlXMZaWbwVWeHDg1godoS1IJn7E4aQmAya2AapsXK88mWHq+CnIuAOywfb03BathNHAV
fyPlHjA2KUgnaufyY4MsAwfgiV4ZRd9Fh2rb8VTw3iwVGp8MPt+xwLMyEcvIWeShES/ADdbUkcvt
Syv1CADkoY2QK34EFlXTn3UV7kiE59RTQ/n5sixI/MCvRKZt5nkAKdBbbdhx4eATmfFv4FxNByDB
LQEUEChOhjKPUG0gIeE/bGBGhGOdQO/4KeCehKEFEN2h/B1fIiyukTQwZK8NaD9MDBvpb/vFDuWm
ILMrxgSDMdWaGnza79fU6Fw7qxVy+TjXuP+jVoUFvgZdvderfhMD+ELwttW3x/7N4wf8aTDz+blk
Da2XJiwEpajv95y0LQVh8hapGz6ET5S7V6GGMM/EWv+eK4aBWunZS9DOxwqvvYKPcMCDmkwuxWVz
HD1wb8mQxTf60iN27Uonm0QH+q8hSwhqCh/5Wdfai/BQv+r9kfMApukw12eSx0L0vTsZU8gnZeH5
EcZ+wAvuMascSfQsrlo65v1PeR3kEI6baIS97uvoAyNaqbTbh4srvTNxdVDau3QgL9yP2uAYphfQ
Py4yAgDpdNcdyvXRTH7wJCLtuKZsMiKj59R2fIOJzcLYnQdXJtBVgirLA4knvJBtvO/ycEC76+C8
11YYshZRgYRjh+DqffjJcgx8hveYZSytKEb9/Dg5J1uy62EFSLLTZI1NR2ZbAwrINPUZ5DltSZvm
poBo1MIKtyz4cNN9BR+vHPr72Ii1BKDTDeUjG0ZIqH1DCHaM9goqWmu0tBaS6kcbzynKMIum7pN4
2YarShNawH3gVQDcuGadyG7ClxN0YMUVKYKlEPo6VcOET4YKblzWfJHGF+g+ieu17ADmrvKYNNio
faxVCOa+Kps2qWuggy+h/5q3VchUqbELFNbrbtKLLcqBCgSd7NzkEHJJgUf8ZgEmWK2JczxkyswM
Fic/V9ORhoTuwDh9LO4SBpZX0dPF4mZwDqAFSwlj4381vORTimUjWA7JmGITKQJu8m1l9UytHXDw
zUGtFNvTojjECtzxcrkIAgV6qiwXojVSBUQvVV/Bnn7KZCpnwvNF4VtYEAvYsgrPCAOTHLkaUeQH
AiQn68PrSy2N7CshM8rzxAg/kNF+yRWt7mqo4qvGEz+PpqUbyeHLtJDLY/ala4NNi3CIi5/+dc4Y
YJxflitNCo+S7ugQmwCZW4XX0WrlejTLp/n68lihEtW3DHTLNGVqACoMMVzNs70iJgtN5o6A5RI3
/8Nna5V1KTOCntky1/6Lm5TDfwOjx3Mphnk/qjR2QedS1CqGC0o+NL7T1TCUxrCrdEucCCcjQuWF
HRVqbRe2BLI5VHGdHDcJY2OAtqLprqgXsinwDS38pUEEPnxL9txXWaCfiVUXuTEae7lJTiTA8f7y
pUMFWzNylpJKb9XifYCn8qOdv3khhYBeJP0O0caJRXH4ygrjrTvD4uMHXNPyjScge6qblXHU6LtP
rCRfU5AL+6mCfWLzL6ZUNDf79luKmGRMCdn5Y06KJTTpnCbBfJ/DP8Y8Z6F5bBrzdcmeq7Cp55DP
erEuvYbVSJIYsWrOe4D7YFkqBYEu5P6nuH2/XHYejiMSLWaU1++WNC+DWBYxfXJpVzQpj2jOAfaF
tL84JHEIm0u71Dk/OQscuSq6tOwZljR9PkRCcfdSUTvvMmvFNMaMuxFBjbuA0fV9JXRiAN5qI4+p
m8Q474BBWZsJto8Jj+lCaiR1vB1356oNV9zU9wvx43WtY3i81VUUZZDU36uFxS9cZu287vfkWXKp
xdaILIRhrSbso2Qnsij8QD7TTyQEhCOnkO+UPlD2DIYNssQowiKjGtQmK/u2mcBFTF5xe4TIzGmu
O/fZXN9HqV8+rMVf54CllJSNiXKIk+wvar3t0W/s+Ef1McDsHG4/hPJ9GH1EumWVL4vr3/0/deRs
AJH3sv3PhzYYN4MDMWhhofzyMOdEm+4PGVDJlpCEQKnJup6i+iM7i3cFXJFxzxFqJ7RaU9357zEi
eaD0ris50nRvg/1BrG1ENouym0lOAAqBQvn6SH+RrWhZBrPS20hyYMx4ZcM7wRsQPcjO85g6YX1s
B1ZdmEBXRqilZjLmOPEDi3tiL+gi9hrFD3YSGDpLj6oUOT9dC1xIybAtfio7btCVgIYe+DxAjlrj
8NNn7Rls/hs58WvBm2VaYWbfptECM6tlms5mPeCMX2rpOvoNIQlk5RDV/73AHkKNDnzHEaGz9UfZ
QAZJhbpdqx359xupHrRbonTt8FUDOYAFxSpxzDbMi3r1zKycLqvx45PeQ/BPIGH+ZoPn7m+nnC0p
4nSw0ZA4sd6UflDtTxkW2hrkGZNe3o9EaV4HB0dyUdeqw7+ZhILjB7rKMqtkPXmO2/zMA+4qNI6f
GKLzUT0WVyoWqdB00GF+2nmOIu5XoMU2fqqTbmtfbrl9MOCUZivMbihx/iZKkoj2fZYQCY5ZUQVk
5/3aS7MZoPONcrZCBXYv6K852GQQugbU210hjujFiWX70J8NT8a/aRJwseoeLp6tHxPpOausEof3
ozdtK8P6DTjLl+F7bdMQlFqQywQgSwxUYTS+YYV0WjdGsPg462T6FpFK3V3vuKU8sO0er5FHJ28j
yOXfpNaviqYiOBT3mLqoHTIjUUwuXOCLisLuUjfXH7OT95p1vIh2FRktCZ9QdLyJRBD/nogQdOiL
CWyEXbx2sahd0HTA2exDmefmoy2Ial/SOwjmIvnIlqEYxcqU8pizfmbZsuMjYe3SD6gGM7Vfx+EL
ulFRX47FiH2sFoChGQP+euCO+TL8CgZOJBPejd+B7ehYcnGak8ry5FwpSJZ2BhyMZPz9KppELFpL
w4FQR3c1JknIzi2NMCO/X3Y3JFg6bMiu5p+jlp3CibDuUp6QXOcChzFuE8/kUHbjEyQ/bwKxgLUT
q37AGwdaFkdpfK8Vj74LBICV89cliPBs1OYeUT68YxbktQ6uYYtTnKMKn21lSpPHC5AMdRUh61Dz
KXTT6x2yssLdLnzaH+qgwHOV+jCr/Z/cjqMqTXLHinDxIet7jTGP1s79vZKZnM9jTw3QZqQZm2pj
1zQ9+FY8Lp+ZiG66VH7biIJaydkb9+ZHHRu3Ot6xX42JTS4QORxcK3ckwzVUV0ekliwMV9AoOeV/
wkDj5D/lulQSXhqs1iTCKnJZBKxlvAycysO5hiuOMO3O9a/0iyrWGrVAoQnM3rp3i3fJnvJkuemE
j/E6C1TnrEPvCJ9oE14zoLX74zLbFnYmMBTLEcAKaU6YdHQpaXX9c2AQZVQ6Jvs5Xfys+pUhGh73
JXg6hsqS1guhZjCLacvH0h1DK6b/J+QjhJVzGngLv+9ecPJrU1LUC8bynZ2I2MMi1JHDvbehBtB+
oACk0q6jSh3VhZGwtdm59ARLDqG6mSFPixmpBJ5aQczpRDuQKkVHviuyx2M3AGybeH4/aq8j+ywg
qijG1ujsJW47kmDuTSAG31YpNTZyRzEDbzyTsH5BtQDEEbrKwEPQmDAhkldgPtg74uQKcO2uaiUK
LjDuqT5Lr+3R10rorypRkOYYoyTlZbDKAq2XHBeAaijevUPz9SXyz9WIB5V4ZjntylQleaCWgjWN
Re97xfz+6/4Z6wGV1MUd6kjEvo/iuoo4sQAicwA57CINcFkQ2ShDdyjOU1uWNFzItnaR5R6R4Sr6
jbFTu5SxIJa4J3XAWzKJQDHrA4OThM647TKr12JSEcrbAOhCyLKCiuLZKQUW0CPy9QrTQgK+L9Yk
gCJ5Os2Wg6RA7p0hpgL+Sw3ZTIqMW4L2f3bhdq/vSjjzrDVBrTZlfeXyf/9ExDNdg6GgCGrvtuJq
FJc8nEN10Ez65tg8InVEIU9Ww3p+uYhLGJyWS70lg6o78t31MMXhHdxpgVXBetfNBkSq9Ee+Qw9/
1I3zWyFD2b03Yf3rtfaO6wOBiQMtMjuLHMJ9tpURmnm9F/k33x1WT2b87zHAk+c6UiYiP2t0ot1m
qKMwfSvCtJhxBeRsQQtUH0MNdCBZbuUgwf34NTaq17C4ZWLQRDVJFa3PTVbhoI8VnmQyg/N6WUID
+46BsOJDNFcm09I27EApbiSvPclgCBqab9QE8FS8KlHWRYgu90ZpZnOAkpAVIOJ554eLntMKHEZI
3qRpqeazobtM+fsCqvPNj3UnK12/ah9/RQL6dmmCzgtBS1BkCUZ0q7iKwa8rGgy3yc8ez2x3Mdmf
AczN90/vbz2IaD5uYPNvpnWVFYrP8HqoH507QdOv1bEc/YKZDJOH+7q4HvK3YA2Yrn83ydWiy78x
qWwJa8wHvcELw3Yc3o+BZip1CL6FA4wxXsJQICKcPX4Nfh8pDDk+K6Lu7v+DGsdZR06NuQunhaCC
GO6yfBWDFxiGHsK16KfK9dsaXYpLINYAjHZlHWP2jaHfbQDUypmGsRorK5hIP0xmx9j4LVMTojQR
mzL4Qt400ySzHvnxLl8k3G7Y97L8sMOF8adPEbG2OeL3KwNz0cHWKZcCPPgt4rUt0CHXgxEX6uRR
Q+q0h0BuNJT60h7Mi+djVIjdsgUuoLyLmeVu1Sp/frmXsPxeWVSYyL0kJgrzXtRmZe7gIBKz+aiH
Y8htUdeyuANqX7DmW7efTnwT61i/pqj54LbW84eeaGw1v/+mYBd615PkpKafKDEi4wDzFUuTpLpc
4JDZhnB/D78dXuwMsQyELvgyAq1iBwtyPbP8vzqLR2tYbdIk5QcwvIzZLGHtQETQtkM04k6KN3M8
JpgSt1dS6xlbL7kdAWR6Y3RCDbZoWvrcwGrTHqGMzZoWfe7GwaoLVB5MwnP/jGiBIq7dzhKfVCG4
X8ZnAerC4Rr5M3KswHG5qljLjaGHsSUMm62+ti7ulPd+OaV/nCdWxULVOU+YsJLzsQmedaHZnnO2
NwWaq+msuDRBZQEATMf5hNx87kY4OJHwbu2qWOvZR9jDfmum0YtuDMuSDIvVCKgGOnljzisophPV
ZAepXBLZg9uBj6MvC4WRZqoqBwGbq1WRaQJWflWFf/MCqP+qz3zr3rUrl4kAW7JMLa+LqvjjBFUZ
20AaYUdPKQ33kAC712nP/O0ayakc75PRtrQ4pXjgDaOby0NlBz/FHTw/r0kPk/MxOaw7NRXehw/6
0ozM9+2nqK0nXpwNzLT2EFpxUAu8CgTGouLSdaARti9y5Xukjd+7HeXxerHQYIoZxRQ8YCPgCJn8
SJkXGa3LoXhducCnOuw58kPdWK/FJHz+Si/a+FjrBIxjwayngm7ryJ+pgO5XnwIQJcStmsbo33td
3B5I/+dM//48hJS3HqYNsdo14Kd1aRptem1/zWiGdf2bRRQX2zLuKeg+p3KZ+eU6MQTsovufpf2r
+3+3iVuXD3FHSVMC1THh5FKSxjwOkKOaAN58yUMJTD86NIRXAq6ISwjXqld4OGji+YpcxjXgjte2
yqHE10h0aXyyFhUMeGwTDebZVo1BJXFNjmos0Puxx7KtxC2qdprMw92oGGfJXfWUjZYVT8jVIHTi
mlNLHoKzH3y6HMbG0Ld+6aGxmG3lqBreoZRe6soJA0142LED9o59Wm7bLJ8WmSbpQv7e4IIZNxFR
lQATdkf64UpIiJkkW1tdUamGjJe1dCI1CU5T8ScuVq+3bqcjIynJchZlPbBKE+Q2aqWN0VySRpmZ
0bfYR5lWH5oVQQZwFuPfpkJF6Vz8mKI7ZUITjd7h2YKOV0H568sFBOxV3yWoQCVo19kv95xqM2I3
FpwxVSUydhtZ8ME8Z8zBWKoM0QcuqsVc2tXGs5iA13550RBLew1xq+WF8YfMxy/LBgHCaO+fkwmQ
hCzbTlMBKN6PPpoOckE9Gq2IDmFtuCMP1RD0rJpIhnn87xRO9Forpx3yOOtmB44EoXKiocHvB2Y9
+FEjrIRotTByKCdS6j8e8AQJjKmfAoWE+X+tGBGzH7k7r98/9i/n56cXV+ZHdxwFw7omrjIwY9ni
c6IFVcCyUwWk00lCbrzq6znZ/cJaB97BD+uZpOrsraA5vb5dDaDbgHtggGeOmP7kdXZkExKjZPyn
0PtNrP7VjaUeIJl6MyV2E0Ely8i+/XHF+Boa0rAREGeTQ/GdG4hoqJSR6Vnmo6aYu6td0XUxRZ4a
r5KNNDE+S34Q0zfQ1wSFKJZsxLudyl5I2uTEb2N1UiJjAzTWjA2iysc8ClAMF86wMNx+6u74NEe6
QuMh56IG0H6TIiagvI556tNfIYCwoWth9EXUfy5x1HGgyEU8GupqrgyoGH0DFM8gl3XadLgkjfn2
Kj1/xx3G98iKzwfqvCug+HgnKT1EFRl43Ur1up6FV4Wcm9xdiebYuRvgDScTqxD55h5qrFrobdt/
cgc2RJ9UWSy8rsK5Lg7iTppsqa849scEyUY6GQmC6EHXtxmpyX9E4ZMjkBihRejXivUoAkFdwN89
ynBzAp8/L3wLUpx0Ia1E+RHKc9HLHt01OgRhk3DqeDPP2nTvzU/ggBnI2c1f9dfa8S9x8S9WnviJ
VKA04+THQcLTzgX7I3/4J/FZslYDQNjIfj2K/0OHxjbOLRgXN7qQC08jAqyktQRP08M0Go6u74kK
xgEu88AHDKT+yu1xC8wu2lSpMfmTRDI6zz1yKbxh48Sj+ZeWlmihYV23VO1mVD4xyH0iuK5yIcUr
fg2aDrj9e9YUkny9XHiSkrYLtqUhdJNEK74hgLdpAIDnXEnR6pVAg1nYOtQGuAY+F5nw0PtITJ/N
4zivWuyvCyZEAcj+F4PtFF323caLAGNLDjrvTktyiBvHPQlwI1FshO5UYsmogR1JT7vvKEfwOYQm
hcTZwqsDNW4s4G+OO0JfQu7xrTkm8c4O+4NMpuDaSFA5AjtM8/0QhdJ0l7p6vcWHfNpb18aHD1mi
sVQUpI9nxtO39A04yqikRyY0g8RnGYcRJ3pPEgBYYb4Ma6tzSt0jT3fhY+XW98T5kKGN2Vzbu2Xj
iypm/qA4n2LRNME64xYQP2aCmb9CDJFDpnk3SuVhVnfnZD0HlH7EsuNGelrOFr0RAPkLbwUnEXKn
7g9+znSW6vkv0zF5VdC5v3ZtvFwS51XwJGBbj2zSGMBm32RYry0VayAi7CammnJDbVVOPHNj9OVJ
0iZUUeg/BHt8n9f9XPTqUFP+2Dei8YgPfbccpTiXDEGY/I3be5gA9ByUKtWYhdpkrz8c7ujCB/Qd
92Vy6Ba1JNMSzWZTz3aV7n4x2skYOWuX/FnIoL0ZIDfApQRGvaE6Mo0wlOO5/k7VV3vYK2ybX5Hs
0YOX+/4C8OxYp1S6vHNLkxlnq7ceH4LePu1R2NWKchuIvyyM7vqS3hoBifsNEr4zbejeFxKf582l
pAWiYfZfj1JwMYLoICEUkI3+rmdLf9Vw2dItb/GD0sUzgkS2oFVwAxghyfFh9pbL3MFJaleO7THq
P51rX77O/3Jtxw8tNaz6hmLAQCmYRWqCYykn1V3mhOTbSA+OKjBoNa4HfoTKB/f2pA4jHzjEUp3l
ZCLo3XQmEjB/1L6BgLTIPTuJrPQqEfS0Sn+B3cuyMO8kqgfuSNy7tl5rSZji3OzJNhtR3W51xPei
HOBwdw9qGQW4uIULyfqMkpjxfhjlCwreYQxQydAqFn73W3kC9lXTQxSaE3bjPYVs2FxhnRrnSYOY
S+7WCcFXRu7E0EGn5G7wZ9cdt5L3dnapTckOvi0yyfPWL/yPwDQEqgIgOW+zPwdUFfDBGYkzRgTv
FpkEbyMuvF9g+Uo+jLufGNEYsnTJhBwO9incj/EX/VeQ27rIG2fpYhwpQByHLIZ114tf/iFsxSN2
FVn2oX99DVVNUa+ybv2UPQssqSO+bPKHhvRvIykuFJtaYns703thQlTHamYHqsxkDe8eOScA51vy
z6AaUFl099Ylu0Y63tdSRZktDV4wnU+MyZ/nHCqWpg3vF5aQXQdI3Y7qabebebBeUeCz/Pwq7TeV
mHYymEtUKVCVQYmDYuCQ3NHew7n1g+rdoUUmPbAdVOEOvLKjFtBlavVSgoE8Vr/3hcZcy4DYQknW
FNV10wr/w+pChv4LQwSTuXwP2f2nl2iaVXSUtIjwvEoz2vJugQxiRTRb2+l32BCcbCmNbqc4q7lK
E/3yFMyeBDlou5d0OZLEFuLfCu3KONwQsjaRtMDYKYI6o9I6/mjxwdoVV5P76N5n9dWtzdC/nzuv
3tsQ11eVNikFErsM7I5QEFCeUsHc/KrnE5iiAdVwB/3H6iafTA1+kpIY+nXVQekw6KNehi+fokuj
MDbbW5kZ4wKS7OKoDZqnoVS9fMOl32MfFgNjeBUu5yqNjUW/b9bKNZyf/Yeorx1GGiV0fWzP8Mjo
R7GHdHqjVm6fYU7cUxTtsAcoVzc4OX1dWUr3o3HaGING0+wIl9TvTEHS7W3MvnxZqB2r0jRCO9iu
ugN2ny6yHCFxNuLjgWeKOoStcBc/hPRArDmhfvZpJ3BH35JYxiQY/1M/eq8frPa4eK99qupMHa6O
vk/FvCxJsZohkvuWSmGESW3G4ZqQ4SVTRcwd535J7kupatODj+FuWm4cr++q7pvhtnEo9T/cjikW
N5/N5fXFejwwRfLDd1VfsuB4bthE+utqfiEm3qjs7wU4GZn+UqTGndniB1uiuPqlstCHWdafttDd
6Qn84wp5I0JUr3KfvgzCoAsyRKUFf2BAk+K7+d+DsdSoHi7Vmv/i2S86MpX3J7oPjXLKJIoaddW3
ZgJyify+CPiNT6GC3nPD28KCt7Bi8Eiflgt4ynei3wj41fa/2TBdRaS0trPyIFB9lDAYLvzvuy2a
BfEBRKHqN+AfzGuaK/gBUBuiT3wbmWIPNmykU2f1Lvmr0f5z+VmREuln0AyLcsrkc96mxwWkPW93
bsslriXfIzpNbAkPr+wYIyXJuxI+Yfbju6S+AhT+sRuAaAJgNWKrxucWYEmEjGwwU2af31LZIqP0
nSlDpZK3qiFR1p4GaB5GOg+srh9PlKAZRqbLnqCS9ETOA2jVORpSqBUQKKlBU+/gIgBEo7XT0RFY
W7zCFWh0f1TXGcRTuDPhsM6nF/YRxjuL3aaIAU9gIlRgmrkonDgREpYiHArehf/XqpCy4KsHQHb2
wdCqOuyJsFCS/zFrzM0bGuYY3yXdBv1FEclyRaotelMVyHYVR6iFLpQhK7dxvr2zmxCwYhTujbHV
Z7xB7Z3Nc5WsvQGLvoiDa2MLkKDmUnJ/hs3WU+gYMSeGuJkzv7yfYe3vKqM611rjW1entDJENt6g
64mrLP5zdQm0QsF02FRN2HgU8QZaZ+AJrPgQHhP9BAMpVtUvvMomiychHE9qxi92/qxHF+VbFu+L
MuigYlrQz17ptRZhVT8oGEeq4d/7jkR/uZz56DFdDwmclYvEe73skTY1FxspSLzcwOG7eeqnmtIu
/RGxJVG7kO+Fa0m8LQFw53+SxdAYVR8kF5fDNZBdXkQE+ZzjqhxDLi2kxBFkoC50wPWAsNNjBvi2
nG854IhG3WwsS2vPdw+qWB+06vE4X1c81cgK+GWYoJpHH2tNxjXAd3jyjkIDdubjXfSjyMWmxwG8
ukQs0YidONARhVwYjAepH74nJb3o5L0U2xIXRGlVu6vPQlDxphAGSUqzffk6YKzX7fjdM7LBi0Ux
NltPGhrTuH6q6AYxgBC0gcWaaiMWFEOjPzqnfnxBTYw5NIBKqzSM7U5vnPpczz/1Jg111uuPW/xn
55lNM913V79IVCsnJ2BofVsPArqircJR9XpJFEsvIx1IR74CEXHu2XDviOv9sYCpJEJyQKGw0/j5
FE1wL3y6MhKhyB61PTuYaAs9Rc4fRLedeE0sqQynjAWRh/mtciCZAbqUDRKA7qHf39UmziaLcizD
ytKlkt2Ta3Vmik/NCKaBFJQno/u2yqFuRLsZgYfXzMWlA/JDP75AxPZQzAbmo8Kc/CTIQ2Ho5bA4
rbmhp58Y7b79DKRElnlbUuSNODMsTCs5YghmuPpizOQpA96Vnyv4UZfLiexCirq6axiUzHdC0P5t
QiMJbDsgCDRGEc65DMvShjWCLH1gPFhmj9mEfoe9fZsdndWhVD2tjOFpVGeGD5HhZRFAif7BJ0ni
2fnYCinaPSLBOekfym7sqFzaa135gPdkCFgQ50EKyWRduPtk82EO21D7rybwtyjJIK0RSu9hPbqG
hoUgPdmMsCkG25dE+tRr4ETd8xfRvuK1lsqOZW9Y88RXMlo10tASyUl3+oOpCvCVJV0x78G8V0Xd
IFJFpEgpAHDY/DZBELvj5sLZ/AWg7ercMlYbIZ5OQHKYm/u8XmKBwoi6GnUZaF2QVO4ulPKQrrk5
HGJ7+b4TlVc7LwlQ7u8MYEAao+1YfxC3g0clCrhtt+U6q8kkeW/auEDs0SJ0o8yq1TKuJtDs4WOF
iDSPoaGZzyJIYq1AkAupDtcdIiXBfY84uQUTn1EOEswZJz064XV/2KdGGsWaRZj5YEWHlqGSRBxH
NDE6eo5bx3cyACPUDLYapt15bWpFjFjocNz73wmkH+Qp7RgPl9F5LKZQQjo9yBY770LLM9rrXRPU
XOYW7sytwcsvbTHNLcSOi2TFoLkpI24rHrkvJZ/jj5tgbQofu6vo2xIbvL7CoLsjedjGj/DurXlR
WbMR7GZ1GVOVijaBUNJEFdYMde5G7Q4gq05CN/as8A9ocuK68f15/unuvgpQc30rld5d8DYKtzqb
9fw35ht7A0vx08+23OXioSi4ihXG1slBce2tPZ6VW0pMs91uAryF/YJ96OAFlKX4r4Tnrsb9xBMg
D9BwgrhZGNtXfm1UcNeUdK8ZI8qFe1jxaezoylGF1gr4nPVfZz/E3Q/uJ6vTFBqgMRZdKF9Ay1gl
0JaS25hlov2ssUZz7QLvN3RnP5EiTxrXb9zn2CsvWabc0yI2kJomfIJ+DJoGo6MpFp91jXT5xA2/
v2Czp6KlmrHe1GsDEJsfLR6hPoCNScXR+2HJg164pqMnT+Bf8yXA2pFc7Sb+cZa0EL60X+HBnM1J
4+GUYBTFhSc5iPq390DG99SmEQp7xzqOw2sthV9oFiC9CYklh+L3+sMSHUXveOb8au65q9dzjisI
PluwcmbHMCrvLGije43kBCGgJLOCGqO79oZi1iw8vvBPwOxc4cz12cYIVhyDhaai0OYhqCv1HBoT
uueI4cfgpcA+8ucNits9qg1h5e/mkCbhgZY5Ni1YqQlW1+iYK41VDJzASz7qb2IDTVWIDoPKM78Q
tF/tDP3lULlAzGbHBheV76vJyI4+aktL/TBO4FZD2XoW4tr5noE70GTjnWX6OUo1nJQO24L6xL0h
ZDBzgbwiJjHV4Ctnt1tTynP90ytS7elaVpVdJPAj5zS7J225/A9VNUrkBpVTgGMlhM5rEh8PwKxW
gEJ8qxErYJ6UK89R6YKlbwERot8D9P2Woyw+FAvx1q1LETxK1rnbe6fGchLV4Efzv6sLm/OaQfA9
7Kx+yZeWDemj04pg0leuk8jd3FyN6TLLXnmxtQxKc0RruAE0AKlaYNvGz7aiVRdQxqjdMLyDBgxo
lTuzxsBloRaoX+pmhNey74nLMmEr8Gw0uT1PTb65GbmHszIeSliyAGs4DDQdpNDxT3C0yuaPtU/K
XT0zs8kZcpaTgJYwh5/sSUczWpdT3bOMMH8c8bP27iY9z0lLuF61pKCg+9LVxiB5m/nqP6DEVzcC
C2wuvyzYwttl8UvMvs/WiQqc8w9tPcwDmM4VyayXkyzjv9QUKdSEak2tpJ6TQ6MuE3Ml7E/xauFl
xUB1J0p16iTFk2SZR4E3iGY2z95CxA+y1p05EVenseCANC9wV8XYoWnWtKq0GMEni6pRQbvyFgJM
MXEbLrv2FOcIUz6Qp+YsBT2E+rFxQlEcGSp83x33r99N2mrecv/ltwW1tWCArZKH8wfHEvsnubnR
4UX3s5BO4t0nTW8M/JLMJX1n+qnM2H/7kqs5fNEwuneVDONI1LzpNUEoIYvrQ6k/BiIvJfrYrThM
/A1kw0hXqEUon8JFhqU4rNjR1TPuKyZ6btw069oc0HBhWWOhUXce/cUx9xjvWz+m7wi/f8LaRR3y
B6MZXh8Up81bsr0zWYbytetlOIhGtfVhnd20lw8urER/pOICcQQLDV5KmoNQrDOGmbaTfmAH0DUQ
W7BEtwrhjEQ09hXbQs6djMcRrA4GMK6NgNXCv4mD/HeKiTHQv7dDxoI1CcTobvOxFYjoIY/g/G5D
PPyuxLyqsBpNZjB7slGUZeXxtauFMJ7/WQgfyZ9F9NVP2izSstTQrufIj/eiPHi8RHAZVZI32Rd/
fHxjyCzdpJ+fKXszxFPAMclODXBSwRZO0Umi5ipSME1BjnvC4ZBNH9Vrn+uCi18ZiITMra9+2P8V
lY1oSGFaHj9WwwP7tMcYdlNf0vQYbsebWsdIXgj3Ypu+licZrik1wHziarHYvN12Jr09hvIjY5qF
EDxj/0N05mLS/k0LOJyhE88EHYodIdto7NLjDZ81wc6ipqqH9QfPq/5JzvUIbE3QtEbkiojEvx8J
E/4xU0gQ8I1fHkZJu89FLzky/9AvmJ3dl3A+mdTIn6WZUyP5XY6RuNPrzTrDRMBn4hmxG9FH5zYK
VNzetdA8RSp96C6Blpfy9wuUJzrr6ndWOHI+9R5yvQOnCHx37nqxvenXxLGtZIAUlgB304CqglQF
tRhRjDK9QQPFjAb3soc2NL/5tMqCWq34ne72Zvo1zklusgpa8ic5JVHwVWrWnEFh2jWgGUWCpm45
Om3uL8OI/2H98ruiKAoMAZwRfjN8Lzu0LCTKPMz0AK5H9MzvYjba37E+R6/jCkjka+2OTIFQKrl5
JuYPR02ilZV2U+Iiy3g8z+DVDBxT9CedllOoWi41q3SM/51u28rAzPeVBglKlUL43BDV9rb57Uyr
SOZcy5PEDc9xU4bqK9dBxh06mAwkx1VatCWQs5wyxnJNo1hJuNAEPTN2aNOM6G7h4wfo6BJtLkPX
qa7Z8vE3H9G2FCtbsDmgNvmzp47GLdw+e0vAo/fQsfKLTNLIJ/D91H8qwga20EzV4iBKOQVR2gh8
cN4vx4R8DuL2nL9v/OtWI+ZnGU51QQ5ZTbVhoxRxe7FOEooB8yvUm9+ELrQ7RczmjjBSbFG5oQAM
36okP9ViR5f/41HVSZMeFZM7ynHP8/ewIyR/tSuMFzdHf3ZImvYCdeVXbaKBbd+PmxqKlIXFm8ML
xkInH/TvqzOczT7i4ibqidRvPpOJR8KKYKLxY2YUFbkwRnoYdgv5IzQ8d0CnCOADMduJWsAjkWds
G5EGgG8ifQtXggxgr+kiV8bIAXyWTMvRue8pmwHaKva1utzM1q8aAL4/J8Di/GMoQiHGh1Q6PT3l
wih6aLQBl4/CkEfFDAQ+vo1EGnMCpBIvqRB0KSj33FDzNMkspgVUftVhgEgwpUH8zrIHwTRJSy89
9p2hUPm+Uc4xHi+3EeEpp70uF+WOcEkLrEixTWyaVu00eC1TRWCIvLdOnxLom0ni6XKhvGDPPYjM
XksFFTMcoD7d0sLR0d0C8zLIZTmkegVTted5vKI0GGq7OxoZO0GAObCkHIB7lMOev4qknuhg8kIN
pZBbrR/qUOYQTsnEMpt7Rn3F7ebQJ1xo5OIzHrsqbZ/ylowCUebjsylyzNLzfz1DBTlk3oRZvfSg
8X1VoiHanPeEA6mDKghO1C4RfkEBIJQ/6wjJDadtuNfWxpsdbRsQmL6w5lXsJFfk1bpCbHgSyi8j
bgRdSyISdAPGti3pGV8ZJx79pR3llRo8TZ+dJhrvqC1+erNQoM+TAGhUk7NpnQKfAVGg5MJcp3We
XjnJT6WhxEyNDMNx5h+46BjgCZsfhh8n6yCwCvXN3ZTmVFK0GOhpeU3uKHcPA8JTowIbT1RwGqED
opwwhZUYvtyJXguZj32eRvmn+fr9kptr/dWB7Dcow9v6Ei9vP97bNZr17V9x+L/hWo3eGXYCZLOz
Jq5C//1hsE+fWpX+2Wu07rVbmnsILXR6JBH1uVff6HyxaU/dd+xy6pg1ECfFwhVWf7RcEnkbm9rd
ViDr7125V279dMUP0BLvHSvPzSGSjhNhhppyvz1OpQiCEz7MB+pvStq1H6nN8lTLxjYFxWUC2VHw
4DdayQRni9o8dK9NXzO5yo1NgXpP4D0ppJPWPx2C9MgBLIz5H9sOiLr3oiphnvfQWnd/rs69TUTq
3vl0lmunRWxR9ejyd2mPA5Dxcv6uRTFPQZF7jJqK+W7+gEQInjWaj37xPXh20f8s4dNvg+KChvnX
q6SrOpuXJEaLlwRfdP91vxb+PG2I3KTTYJUnDkb8ceUeWUk14UUxtWZshAbNIXBtTsZvsWYEx3Hy
n8M8iHgUr0MXezpW+4YyKvTQdisr3i6+prsmCbfUNCnWFjMExP1Ji0flx9mhk63vbOpHIsmRtyAR
gE30QtGm6prUKg+wyAxfUHvTuY4EmHup2m8WlKaE1K0ZfjxejiL0kI5mdBChjIA4JmiZ339PJcTJ
WpoVMp2Vfniiv2eeReaEsH60VaP0kME74tj+PkpAbALHOuar1hDAI5CkSOVNv7GKy+I446pHwCuF
F2bRur8mEnv87MfwCyQ1dEx9N1kc1CVZ0jKXR94dJtvcoOQxGCkSyHFOxP/i+1jcWQK+/F6E3yGm
KoHEJ5ly63JN2uE6vG9372iTwsHnnlFqFucT67xkwYkt65DIlBW8C3zRUF8Jk7sj4AixVJgpN++K
Q71nD3dricTcwtNloSTvVn1Iny8WZk2k1bXWb75wRzOhQZPcpZtH5LYnahujyPYOOEmP5zARQgjD
m+e5tdrmUFYy07VwBu0xzSFCwktp/V237fPtsnIDXSRbpal0Woik6n2fye1opO3OiEJkfkmhiBfR
VFfk0I8Kq9ZMoEHpzSZTPPCsmvqMvvVFBzBdVzEJc3my0p8iIblIwxpl9ikaMZm5y3UNCcD5pHH6
ratWpnIculk8xplysjq6L9l7ei+l6lau9hpOnLMERktZkAXT1DlSWUGy+oGd9EQgVAGINCmPij5D
u4/maoRIQdh3M/hSW572Ah4B3/jVq+S8X2TaWscwYg5JGXpaAhgSvVZsAMuQb76d8spXcUeShBvR
o1jTNZgAFtdtjQ0opmmzPgwaZpAKmcv+mQ9QCVX2d41gPmfkKQGRJwUWXso/eY900ZlTEWy87Kl7
uD4IgowFspgHtdV3nGaM4Hu1vIeI5u2pqdnpqV8B6tpZ2Z80favQoHS0P5jfWt6Z0vKs5hWlHHwH
O5E3b5Y3nWZcSFzIqi+lLb45fYf5pHePjKi+M3RWQBqAUPsrV0ZQ0YTKi6Nd0V27F5bvuGzzNm6Y
VmjIMs+zvVO1By3eAfe1Jq9BW9EMTd6w3bhn54zH2eaUdBfsC2ORo+pO5pGQiDkQ18vvESocYkMq
dDM9R5BDEtQxNtoEfzLhDj59oGKegW5brfjdg8ID9M1FBMH11onBCv/QAvLNoomCouKMqyOexAaF
NrjKqu0zXDLhFCNFMwK+pQs9Lslq76WjIGGGV55lnKuj+bIBqoygcUL0ILyYu6opNR/rxnih7Odp
7rtCEMvZuX/RawSAUpyBW2hJ/tYZ16gj1TaRah0M8PrbtEFIYCI8vct2h4pDClhkg8EpQW6mArK5
PeupQmI71+gBKw8uW4iXO1aDkPgkHYKptp0m2vlzKqQpVwOm/P/UR53D6FmZ7g7f+XHKRzh8F5TU
ojAMXW6Qg4FN9Q4oe8nGzVjMUvwUufcI6wymMKYQ45lA8sQBxKM6ILPoBofoIbjehpPA7JZciCal
uBCcS8tcVLSB3mJwiIGg2iRe1IYq9/q5j3fTfMaK5gY//Ndpz3FlyHXnN58j+Mu8p4MtTyE93vVv
obzMl/aQlB5pj3NESU20nfImQTo5I/wxMAGidrL0eWkorUhea0kq7As6BFJyUe9da7Cr1ij/FyCt
wR5VdYOkAtOCMcGKEELHH5v/IP7OqT4v6KPWTQu2yJCxbZLBwRIolkMazY/3JkINSSLEcL0o9CDS
gXofStAttoHzbFvH6VZMxT9IPVe964oi07z7+zZg+IbULQvAfdrxSZWPGzdTLa6PWl4Llw9A8F3m
Fsi1t55fD72v8teEll7VJLL5LgpUc3OZ6dc5xGsXJXnUboLxkJ7YGOXeMvUTqlzSr+D38ApN555d
ajOtncDhVCYDuahwRdF4jir4NkoV2Ozhcibnaz+ufFFUZx3pMY+09V0qGoSp3iPGRjv/1eEhlWtk
jsC3MiU2dWqUnGUnj4/n8qV6ygsIhdZo7qQHPUatNgTQWZsqqZwH0Fj3wOAihStRDzlS4rmYPO1o
S9drwnYUrotNzJEULBOqAABMZ+8XCoZ3fgXj5zKiNiczMbU9qh28W3GhgQvCJlRpeqK14Ure3VYk
SmEEfSn/wDFAvydq4QwXJpvnU+CjwK0p4ptr51nep8oNwkYLbTGZJlIjEVLzo//9iLEVsYTmEAS2
OULst7HoHUAMs6MSzKWPF2iJCAlY3gVXUNkUfRki4o1fyD+1ZMWVTJdMmuhdH+rAxjLGi9BrXbes
CcBfqY4a7VO9oebsNMBMxkJj626tGsyc0ktRu1nyX1zgQiuYmFa1KbLLqiC5QClHudLxiOa/oE+U
/nlmuDsC8k1HPznVpeJ0TCjFF9JgzFVl4d9fhCPk6ZOFqLFSKHaFUkMkHEmtnYRYmEthpWocyqKe
D8CZvej6Zz8xyrNnAibjA0w9IP3ry195t66mbBnG6WLvQzAZrWtSLX1xYzHif500H1B1EJyaVbEf
BfCbsRxWREAiwH0h7NB1soOA/VNXnTyHAqR4+KzrB4JSVttEALmk9uwdoFW9YwqEO4XueXp0OkFO
dwUu/8dV7e6VKJGYw+JwM4ynvSn0UPwxUFQw35VYDIbyi68jU6pIwRcSEGOcxuB2z+Ytdfn8FoIu
eq1Nkzk/hTsMTchu4Fu4C5FV470/cOyd92Fl6fIzIkSu79qzluWyNSmeU86m/NMg5gfGn4XiqH+B
eDhJAH41MN3fJaNgZo31Y+6Gemldg56O3GfMfzm83dLHAeOuXxTf+fsYerlRH4FkF0fs1Tg2lKLe
61my4Qz+EQ2tt4HmX7nXAFXqOMnN+7a1DwmSaSLgJSG/MXVQs2Es47yq6XzE8QT2bzL5fjSx5cNU
373SYCbwp///XoSbQymwUaTen+Jk1Mv9fGv6ENQU3yt+sS4tAquOxa+0IffCOSJ04DhC/symPbtm
/jmL9nj8lkr6eZwNzG5HYu7YTNfpIknApFkUpF71aNxqIt+oP3sewEHQQVExBnC+yQEU+zIumF1L
tOBi9jpwN+Pst/BAot1Ul3jEzvZx3MgltZEcx+62bmlEKjFn4jHv+/H00+IdcYHJ6HdWvHA7cuht
UlLesKv0lZ/02UDL4cokhEnwSKVOG0Tu+qXTaNzRbdTFAlB2yavwLREhxU85PECNsFPoCRuXTViA
MU6mu89ONhtuVOC55TewJr1PXiCh0Gv0fB/LMoRteFHStMcpsrQmoeXEEcngm+B9odKlVIb7yVtG
mBPX4wq21kJc6eEZacKSHwQZk1H/aktXettREGkeJcnVrz85JK9PMJV3yD9AnhRT+YVDQaPNNYB3
54NHnT2y1Zl9xHnHmSv5dciIyhOQZ4fNa2y3R6OT0CTj2j+sTWS5dDk1cmbN1uOtNffN6WX6P/m9
05SlVCdwXjAJ2JcPvuQuzs3OFCxI2mN1iC5saFp4V+iBYwWpzSigXY67S/DUdLBwFkdpWDrHnxV9
o4WsoObR99eOBeky4kAAiQbc3eqHyrteK2aI4HmhBIYZGRPnF6XGkJi/LMtaSccyf7x64x8+kiMC
irgQV345kSDKdrq+kQ6sYR1Gtls3tQl2SjZuW0IEjTUhvM55jEwVI6Mf576GLIruEbGKBxpvIKdy
tctEmvyvHFXrF564jijRAjN1xcNIieE06E8V/TYZmhuIZsHh75po9Dg9/6qvJ1/SOKhUUo/TQeg4
6EtYcb93JjjPQCMV0eFvoggXEVPeH1vi/M96SxdD8ftqhEMwUD8rAvrdV3eCsGN3ILGWquDNnbSE
kTSQNxl3thU8k2RUhLf733JYoASj+bcg0RZ+cc0iivEE6i+/FonCC9KIrIe04dknBEo5Z2CPu+tn
avvD/8uuOw1T+ZI6hNlzGw271jH1cfENAgoscVEksoB+I+zLp3ykfgXnqhcS+rEFHhrX4FSHS4T/
4W+ynrQszZjChzzhOMROdMo+65xgEGfKsO7G+rsqG1x2FD9W+9uro4bGlyqVgd7jPvm8SuO7pUYr
WI+idZA4DECqRatCWNCk60eEsWOWPB0+dimWLLXGDNv0TmD3uclUYOHuDIkUnbT/QuUXQIteZwdp
8KNzwldWtlpXQ6oYWrMJ+oQ0oILTMNfuLDUhsZfmK0I68veWud0Mz6mvDK9o1l+jfjq63FU5LTY0
TYvjKwuzilxVhjplk3am9sTcTQbkqbb9lODw5oeAXL2OP0EBTOcA7Vd3jFKM5rULsOjiHtwtcvdL
EYnZV64Nhejd0al2NVJ6H28s3UKdOIofztSZSJMGnOhTKF0DI07+1fkH/8ujWTh/uhMZTSxEr+kw
s+iBqddZrwrjhyEKw/LnoZoPbKO5IyiPCc5Z8p4/lbL8eVy3bg686WYOHyb1foqkDps6kl/maFhd
2Ic2AWRaQfvogr/RpT6npJpwHPxThWdiJK1p5sv2QkfY7flTAZOGI73MG5XHNc/DjzzJrdkHRCln
qIJOIOj14ZSJyUnqAth7Sj5ll/neKVuA4OlGbuHouGUELiTCgTxW/qMISQqzaDiCGm4nz/QzOxQ3
beJz2LEVI0JXJKvaIiTB3OGIHIuEJKOq5rB6uqf5tbjay6j2F5vy+8c+owtI1tnu99ZLeDfuXY5c
cXRjjkkUx6RK4ggyOZir0UCqBoE58yuEdYXEQuBGMoumlONrWqeuVv/4OVZjcgJIeJmtsY9pcgr/
jDuq+cxsnDFdGzdF8LjXOqjooQu7QnN1pmW5BjzzCFhg7vn7HavJ1Xp+WFvnSEC3Ck+4qj5c1amA
qws/Ih5GYzqS4k2KdepQqhH5/LfRCQiCFO8mntkdj1VI0zSsjCHDUP8oSyVFndHk1EojJYY/bBhO
kC1B2ZdBWtr5d7onHZu6ET1WSfxQr9EBCPd8QmwXrXLWEVGVuK6DpaPQyfWjm+9m2MabjZ2P+DKi
1ju03hput3h0uAgXjcUiG6F7dWYlCxABo1uU+44EcE0gQyT0F2dRMaJaL1RsKo3T6WQddu+mVckH
rpVxNlvq0qQVbDzjLH50k9wzLSQmCXpWjNbKZvbOJoIyO2H0Gv664RcYPRChVbSMl2/3pAg+T21f
HGjDGi6i7HnNAninuvbUhaOULaERy5B6Ge4QbvB1V1H4nxraeND7zAupdbSyiBte08p6SRSmkdik
NUdQbMQuNYTZj/6o46h7PEGBFxYpPKd0hOuGiRjKpWJvPkBn5swN00oX4iyXXUIhsD9gp1GQEGtW
6WSUF6h0t8/kl0FTQ//X6K0oB5gwC5ghbK3QbMLaXE3RXrcd4obq8loemvT0DLAmswY9V0H6TG2V
a0FZqKgfWQVZMAESQrTTwCxImsLq48I2Je2WdemAQaxjP8RBqq/CODaWE5YwuuH9LWlEJFA6WSMP
BRmRoRJAIqAAIz3LJxVXNufEzSrAmNXwu7VW/IX9CPtYh4L1f0b/BBpW/UxKfcKszB3SKoDlK8l0
JCROh6evBjhiPPdXAAAA/afhRCOjgmLfTQ9t00SF3zxyYwmM60xQXWgysgEBWxNC7x7m7Cq3hajr
TIcuvQgRAnj6hOyw2R3aRSa3SZb9asJSFUlhx9G9JefmyyB998yo58sk0QxcSrsQogXCNBgwF1cA
ZbTUEwxWCiPdh2an/r7td7b8W/MppD49wRuTAgBbfQ1kA01dh17p+tSI7u7XqJ0QmqFGP4oXOEry
mcsuMZVrxqaLv9ISiaa/Dyu0hLLIH83RoYq6EigQRldQlVAwdaQMzWUJw6CvZexHs0oJEYqAp80e
CMy9z6pdsxC4Yq5QVZveMFJCq7E/rVfJupHVZPUBFnHTdcQq56LIvhdHqHhtTuDJZyC4eKxkLFuH
lNhr3KmFOK4Ev2YknLnoihK04eHN8fQAP0e/B0emk+3f+YlfPHeuU0ELIFHa6Hz/ns5HLD3owg1C
nZmQGIq4NEsrY+agpx4/DZdo65MoXlS7Fi+Wdw7dt3gUft1i+pgXO3HKyP3Vp+tIexsB2Aorwp1Q
HEjycfnAJNh2xV/ciVQ1cII/UV1bCNdgX57X1YySCZAYANcc1nS2A9vl1Wic8926Gd66Ajlbu3Xe
8VOxhl9k2YrFH02mhBQWCSnqDtwZ/1+E3HlBEXHVL3Aql7/5L8P7lkB6GRU0ILBDgnVmKw903Xwy
s7JMvRPHI6htbssl5H7YDf3ctLL/O9YBo0YqiKJkOAGIdAYuGc09lwqthZuiX4HtgaL3DySePKcJ
Ryu+doi/x55xXdYWc11jTb+JoFJxXQ+F0/DLgQTaBoARwhwryCSp6V2/aSePsEefcOFLQVNtFYpb
1H9crBsC+zxw1LjV5ewDz6NoQStdMo2p/GQ/fCktnBsY7z1kSq9u3KJCOdUYke3So9Pluhrc7KmN
Ti1O3CYKRuqQiBWZOrVgkaPRsIrC8Jqqp8Lm0/SWIerJc2iRRN/LFvanTDwW4st4PFmVrZ3J1eFK
OTtG1DbtORrW4otxH0bU24a39qHcJ+QrBPUU9gId/CxDABxG9LLzWvSLQ7G82x1l6mZKhq60vWMc
HG416pFNSBm3V4XzAYk8h9SJZJ1bmJUCJYXR2HFW3241ijLKAlzM0Sn2hEKB4svDMR0vAKc6Nqr+
OlwPqqoDlkDg6gqkY2w0/TJsSn2thx9Sqw/kkttcufhBbhc5AjA2dDdSvHNJuzd1tAM2MM/ynYhx
fl/WBKr0On/8q5YLDPtU+NlgTrR8JpvEZHSX5Z1xtcMt6Lam/miQNqEBfbKE85ooz58peDbgXU80
yoAgOHHvutYkoqZyM0mvRVO3gGszSws+2rs6Uiw0yeH4iY4uvIrUmsg8T6zKchoq++XfHn+P3epR
Rj+vpL6DF3kpbk4DfwrLJvbXQ+fe0neXjUm6/9DZiQq6uiYBGyFh6C6qSuyHqKaRMPTDA5Tkl9Pt
WCQTi+XlVQPad2JHrlIxNzGUdkVCA8zjwhRUgIYT5AN2jnpo+zNNvJJDv/eW3vFE9gmZerbu7vQy
sLtmjv2fX7sw3niCfQpu+JTrXSl07TYpiw4LX4VIgGcewqkPWeM1bSKMDdP3s61NfLCr6raI78fh
PosRDsa7RowGPacMkhw5lkf8zgjAZyZnFFWAUwzxErVCbka9KWlRp2OFTGcS6p12zW9ew6TgHB7/
7wRwkqkgOGZnhNhDN3lqqEeLykWXVhOESlwE9tnj0wW/OIBRU4mc0Mzkd+xqsP78dcHuhtVQGUbn
bAAxEkAHeiux0wjzLIqjNhvKrv6n0UJfBhNlwSSCE4bjyU2dW8tx2gCTCfJ8beEeTju+hKvT2jgk
yFWEv90XfUJAt8sbQ/+uRtLrND5FuH6GRpdQ3C7Db+l0pMZBTQ1Q7ivKNSucjZuJtA4ypHAkqdOK
OahsfQCvjBGFyi1EhMST54puwH+DOPGsNtqmGh2b5DDxPrGmWQYczU7OhJvdcj8IT7cakvZHHHsU
a8WtIs7AWztBXxDl386ofQheA2rQp4t7NW5a0rHeU6dvciSjRo4ySxxj5K6coC708UG7GuKpP1Hh
pJD7MqfL2AvycteaYimDfw1EP82M1HC77WgKxf5BNuf9iKo8dudSpNGSCfirDVCafdmwFeF11tc8
LNOw/lp7X0jfaMgKxuzT/tKExfTqui0h2uVu8hkzz2LGEtD5+6v+Qb2tskk7QvEXv/FYwXjRlkG9
vrCY8Qmg5XNdyX4rmESzlgrilON/rbNLyzvD+HITF9a4iri/EwMXR85pnIWVkuWysLEzRwx0ch6j
/ouah7qAGE5jPWrSvzepfZ7dYlofNYbXhyyiaUQKulmgtqpF2yjpNVPAh5e9HSkx9efJP0KOCUXZ
9TlxjG0ZwoPCC4G/5ILL69nkvPWE6kl8oHxkfRXdNqdaJ7BEOW/rQgn/Cgc6Kwxg2dFGMu3z46mq
kj7R8ITLpIiFZnRfZdlGhzeg7lTAOIOwM4qq4eqtahf1QZfybD02mf5NnUkVM3bGe4A282Xbl91x
7k7aewd631uXemkBcLXmb7LA8f5+FKTZEhSiTOP+MspoPC/Tc4LDYXAvT4pNTOPXdF35v9J2pHe5
XkRmmEenKfLo0tTRervTMfN5YIrGhr0DSffY2usAd+JjT0j+t+iqnZ/IvJhJmexDdlV5otJi9lLu
OYEKLXQq0GAE4Qj7VT1Qpelct+9XBw7iZKSsCyDEm5BiMtnKHKMyRH9I3xLe+8llYcnWUKHFPHzk
W6n6ExbHIC4jl6l3Dj/sHP7jnFrWuHxJVg7do2JkuGxUQXnnTn0dPIjjdAyBVweVQJl/zCar4Ujk
F1d0Rp44V9eHmqxCW8vRKBeKh8QiBHqnTSVjW1SL/B0FBfcuyZt2+Eglrn3QXmQcXRrjdtmhcneK
AsodBeUTBRmtT/fLHQy6Go5JJAwCpmWfc/XG9YqQGrJ/fOL7ZHkxMAhlbKkn2WMBGi8Uyl8zX0cL
qxwVctSDUrtB/kBgoPWKOJVrtMVz5mna7iaxvafbiaY+DONdmXrRoYBoPdwMSwl6oqbelGS9FMOh
7AaZYUv3lNr18FPJKTXoZCxPym4ER+QNOKjHo5pZncDQoXeNy3zP50K/J69LB8gzbiecslBm0Mr4
G6kPlpnE1aV5L0oCgLR6gDNh4kZZTsvHZaok237F5V9bonG83C2E2AS5xG7l32khWh8nyNFKWr2g
6yDuvLDDpmyHln08oPlQ6MxNZ+0edsGpAT/Cn/Oomn4vUFHvVS9Mz5vrPXyl2xy2vmr62h6cN6Jd
13UD2VG7bxIA6Hvz4ssWbL2yDJUrs2LseoYrypMdso8M6OKcGkuZ0w2QfiFLvMVfMm+1+twy6JG1
GTMlmP8UA8qgYchrS7RAKglYquUGVz2fn7FeIBMbjROY2apFnS1+RFx1V5jSVycTFO0c2ZDNns1v
DVg0wj3vljT0P8eASb8tI2ujeX2uGYyy0RRMGvoUprkb/PdDXa4wHAxhc0/ofbt87eGdONPFMYXI
D5DyhShDfr17r03KEbYgf0kVjMvMHEuCmRnqc02T/NlKzEXtZDy/7OaVXDxMeqZpdst7Ihba9PXy
6eMZby5eQutF8VirQzoeB0mXjsdGzXB0+bkmsxVEJSPjWRzch1K1QmEAdPtuHYHq9MJdv9m5KdbE
8kfRX2dr0nbn6HoIccyJyUv3Wg2m3juECk9o/9nwCCFz3tH83e9hHmxPSH+rPZhhTBTQlu6fuZ4F
k6spCkr1nkg2B6E8TPv/qEAhbarzvDKPnZFcSbs9ojOeuT12U00ibMlSpSkLbp9+5s2mX+EfdsF3
LXs8KlLyS2YUESowgMxb60wFl1qZN2bCt9R4A8WOeH8ixSfuv1c6VIImQMoECuZ5FZgPb2Ir1pVY
RTlmO4nGdCbYPiyKUpzo1uK11ucYXWCpm1DdUORTuKC0hC9VfVpDU27aWsxFvRvc29yzY5jLBFAQ
9Bn25KozylgDD6eS0RoByXJm4+h7f5qzSjSnF6cxfd06q07a+rZtiu7ju0q/kcUdFlCs5jPhuhlv
qe9a4Rx2kEE/F6a5IEyNssoG/mw7tNrQtG5ldsLxZ4sgW3qVw4G5OOiPvGfiJwPBwUh1Qre711S9
kfcYkBY4FmZ7DVQtWvojLNazuPvKn4fNr9EqsmAAz+22SgTQO43RdLDwCseNjcFAwOP8ELvGRx2v
5haqBJhXpACybmgkvrjpnxf7gfAOVhTLHQPCFJwhmqdpBG65jQdHTj9q0xHFvOyPmx/AhVJr1RHZ
QW7WK8wPjAbzsUdO8KNDN5yyf5fgwnwG29661Rb/Ejys4rNylP1FpIfY9lI0RZOVD/5kMBlo40U4
mRosP0somcH8Ak2mZYv5byYIBv45OC4iX1ZumHlyS5hz8jEWysgAAv2gRsPakI2v+GqT3ab/YcF8
jkLQsvjxL4S7+IwmfBl+y6MkeuVFjC8LAhRo0fm85KZ2z1duxmcI4u7lH4DpIfvTITGY++0CXkRn
CVhpXSzq0D4TQRIG+HJo/S1w9TEi9bAuv9jNi/3whpWQWrfEup8NTQffqUonCjN5b1JGXHMi2I4O
dtLfFgoZJWfw5Gz5XngIRRyjeE6GCwc1Ee+H0PhLbWq+NO9nBYWB6AoIsE8J6nHIZFXzKnj0JvGH
CRMvhnqxa7yOVLBpPXmaGLtHAqwFnnLeaMlEoZcMEjzAa6CicL6T3RnvG3purcvujwkhOpFPyt6U
mtd7asNrv/ide6K4I5ZNeM0BPGmmzozDLcroqo6YjGUS8kC7p2a3pt3dsDo1Grm+Tw3rjjxtgYXy
+wDcGZQqtWCyxcF+Ypj9zNcMbSwsEkl2PM+N/+AeeVvSyt5sAVlqK1++gP62NwKKb8IAAm+bVhWa
T990s8Apopvw3kUamQgfScZezxNpC6q+h1HdHlngGYfpc1IUqvp3H4U7vbwOrFgd485Lc0cwtG2H
cSimWDQMFTJyLBLCM4f7b40rkjB92x1mPgya/CmtY9cOCmgrmMF1SHuT+grQnIBgYszFvY6swwwZ
43Miaie3z4KiGDMJM2n7EoBG78W/2sEAcdIj/cwXBcuUjsHcr6LBxh6Zlp6yhGyxUa7E7OcXTRk8
z1EMATg4kDAOXZml4aSHIJsMeAtSkooklYldGlYTy0M8M7rTinFtUYq4HWX8BXjv9rGbp3R6Hc+T
l9PqG43C8F6J0Q/mg2T97yvH3Bofb6N8Nj3KniT9lXG36qruTh9Ca26wauYf/3W1ap+FkZF41SNY
zEhmJyJ2oRO0oAoi5N51b1ULul/pE9MKS97CY+v7A2lIC2en2d9wcwOy1JsHcXu7HbvE7k46Fyga
9VYX4UIJRg+UkbPCSb/zYR2rugjcQQf09RT2nV0ZhNt536TpgY+M7PuRDDMLxbOk7ftCI9ankLmE
p7RDfqTvRjSjqY4uNGhYWdN4jd+AlVvuuCEeZX/RWVM9TTH9SoAsJiWTa/YA3IDIV8B8Q/M6jacN
6fnYTELScOQ5VJh+xfP+5L4YHBo130zNX/oFytW7X1xLozVSOHv4K2yNInqvNPiIJzPejxmFUHuA
1B79REIcfxJLTjYIRfbQd9ZSufUsorPlHuzlaqvPbRtCHiaO2dsMxpOkEz2B9aDRW5swV1dXBadU
yC6dy/eBdNH4oS/jkM9/0NVLfN8OZ9PfZIAY8rfcZ03/pdftVC68nmYP0IeQDeMWY5kWBWx7PsZb
YeccWtBYymzwUVa2o/9aMNz9EXEI7gY3m4R52O2iKx84jK1kA0c7YWuk44HeQikFZ2RJM+ViVrZP
deQyL/HOGVTdJ5P+ieeth3rC/6Dmqp0xCXLt1+iCn19OORI38n8n8KuEOFK5DQ5Cb6lbPcjZidM7
55/G+VDf2viumH41+3H4sJXBGnPgwE47FkBPeSccqrK469v6MFnUvl/c+aERxhdMPnSTnUvhudbU
JIM9yMZslgm7BEHhk5HzNRCx4FbxW4UrbhrACQJmrmZIxEzTrHHFGLvaRgUhbwBAWfov1ZGyGNis
clWaxLz612O2690ZqdI/C6h/F++T9XlB4QGY1pBUZnBP8I9VZm36twk87pkaX2qjUhGY7iDVVJtw
qA6M902eIh7PdYcSQ1bw8kLMHXC2/GgDFTK3XAv9jvkTP9YVuZbxaGdMEwaJ0w5mc0BxBh380Tbd
6DcVJCgtqy01gTfw1+CdxhPGgOuqpIH7Qf+rsItKxv0tpub3lKD6xjZ9YSyyYHkeC2+riA+9tz1Y
nboieF+pHLCPEhs2jsN905lUdgD6us8kEsm9zgYnoD/jrCSrkpMG9gEq+nbJgruhVEoTr32u90nw
5956lAuOTt1CWCBcDACvuKwzJimZ5dhjINIFX335EWUG3N6+4aB7iuiyuZ1/4pyJB7cgZKTospqD
wpG2ZKdvYK0Tft5Lnqx2a/32ashPWm+EMJ06oVdBTUkb7TMDnCBYB/XEeDl4nA8mvrUSnHs/n+2r
h6l5p7L/NxVYA78ooukXDAcmyQop0ls9WZe+TX6CuWZeC44jzOly5yDL7F6Z+WO7GUxl6z1gN8Nn
YMJ3uQXIGr0HL33BX+g6D9c85mk9huJ/4U82n4N4HfH59XAeykqq5+B+7E/ZG8I9s9JkpIXu9QPR
jnfTxnvqfwrPUmQ6Gqs1QUF1R9UHm3MJpadlmgpB+qA0aEZM3DlBOMWetEjlby7gLBNng7NNU30c
1dRoJ05S/lEFd/GxH6as+8XnyGb70JuGAgoiiA2qimgjU7KJCuN/6r6m5tHXcsb5/5u4Qro6LXt+
BrcwwHK29CdZbBh0ct6oCi2JYyfPKfhOldjHR0ldHddV75ZGlnBcgYDJKErFbUv085ndfpewx2/+
QbGLxp2uVHTb+FO+1QqY1pT5w1yeeMmTcW7unuzvpATPdvgWjr0zYM5AiLHLRVdEVaKyUa2/BBYd
goG/6DTiN3d216LnGrNVhf5X+QedXKwaMGEGuAAwIVV9t9Ag6HFaCE4dZVUv9HPuS0jLkWiZMc4K
puATgDbOPXt+CwACvkJb89hV/kUijd9mqzP2w2rqY9137Uuz8B599q12UcBYpMhGFa/fIRHB9rWD
ODLF0Uphj10wVK7qm5fMAFHEejs3xVKiPG/K25fI1YdX8cJqDMCqCDQ/e9n1KKBckeYNh6rWf84N
VfLRVP5ABpjET/YTm4bJ+a8UbVnKHsxc3xoDree5F+L5CmXZxYwO2JWH6Xt1B6m2OLiVHahbB4oG
vvZ9qWwUcOt+ZfwaQrEcJJ78XIrVIFrhPzGgSm4hz84JnOjAalhaGtLZtyYTByTcFQZ3+KUjWIb1
kXRJXmzsAz0D2LA0HsqVxYh6/WP8E83labgge2QW9kMCo8kg4w7VRlKHui/ZDwIYDntA30TF7Oe7
it5H4BnUlu9UGSB0jUvvujWl41L06AZ0yQv8TTaD+lk3mUiTzd+uxdWEDWAhRWvEIMOVEqhIeuXc
zWmBC78SkMDUigM3c+wVVncHuwD0bCxty61NmpElGL5wAKO/brBtldf34v/7SwIt9uqWhM8H+xY4
imXAoGpoEPS2ot/3EjscxGJzxB3wbDEC8bKGWIb4Z9Q2viuSTAq9MEDENZjDmDVxa2W+n1dHnSXZ
rQdMHHMyAmMitsNHXFITLt2ETcZ63QwEw3vEWCr1R439SsY/bneBqZYiJjWBbpQ08B6U0+nPMvb5
mlW/wiAlLmhgbt9fq/NRX+3a9HW4EBEFN8KwKmaygNa+pZgxioXfAGFavuQgcVhpH+RfSbc8F1z7
pJ/tsbVByEsSmksr79cO9n6MxJjIsX5IvZgh4pBHX+WkoqFlrRkiipB1OlR+zfl8JIt2FGBvjFYj
0GyhXoKCCK4xN2lwrDfzWXv7gg2frQD61sgXMEbhegkLdgqod3sxANn8tR6uw9HJFE9f8NL1jD1o
6dIAzLYoOWY+yrpaOQ38/FrSjKNptCztpL6WihO+oITQ5el/RqfDagXs7LXau27lsjlqorQBK3Q4
UhifvRlxzt+KPOkB8XVMADwKLdWa/f5RylNAuDQk5x/PESeX2Uhu8jisyyJ44WBFn3YP4WnVm9qK
x3a0wlfchRT25w5PRab+Hmubm0AT38+0Naxa5J38slcf8WhtkGHKvRmkrz13rba71Jel74TrAlIC
yJl3w0HwSXc5UfePQAZ4fGxwKfuz+fcqSyULgRn+/G+DNDlygIz05inkULmO+mnY0hXmtFr5hUcY
GXA3Fu/dIc7ZSOFeKhibzfEp41RoPFhMIEw/OdBWLENZ99YxsMf+Y5QgYPhS6itYhJvfNm5soCeX
kts6SczAUDxDNRoMR2pJ4kPTic48fO54i9MZsTA83Rox9Z5RwiW8buDezHoJ8dNMq3tT0S1m9Ozn
lt47EalDnYsXTInqlugMijXEcGC5VZNwEXlTALmmqIvdAmrmnP2O6cUZOTLIxttjkpt7pEbRPUJI
DnRsoowuyviaTwfIDIKpEg15waIBEkK8Jq7Vq1P+8uFMJtIT7YNnDmHKEEKjJL9oNoSkPnpMtBCA
4Do2io1kELeBKte4GPhtPi9pxQhATT1Sw99YF9RsrULPDBx6iG7qir+39/pD4ioShhseYExkj4Dv
l15xO9LgosMCax7YdL+B3jS/zH8xylP1Gg3tEWx+aDtOvFixTZcoRrJ9UHh/zxtKgCorZPjcLtaA
ESNBF9o3EaHE6RK0SQGUza0JfSShlQjodW50o+r3Z3VypGw0C570nbGyy9qhKWgyQS+ikc0Uz3sl
OUGWCAcjKgL/Sh1nuAy876WG9gCzYzzxa3oNK44xT2MLQgPs9o5baEOGk+Ihoo0UFrpgdFgHY87F
udqA2n8Oo5BSOzWhv1rD+yB/KiDjMAh6flkxOA3HTTpHqhk/l2kXqeCdBovi3Rkxu2RnMt4tUDNL
gnvvDPKQlnSDDTzi/eiCcqcQBZUGX5JqimrFtmeAT5qZRZN6d6FGASm6DnosvlDmrLR260RJ+i1W
K8gHx+GrmNEFaAD7nmhl3elJnEJrnMYjADh9ANdb0+a+jUkWcSAJKJuN6OeQOl4XLbkZuYqwqecG
EpKcAfgru313LdfH0uJLY3QN8aHxA1fS3AGjOIRwfo+3+xwvs48ofHcm+UzhRiO+zuBLsSn3l98j
AfyO0sk4hxYLwStAH8kr43iMXzonGbWG2P3B6ASGqzXdmedhsJBO1o9iI0ODqUtkWZtX4+G1hQNc
Dqi1CaWtZFKklbdaAKDamXpjrHaFBocNjwPtcQgQjDOXHuBWzee9v/G1KGhMpPw5zzCKFlroF6Fd
frlMuLiHE7VMst/G1p/h9riBwVIJ90GFZ4e4nWqbgncBMrtswLarzfvC6Y7lOsBcqNVLjF3igWlF
a9Xc1YQ/DuDEHik5q9yhbqesODSOwaos3w2+jwuegoBGzyE4wDdXutdNa4uQ7p+EYfKK3hjjfegz
+5fa7U5CopHUK3zmQ7ywdoiHGI67IEid0PqUZIwKWIngETj8jDTfUqjx2/TAIzsPE3iekrNS6B+5
J0ZQlzgNq7vYP0eOipuMdWX6pgI4dUQlOwvAX8u8mgocDRjB4XqgLJpiCpu1N//sOUV5YjgWKQUU
oMH7FkeA/JIn+70x/JsOwTRKcPdlJ6+ynYpBQYU5BmBOq2R0YRSHkNcrSMG8X2M5rtJhDQqUkHIS
Kidy9mt2bk980QjXYKem3A7vrxj8EZKWhJQYstcXKRKQbTdHC/gmt0MqT5PXeWd1vGNloLr9rxUg
8JWdDKv+hnkMO/5x595zQWhaMwPxjfPaivy/0hG/QcUBHyMlRalpYkIiUZ71klDV0XJRGI90iQJx
FieRvjs2f6JXyHzrGdJTY0JxL68kAHUK7HUlBOyjy/PcZ4aEt7TpnO24V7IjNVL/4qsNPcU31bms
l6Q9gUU/M5L6mjfY3LWVOKfxkwAqcX6Gib9EuYezzo1T6m7PBrMWrgeYFGffn2m3FkwEArQdZotM
IauQ4upgalDMDmIUi6YSD1kvZG1tpnMGL+f6FF/9X8xskkwOdHUCdNYQuFu8XFQbC7h9Zi3hY9Wc
tbatAc/Id9pXcHvqWHqfOeQinnJKZwx0pO353/XV0LphLPaLScj4Ta6oTGP64Ypc1huwlkyY/FZo
r00euBa9DkWXzaOIFlkssZugMhD0Xgi2Vxjp3dyejgPp1uO1heEc1qGVnCWW4sNaoHVk3L79FVTz
0sv5QLbDIgTW7K7rjSs/HENmOeeH58hkoaxLREMnkIXuA3XQydxfCqnrvlWxmwJkQxCoJN5hjwvC
JOrp/qPMlJsD3k1aZgM4rUWQtGVL6+Ldvv45uUisGzx+a8bBmUJ34FPKnt9Qq6dC3w8x10uzQ/VU
vs0BBkSz/VSNs/lcrWaR68GbxOwqftrqeO+uPZ5awWuCOc65YW03QufQOOdU00cSSgG0GuBOfF3Y
JFq0fcdro1DsU6WWjFjp2SoOaL22XUtkLjshJcznPZ9FpuTLXCSIusUjSlM2NkGKHOPgktOZPvUf
I6ZhjbQDqSYlu2w4VVXL74MW+ImP2YVThQDT8+QhqNc/z9D9T5Ct107AgwoMkwPH/u/31wkoeJU6
ZNRaGS/fm0gegmFXQnm+LkMbtSjgeQJM0b++y7yDgpwnZX7ybRX4vKQR897Tvq60iVNhPczEi08W
SjbDoYMaI0xzEP5xr75xcwabPIMjdFNOj3B0ZzUJHSJEzgBFnwjXU9t8ZQ5Uo1xwNGlaj/bmhhrL
pzRz2G7iXSzR2aQIDvpYHaw1H78T1ruSRtKi7ZC2x+Ve6FBfh5SfAQZXdJZhiFujbvAD1tMB/MTA
n0/jzEosHCwfN/rh2BqHrOkUjg0QydeLdaxqmql16M5jXl+/ffqnGJlhUzC7W3UC+95f+fE4YyMK
j6VN1G4sjBv/nsfU2IPMaMgjWCI4KjfnZ8kv5HIA7J79EnS1BYRcebnT6YmMDp2fozi2d/5XMZ/H
Lev1ZK109FBxEexTwv4YUxZ2DE+MZm0dBvXvL932ETnU7FEivUC0+93qX5rb57q4t9Q0RpLGCmXD
jpZLQTwImY/w9Yrf/WcatE+lfL97+I5cm6G69BQvzhnk0kxUTYBA5MKsa65ydDGobMp3iRDH4ZWU
DOP3LNgk7QF1QO0fOVcG97nKcjzSe5520b95EToTv8rHyZxNoVPtKTZU+rVrUF4W8fQQVWMKeYLQ
LYwTi3T0TbMXY0ajaoe8P0T2kJvBSLal+5qUJDXOmsv4q+4g1sYk7Z8zFLrbzvAqrkUPeCwWqn4r
YjUlI/rPkGsjPTrz/uHKM1yO/PpbL2XV+0DtAkiWUt3rurTGTHYK37rURa80xmRotGYfi38D+zTc
Qu1ijOMW25mdWDSW8zfS7ocGQfWuQ6RD/4t2G+nWR7zLgs1xJ/J3kWfkUaldP8MPIj0WEPBbwiWd
/bBco32PhBalhfPSQ3LyEVLUeQXVmEElCxljPVefsAxqIkCdSGqURQsBzZdNnBTaqgaB9u57FamV
iFJ3Xn7nIL7IxOGxYNj/RVEINsWYSn9nOW45hY38yTT+4BkerxEVVKl9fDaAmUtJkZ6qngLVGyRQ
gCVo3xA8Nb8yEmCDWuzgk++dYcLZTj7O3UE4pp7T9mQdj3EWgyay1JJ4AutdQnp05pB3Yt5VuPfP
zk6uUVlJDI/pQpqyQCaWFe1ojHdADRdmcXY76M5TAPChC9I6TOgAjx7adknV0YxD7H+30/IeeA99
TEW/xu5udpmMJLc28lipPJTmvkEBrmXXQ/AYwRaMdtbRQReqqq5Pgs42KNG5CbtwKqAzh83lBncA
Ee9WwwLa2P24ttq0ZRBQg38KgeL0JHqZ0sVBc0hJVe1IcNOct5grRnDymtioJztV3/TQx5APeyqP
Fx5LNILc7ArnoszYfVLskwdBkxLj30ydHdDq+zmXa5HiNw3fmRf9CxFVsQmlJV8zTsjQTlAqCGix
xXL3nsgCu3jzLK4MvYCtmdkuj9ajdbN4S7gsaGsyP6IjJiLbCgA9Dwr41qPL3MBBOTtIluBVBeCp
3BotlKm8NvII4YHOLUUV04XTu4b+CtZXdZ+n/eR8l2b6io41wipevi9X737iZjA4iV9Vj49gBxKn
DQQ5hO5JjpGqxej7Y0oVa15R/tXXQajwbAWAi7+CJdhxV7kGr/7NZcNcTGeaDzfjHHXjocsvapM7
77D3WAra6CDHjii9NoPwbCXrYvT67veyoz9prfhyDmDc/EroV6TtPf8e1JfNZhYR9RYCbyHQ+qYm
RqgEmMvPkbnQubxJNk6943yn3/MWsdeAGBZWCCo8tGlludWaOzl/Lqv5rCyvqVfEUEzFZdTUjak6
gkyOUX24kZ7AqtZps/yIQoe7sCW8VYrTlNtDLLOo2McF71BYAG9bB8FU5ORDtBHUOUnWmdiIAwep
gg9tO/wH7OgXyHBiCHFzRtx6r4qeQ9GmR42adsgO4OfAkKUIvw4U8HoIhv8nLpRE7emTJ3vRgyp7
MTXlnG+4kUnjlxL0FY0EDUajLOe0c08nd1xhMQMXft2VAGoAYU4mtL5vcUuxwpR7gvEKKjECN3qS
R/3CXZ4tT9N3vGhB74Oig/faPDshJQAF7/rH2J29HGBf8qxh+GfakcEORU9P0l5xt1YvUOPJUZpe
VFG8d5Q/8li0uJIpa7h/RC7YOunGtZ9COMPDv73xHUx2Pv9xylcEJjzQ5tAl0kDtvhkOXLRK17Yn
6AcW0s9VhzcgrGRUbhfzsSSZQ6Otqz/DdvLWx/ETVNXP7MTh1lZ4sS/d3+fbuMMPJ+ksEEPFd63M
E0j1d/DqSlUUZW/Etf0S3FQHJh+RfhhfMJ77JEg7XJzr9ZccpsDGgttD4sumhbHUIZo+PLrsxgSb
kRCOpYHln8jjNQFj7IAiWCAkcdOEEEQAu0fvOeXN38dalncxg76PM6hTe7t8IUzHDHrFLQCb+IPp
s0/I8kJfZU0inPnPhSYD9LcBRDguLnmRWobHrScVYNpmFnQ8w8O3UxCLWvZAro4Z4FGhuggn1TbI
4wMR4pu/Bz/15WsfDhoAZhkgtOdSC44/iPXGTKDX7Lg4nrf+p7IFVYQHogz3FR7ufc/fC3qvA+e/
uB0eayKVBczscsbpRQUGHZqvkdHw0y9FCW7MuPGd/rSnVv9TwFF4xUxVKhFys8OSR5TZNY1t+XlZ
PHYU+K4QZ1lHwis0ztoau73rpc+Kk+B+v8Yxowu4lxB8ZGTtkT+gaX6hh+LrYTNsBn9ZogQRpkni
T+QjwmAtF2XuBnGHlIgTG3jnRfGvd4ctPvtRRHpf509kqKJE23ZI3P7kJFUyZ9eTdbJplXIZpjfw
nhvbToBUFFU/Am59RZYuK12o5NqZ04Z8Nydy4CxHZA4drsz/hyNL1Wj0VAWS6kQuy/LTGRlXN5ZF
4QwOwwMcWn544wsdqsIeu+XW8dH87t5O8AeiBi0moZ0q4mBuMcwNRIE7cjQrRiQOCx2hRrnKSKMd
cqMe0BsdHuQ4T4FRsd5vXk45DOEYPSVen/LeywVP9f6GEFG9gK65eNzvbbvyAGv7DBLNTXrouZ3D
89g2wAuvBqAJnCTGCn2PXha0DwDcGG8FIlyqxc88DhO4dDxbt0IhgnlFe+fEaZsIgqgf+1rKQG0m
ipqgaCHkqxOHYGFdfn+lpC4QwYT3Uqk/0OBAu5duFNHBvegIyQ2ZAdqKY3a4zyZMfQqaLG78k8/e
2s8sACVtNyV/XWDx2vl1g/fj4iVPV1TvQz7ZmrrLIevSfjkYnElxygyYzxvn20OjaOcdhm/F/Tyk
/VeSzrjWDXuJLH2eyFJ//B0oIPi/TxwehD8e0BBmueVR/B0IQoWrxZs8ppTbF07bzmHUPTfuYAFD
1gWx9rN0FTbKWdXrL5IVdMDWXfKrVn9ecqICsv+ZDlKMiLf4dIdxNeQJEFiNtuxbIbxt2SyQyy6Q
4XHJYDKvOLtbAwczOseCsvoyrqNelHuWN/kIT6cVS2WVQ64s3EPY+bY2MN2luKzVOJ6C/9Ih7q3v
zvsjg+dOnkiGGSfOaICnuFdpL4zQY6YUo8PZC1QAxnOnEPsqBOL4IQaLhfKGS0ZWy7htjFEoWUV6
Nxo2uCAMsaOE5Wfr4AcwFt1FKzOndNkNUN6gTokiUkuQawsrtnGH6qdOf93RZFv04MGyI0vS6LRu
18Hz83k21VUGN2ULrxpPj2B8PS5iqkzBI54mcFVesMIIdoKoeRQ+7aaqWns0lOLOuLZWwuaSabjF
KGwlAsra0qUTvirs1iZiqAPGAx8zNycYMtD+jGQXbcyJOxYydkVr+uOmmh7PD4so7xlF66Gpm6Mz
PMTTYqIN8TE6MxoXq3/g8yAhO9yf6sqf9t5Iwjv6pmHHzfHoAW3Fq1wjdJLUYicu7ezJVOl7gtwd
CqM7W8v9QqJvGwEQEXCXSO+Cp2bRj+MDCKssJpW1A6FB3Ltczvh8wlV6DhXz3dZrViogKPeCHKTy
N7WYHtzFrB2YmeQNrE/CA2Es6rzQlwyP5O14lr7GtD4ZFk9Zd6aW173jazkRLRQFzFBVzFze0iyp
xSGjuh3UBYiFmO5t9kKFu19dLTRS11iNvi3/umdFxY7e4SkUKFnOcx4/rczvU5q8uO5PrglSzTiX
q13qnKQ5w4i+xgg1mMckwcPbLfoSGKpn11SJRcWyB9tRIrkx8y2M2bPuEKWGFUTrgzChHPiAgE11
nKEkdNQdqphzCYqcqcapE7078cvAjRtDLGndW2lyiyjCOUTKLnuJm6xU9lLuPuk1DowSMDVQpCZB
240tEf8Ji/G+j8Wjh77W7etitXFE0rtBOPps818N5ZY2dbUjREvpKGEab93xQrlzUXf7bKdZBGM4
3duWW5Tzr8DBp6RQGQCXJRCGi0I2hMRg/A6+1Ifgzyq5njFp9b9e5G7gzdVFHGlwLZRJxu2aPjHq
rFSHv3Cc7eeY81vIjrk0V+C4yy5cHrP0BRBBC6LvvJ3Hoog0W8OKB8qbG1YdzgPuWeL72ytUnnNL
VfqStbCOSfWdGyhBh8U4dU2EkYwG/QWYdgcdBoQ0V5I/y9hDSkkPCXivVFk66uvzkM5jFTx8juZ9
WGEYr50prW6GKLXDl1mjo+Wyh1y4ugSCRybmS9mdy38jSbQ+gp2qORi+FMB7+Y32oj4kc3Tx96eT
a5X3mRrFUFCKY+pNYUg/xrwfAqn1zjQG2tuTcW/+Fw8LN2aH/8m11A8HzWtB2dJt8L2O7G2HQAHW
z+9PSBvEVJ6bm2MQ/qdwwGX1lYCL0vFN1qWKZkz18KnD1HvM4LqH5UUeMyLz9mbDzHCaBuZoQWhr
QnWnNxVnXG0+oUz3V9yHsLHxKyYfV/CTimnRafRgXbjUBdTHXdMt/zQ0pm7ozkm6BaqQSOHQX8Mi
FN3xDuDoNtaFcX8ToJyVygVvsEhfT1p6Da6AEQxqUAE5Py/nYWlJSSXrmvBoVa0Q6YwdC8imanyN
9jQlUX8/Uk3I6gw/f0e1ugXWQmv0LfqQ2mO5He04ilcUghoD3FNZVBHxkY0k0sGp90REpQMBH8dg
hUR46BNOj8C1vXHtpYMKV9LPRzdq7a+i56lV1pzipyisuJRYfJIa7xO8ztnxddXzd/ncZo100bgZ
Ir1l9MvldbZliwbkdn/dqGsL8NdqdOwKFQT6bysyGcv6PzzlSRM6Q+aqTJud6ZAZeCE1kQoeoHwy
xWo3gFU3psp1UdkENHOmxBPq1/VFaCJerugk4hjIT0c775MHGdCVP+5WNHQfortgq39mtaTLjgTg
dqHqjPzmcm+aG5+SK8uRu4+/9Mce12S2MWbekP5vJGHvQucYyyxaJjza+LAbSOXpDcA9Z+ay5xVB
4rXP/652TRglCayU/tLLYFbWmKkIsYN3e51fpQbhyIHatNe0kKVFm9EF5ffRvRiEFg4sIJKdm3hQ
LBYRUzg8ircpjQq8Vd9kK5huwmlP0tW97IJrp1Equ3dAlP6q65p7X0ha4SZ2bBCGnUh04uHEFR9i
NghhzCaaD9UEtZH85GzVEet8ID+72orZcmtzzMmsM27tq4lzKpDAMFRhbv2/GNPJN463i1MjSm6V
8qtklea2ColK21Ee8uGXxR6GyAiS7naDewNjt/PcHtpuA/VxgKVKz1q5vU97cIpeRA1R/AWkUf40
+2PdtWEfXsgJJwo9ceaPciTAxCVpjqzGIXzjT3mYQuRXWEPPOE1JoZY6EMYdzT1l9fLX40vO08DU
vOo+wVdBCxJIfA/zcMBzy/9eS8ltAxgrSWJRYWxF2sUNM5/WZ5SNoGymqWSUZeW0dTPTQjf96MIa
tPS33LSTfwr9oZzc8CLaApxb/esuWpszbA6RL/DlQrBkPUtR6fa0DigvQTdtTplGZKuSgjTfWRj3
nIY/ab8MFrAYij5/KHiBOsgAlW4A254eUtJzsMWodiRF1sbbYCPubJikagPQPXuXyZXOT2+HMAHT
wMCJzwK0DDn8xJ2lCtDVK583Ne2boMXcdj/cT3JvzwSJGznt63hlDits8SCwNaAxxW+AIjBlIDVD
3uf7L1ODFIoEzplNtf1m6meROS6GmE+Li1swfUT/JnuFT2uBVlnaNFp0FcoL7F6AjIAwirgVP6rT
y26LxXfvLoXaF6sp7qYVWErDQfBuikG4T4LruiyvaJAV6InE1+N1mEx6S/Osx4PXZ43UMIqAwRjq
HYxnOLtNPpu/7GWx/Alf/qdFqgwzth5utXozut3GGSydMRNO5IMhBMrx5qV5JfDUDu1U1khyWKn6
z4nUWJ5oucatZMi86eqB912baWuux2HLR8ppZshBornExXNo3jyAOYdFtbRaPB0+6IigpvgfrVdG
3bh9qQ+brQmWRGBfXVfajstTPzbZDJy9ntQ6WOHIi45E9GSWca1aicizfm5AF/h1PJVYr4L4Ut8G
jHooRIavekkFPwjL7DG7t1PU3cmhIRqS1cj0O8eDwC8CCCcOI28CKWwY47x5VRqKYOxvWmQ4+1ci
GaKIUk0twpbbtEpRs8p8FKnxNTDGiuzGctEYN8St9ZrY+QhIHuscf1UAvOztDa0b146VGJ9B77LF
yZFkQf/qpwFsSi5tslr/O04QRJk8z1M43aa+/Aud1S+3krg7k/rupWwOHH21pWW12UKGrdGacZjj
fmYpQw7M2knu7GysOAY26NEOJi381yPtO3Jq2oePBaW3dSQGpqRs8AnkUY9MBPeywNGYDt3h7i5V
yIuRkb0V+gqe55M8Bn+m847kugVYwid4qwTXq1/K5z+QNG0Vm6lXLdAE9Z7t7YMiZ0x4lJrs9QFf
jPWTLYjsbJOMZy0QyEeURhjplw9ZVFZMwo/txMUe9kjzXgIJDDqZAekvWhSYLUrmn1cZZWTjt+iw
KHHsCp3+p4S2C6IHpoNb1U2i8fjU4pRstGWQKiNs5FwoC7efW2KuH9gmsjxLj+m0BABVJF1Z3vh7
IOEj21egLFCoAkpsry6ItJYu67+nkCg9ejrjTDFaR+KkvX9ZcVu7gNIHt80uopzFwNf1fOo+6Dit
h4O7oVv5xkuIvSziD8/cTdjCdrELJgZAYRtjJ+Guj612njHbB6QJ0KBcr5oj26uuB6KDu0UHDHyS
3hVDd6HWwFyIpfJFF08f8QWVTABiF7ERKscq+/sDoPU85zPzheANtXkeYM5cTIIult0pT4whT1EH
FNvAgdnD113yyZjgLTLXlRMgDFkDJ+BAFduGeodTPuiLEMgnEre6mIeyiBjTC7BJCaWh0zbrcNRx
5ClVyOQ+zM/wq1zjI05AykOJH31gKWnceqoeC2AbX1BloPKihjVmfkHGlpz2wm8tuiFZepsC7EuZ
E8M5wjTkHi/x1l+Tx6VMrZrvsdC6Q9fsJsgx2G9nPUh1qrUeBbbZLVoCEJ68ZO7yXu19kwIWTSPM
Hm8jcwtGBMKnxUjgK/MuaqbK5eBJNOofpNKof+2/tKunPI2wnF3YcjsAOKtczx8wmB5Srzxxvh46
3KTQqCBRKWrAw3bw19Af/4hrA7GAo9DDrrsG1c4c9iqtdc93Ii6qz5LwAt+UTkMu9q0qUmxpkSXP
ZJcXZB/+Paz9/wRFmKSPURcSTc+yYRfcaLni8JQ4yvlbYQ1ex7VFF1buYEEqVeIcaOWubkh4xFt1
gkvLHl8lUw7yLRHHC22cKyaSFYnF8rKq/riQ/0YVfQOEesjsTIHrg5aYZeDt9jSWS4rHfPsvgNeC
DOwMIHvtwVbyamyurKbkM9v+OkvwDhZY6b0lCVTsB37wgcoMmpOKudmO/uNMkYfbLynT/4HyAeRN
ZzayRiU0owmalQb1LqXgIThPYwDaT+KeMyIAcfDMTHw6diq+JH8R85o/0OA7pxo2+FbyNaYq3cup
DoIlOX+rQ1EJ3NjrMQ/MSUWx8CIPp8krrXOWaIwRn5S7KUOnoRROg66OVKGhEkuv5JDqUWsm8bKw
b5bRklsUSJnynCCadSD0l3x0wKlvcR8k4hBBtfpN4P6Iv8Opgkhmoxql9Y2IcQqOe/Uig/DA7rNj
u8e9Wi+FkggFhsONHyxUaEvfSDz/WWDGTUDkeSompTZBUvGQuOuDCMSa82m9kUzb2ED557nE81aa
c0hSvrhBVHhnQvEBt2q6MKlLQx+O7OV1jdPlyWHaDTbriQD1RuGwNn1oNJGVZxBgFCuRYBJQ3qIS
lZyiAlyuwgEDaeLvNsfF/qoZMjXgdv2idzwbbUOT4oxKlzFyc0TAVUqADpZWYDtnuC2Hub/+FI2M
tA/AK2BiVEyP2l7ZmZ4LwWO3joDRfuOD8DdfavheEXqmJYXYEzRUwJmqiD9RjFTLUa5NBgnaq4bC
oFsT12+QVdoOHb8BFii6Q8f01iY+m6dHLMnoYTpq/Q4sard01oInOIccQaqZmsnLfhrB+4C1qcRk
n4VXByWRvyrYD795bg9YxeRjPCutBMc3BFA6ZjTiT0gIFAqyBHgdt85VOOWEMcXPnbZuwusC6086
fp6BpbHqaMMbHeU+q9GPazUk/LSf1om2/cNvkY6jQMSg6Q70UUkWAvH2U26kRQFa+NTrwbBYsS9O
h41q6XiRqxHPSlAdjbjsisaqorxmOTxiYzIE0iYvLKh5x0tRgMj1hRJXX4hftEH43obgPhil6A5I
G54s8oxNQyKpUb+Z8vjArnK9x1xg9BwfyQjGeeEZ/F+HKIEiX2UHHNEDn34qmR4ioT6cYW2+omBz
3Mxh484ung/M3w++7Lkf9K5Mig/nBPG9lGwyxPyhEq/RvQXAJ8GV8kUWg6KIkQzKct4IuHERPz2K
zU89pXtcuuZCY3TcvpB2WTXe8UJgE0HubJxPcLQlCQqqPqQ1U31DtAyZCt79TcvjqeVfUNcvCnQA
8eNr0ZRj/IQQTtJqUnPGEPxiuOMVTNQEHOoObOGUO0UsYarfv7Eqdpy1u1cPDQt2aeBJvOo0tbSm
uQ8NkRmG6d4NKVQpZbOc3tsZCZFtlh7H9Hq6cttwqETZhIpU4DHjIi6POsL+4ThUycFfKqfg9vMc
Jo2LEDygN6RTqWtaMqyibO6JXnK0qIDDlr1tRdiZJYu8elI603+cv0IbnNk20SqsoYj78Szte701
jTROFaVlvJEhSauzVWs6xw1r4xfYU0QVtvfUsP/7ifbgtKqphq8y+iSLKTfiGC8ux1hftSu90YSC
AlzbBxleZ1QNFB4hzsLpMWm6AGwGCQ8D98dfA2dq1BGBNJcI2SO/6nI2A/KfwCbvBBfGNbEa6pL2
XUnMcaJpbwIfJ7NTrWq8Ks5wYJmrDsYV7nJTVd8jTEPfhiSMsccEX9Sa1E/54NcLyQ20VbWQk1ZP
z5HLslbcybuqYSnjOAgSN+pXYxBQm/XozJcQhK+Y3d8cNauTDHJ5JeCBnjM40i8fhGxfyK9Xtp67
SShdGwn1yf1RdRoa1QyZXWsXUkXlIBSsaUwalcTlAu415FywgUaSrj9sUEmLdKmprNfOlP8NzQ3i
X3Tpn7v/9T24kuLwMnfsn4h23iQ2w+l07h6bVG75ua006kKCMAmIuFr8XBz9UyvRF7mNCz7LqNlF
qP0LFB/engXSSGz+b7NV3ulBNH3MuIvOmJVyZaNWwor4dt1PNVPuSZ9A2CVoP5KIyVhO86o5aOXQ
1K0FC2hOg2WweWKy6/TGJociibvko3YrCJAezDJoM8fIUUmmcJ/mfVg3Wzkyy9/Q2p0msrOGRsE6
3kMHa2cofu08vPKIMyiaPrJDaZ/VDLd0oK0VS3+S/BqmQsAmuxVAHlqiVo/Rc4LSe3jVQsvQj1TZ
C+fiR9KnXB0utGYpvrYBtql1uuovdW8AIRCmdTCI1q6/TsQZjseudhrEq+cE1IecCSswCnOqmEuj
mWFixqtYM18Tyqvho7oH5RqA8XrF6WXmZ+l2D7Ru1W0IcDCWAOp8WiCz58vHhxS1XuxbAgQBZaMS
FpQWfhm+WRKVnJ7iJaD3OKm6OicJ+xXrIbzK+YA+17BcvxSyPRmyRAu9HuELj8sO+l+2HTmla9OT
GL/k+gcKwCaUs+YB1kTrayeWCnZKQEBKJjM67Wjedt5PObA0ID1pqEYvc+zLSc5ejadWtcEo2KMb
YBWM2O/Eme1oyT7WiBTOUu+uAossXaZxiDDj0X1xX0IyAwYYsGAJDUVlkB15jrWXWjoTgbk3Weu7
YgsvclQ8V8iI5ERK281dGEzuxI5HexbL9O4TuWH9qKiMSjlcDpqKSfm5DtAiDnJD/NIJPV6T3CVy
wSB6VBB37AVHxRSJV4QwPehm+OSUwV28/IzhWoKtrIrXoIQSUI0h2Irza1lulAwTewuq+A/mvv3e
475biE35LhUEZ9r91XiNeodiZB+1WHy2xd4lj04DfYRDg0hFrP8c13wK17vwOrlaCynnBCr0Vu5B
U9E6MC7p/IyFNZUgOsBtOxdDbRlr8UuP1xSWoFNaBMECA2/Ann1ShX/XVLh9OAXPidIz7xMvPZFn
QQjwKNMqANzZ4M24DdmICd30w0DwJ5NCJP9NhvY6m4XKfvW5dAEjlvfMy+XKArZmyAdL0JhdSX9e
wtAC9JcmgUfOLP5Fzbz844kSeidF1bV9Ktp6wCVV0nFC8LxMg0CYwlrUIL3wxFhNte3uvXiBPQ3m
qful46LqqCRf28ju/zMA+1hmddiGmf18Bzl88v+w5PtILmerbWqYfKIzUCNcgee+GLyGJ+hGnax3
64i3W7VVL/lbXjo+6j4bdzpEVWJmK0Q2jdf47qw4RT3WjJn5ooxJw7gYu+Wyr2GWpVTHSvQYTVGR
PeaqG5feBbhYnBmxTRkXXmttGUPPk1mqSOICBMMZrpmmV7UQB9TCCCWMjWSRWz8BC+7mWjyQ8K3T
Mi8rEJyK4/3YEquDgQ1h/bLChgut6EbCjjuJaJHVtQ0Ny4yGcz/e8ww66qPjcHxUCNmko45Dv2Tx
F9lo22QCkoMmJWZlqTIAxFB+3TrmR+VjBqq0Tq70H1ZhyUtYy52gxX5X6bwHrUIDyDelk78OknsZ
oQrNV5lExyGzEILyce/uOReDmBnUO4FzdqnOEjRQB48B4Om3804vpT+MSbsUG/3YFKCLYaoA4KtA
dRBRUOZrHCvFBv79tfoUBV9EIxyaUhhIcY/nP41A1BSDYnWEHXaO3n1iRvaImpmVxe4xBxpXvZFg
mHLXxfd9wGXZbv8gw0dawKxZeALTNkp5+/x1WgVIm3u9qS00vL7I5rfo3FzfJVuIqHBRT09j9zQf
eE9SCpDpLju2dA4gcC6ON0ZN5nhI9NH7A7tUGwM8vKi8bhaLDkpXM6d6txuiQHtbvNfD+jt3w/pa
7arlMtNQrVo5mchPtgYkey/phwiwL4owVHSqgGD2EjBUMKh1EtdaIb682RfHqhRbiBTak1MFiN6D
jkOy61b3fRp2TolnZ+YbCwiNyt6olW2CCgyT0WrKrc5QVEuBxCqE311JEg7YEEbwjP0I0+l4zNA/
dQ4w4PlIOE472Cq4W74aT5R1BISDdFPWII5JhHe5HeuDcQ5fyuCnBtcS8f73NMnCRe+vq7qa5nC4
RPvkOyaRfbAfMxqsq0JEcaAvs42E7zIqRs3WU+M/L1KmxfKSBpfiAWQebZFblP/1inM2zUQ+0POM
8rKMWPcVYFb3TQnWYvDp/n+G8cqdRDlG1x5njGPh1dBrkixoVYbBiwXsPZsOkOVdgd6ob/10aSGX
zP7zZr1KeiF5E2Q2SMZm2zOfnrst6RTznEd9MKChx7w3DTQr2VigEnkYeMwFQxO+aqonTgeeGWAl
il21lJjQcIUESZFbV2WL+6604Qe13+XXKOGhuScOKODv9/GtqdCxVkx6wMCM+GwFAEHY3H2XjIf+
DyUEA7aPqkoBqvmtuzBeFPsKAEFO+pxCVWR3M/xJEYbiZm6j7IFzb+PUQs44X631LbxWSuvehBNd
nXV+Poa4sl4WtOUb+I+rUXFM9ad56UOPcHHo2VRbU6WkNYYbHD7wF0iPrF0KGvHcJaqezUtvvHpB
PungnSXFqyMEPAaWkZlNbvF2qsWJrZqmF/SPvNOrtn5hQb+HA1FWD6JsrawzwWtQj8BnxnQ9kU04
xFqinns9IN6YbeT5Cz1Yjclv0KQKc2pjd46LaZv30cv8WyQzMZK0fOmaG6MJSGyKxYqO7LbZkfRm
GsZJBCnX7HQg4aobBVzkvXEF1PEVaTRoLTWs3iyx9rnFZlPwS2Fw8n4ITXcu55jzRrZ9znsRthEK
XuTYMuKpnWclsyrjLbNx+BYlpodHRz5kZ1sLP5xj0nrEQOWvlslUO6PMMCFDlErYe5liz4RYatvm
+2CIbNj7TB3sybJCQqVFINe1FXchakLPG/X3I8noLrQMtmJB+lx3vYrYSGuyhkgdEAybg0h9xZX5
soRga/ckFTLR7y57F/l8I/4sFpvZ6Xc0k/gjzlGCv2EbSY86m+DXwyLrz5RF5qZqAp8E22TClujG
cqwyhwsWIebhpu0aI7nyXpPmhO/TAYsWPHhB+mXw6W9zdS1dX9XgfcPlugOfmvr0To45whg32GCG
O+F1H9Igc1EGQrwW/ap3N2zTzFfaAgcjbCNvY7po9+hhVB2v6QXciMimwwTyGwnm+wCZ7JBL4ZZ3
FfEUOmjd3zaJgAp96dTLAqefB7f3EbBJnkm6qa157SbS4iJmXed1Wu3Zt2lPzzZzVBgZ4EZyIS9J
v03yuwd96TpffyVGUY/Rs4zZbLwi3HbFGo7qOi76bXMWyyDfrNkXXbNjpMvPZNJXNI0z5SQAxTTk
UCFGz25HCAatYC50+BY8RbGD6T7D5vOqHuQxmNJFmT7fVL5BnqX7utDEhu2xZ0Fop47Q8OjOfWC2
NmhUVMaRibZHqiRNxTo98AoZ1aLYv5s66nMB2LgIqOCfaCLXMKAhfLUgTX1d12QyStuOcH2fwrBh
wVKNJy66iZ4/efKLxcAK9uQnZrfvVTyqgzJec/iI3rEYctsyzpgb7dk+jH7tSoF7s9lsclcoinSe
1sL+G92xzsqmeMxD5qq/kys8yqqjDK+RHMUwu/mVTe+M/hLa/FjG00u84JqJgCTgsz79EKP5wP+3
YIEGwQxn8TKqLfi3q8Wtvls6kF3LuQ1d15w7Ebo0rfTTzticLUWU6g1vdzrkawapfZZnnOPAqDoV
JYsX+PQidhNJxEBpQO+3l99kOu4mqqRFcnWehOhi/8LHufNycaoyC4txNFIom/oYSwmteCRmIGlY
sRAXeg/KX9tK/7XInQBvN8i4weuaD0OnsbXaQty0iDs0tHavkjrPBHo7+AUUgE1nqeQlEobzzhRs
PRuHHM2oa8eQupBjhOPgjiZnlqxc65X87ZybqDpVhlkntpnTS5jLHliqfvIjtRcwNaiDqvqHN5+i
Z+hpbArnnu5tW+Ux4MMua4hk853eLVG6w8PE+3IJD9MKsdS8AGuez1DeFRyQH8nuO8DhyFZ9C1lt
H1yZTzgzfuIjT8TPIwh4sPcWFsoQZs49SsDJlQyVQSx/3RyZ107CtnZHHUmDctjn/dYlwknl0AMB
+lDHW99Zahu2ykfwuJJlQFCRC5WEJBQboFUnq9tJMobeQ+rVF6XypK6i7+FzJOC9R/U39F/SQ1AL
FhO7PEuyRKbaLTiG/KRC3SO38w+GSKwtN1VrEM1xBCtbeL0PwFpQodj1L9UQ5xrU5hJcWFPKPN1a
5nSk7rp7lcnbO4GDj4Vrvr94pQ2vTRD7eJ8Dwvp7v44ffwT1is6U5CpryPNSWUciBwo0g1bqyJJC
72dH+TKM5+m2v+cRJurUvN7pzeCyindGGae6y4PnADZOXaL9q/LIir0fKh2k6A9eejgJi9DnPW7N
cskn/3o1jd/PFGN3IJKi1Z4lkO1ey5kD88R7OxUKHYHS2ZZwYd0PALwclGUxi71Lo5VIehStpjIz
gLjOFA3nfNyL2K2eQlxAJDCSocZURg7/sWG4bbKvet+GsoudpvNrC5js/vRZFg6TIES0r86FbPye
3onMbIIu5RmVuXmLvCSg/z6g8AeLu+F2J0F8VJqWNq5CsMvURdC4xwgSP8l1J6r2xIY/U+X9XFBF
tmjIwxfJIaldgvOW3gdE2FdfYW6jqXtjqluGiRvsBYLFOJw2dF5m6DnRyuqn/iLCEooTOiz6lDlb
R99QVDPnVUYXkxRN4rAm7oeRAZbWEyO3oL//wrlkINwrIWFlxy39lr5AYFH9A5MbFivZb8X+JXlV
sja6rjurLnqTLkeBsA9Vybb8J/30AHGS1tgupH0rVFsl7o8epNlyZRf9TaprE9kuPtGkhw55C7CS
a35R6CnWOHKJUWSngPxhlAHXJIhpitE1rl6bNjFdOQtNSJkA5NrFlZbuBgMIglYFqdlKx9mZ+QFF
5KOQ2AVpTLj76cgfjf0l7tgQbiIFrRUlctiADid1IvR49oQ8Cm9Az3ctn/wBW+CFokI5ppc+j/32
NG9dDwTuq0brFWG3Q7p0MGDzQdzKy8GNhwgrBNjEMHf9J4w8xmUkdxA/vkXbgSb8mlzCR+NwTKyg
Hk6lFpW9L3ez+CLH6fGeTGU60cNrotVPdGRKU+/3rjoI7pQ0L/21hyPQ+xorl9IAL6igqK90ODxC
wBz+KC4zpsjbprkM/854iDmbY8HDiDyJLgNi5tL75i/pqbkvZftt072LDRWF33udlYoLZRrSK2Ml
RUuaKjn08Ve2PvSwFY4r0kg1a0zZDnGxnkowue6DoE5jzNo84PrwMKbi9kEkaz2VN3fjnaz/909p
md9Xk7wS4/HHCZiK3MmYyjen5TwBVXX98SXdq5li7dbppwjCx0oxhh/xSuk+h3+XZEAns+p4xUaD
E0TaA9okfcFIIU/F1QjQPjYWIntc8kt4R6wT5YE0AwDW3Z78YWPeAmrCxXf4bqwrU9x40FuM7JpQ
EsoOiyucDDFiE842mYG3M+HO4408eysElTDdycZDoE7vNq3ASYrCnFlYsE/c+LgVJlKV9p7z6WQ1
xBFAvopwZqwnYDuIYM9vkc8DtKfEKx64oeEp8Ll+8XC6EfR9EYm+bBBk/umryy0pszqBWC2J4bq7
NqVIbtE1ms1/U//UT+AgsJmwkveiGKMsV09Bar7WuCXvkA1nQJtAxeZ/I+49c57do/ptv4xqLW4k
e3/WZMQDHgDBTtxRYnAix16rPmn6sG4HKhmTBMJ/O36nKmwVU3vo+a18myVyfyL2e19wSf+qu7w9
s5fBa3H6FccZcIFgr5g4jEWqkqEpmmH2dK0d/hUGOcJNZKLr1kYL919SO5rGjpX4Ii/Qa9NPXjGp
/uCNGF3W82z9cT12/g9sYSj7KbpUInSRlOk3dybmbLxrCj7lOjthC/1raVkvQbtMucRWD0k4mXyH
VSNMEnhPFnz6LbfJE4FWJfZOmTE09PLSifEtSkxO6XcYvowGK2wlcU9frwTRkHy0yQqKxYaarLGH
0+ygPIYqlQm7M+AJQafGGlMRZSyJ8wohpZGgO96UyCsyTlwFekhpTgk7yvGnQdm40UWRq4/pnC6A
JtqmutBKYwdx+r+mBKYzVte2+Hc4Fq/yGroTuPDx6LTyLrqpbiKLl1KGKozu1P9AQnyWDvXQ+esT
RcEkPWTzv4EQSyj1WGF9eU170xktDvEb7RhJwNQ4AscJPOkv0N/9BnpDO4jVEXks1VYIW7CXuTLS
sjXoTWw7G0UVsZTlwlI9UWNSEP7rDPlzNKaOcXpg15YsGxNwPB1mfijYt8pc4TOBNAAvn3lCTE+A
9m7dgVN4Jjl4mLZ7zbdCazpxU7CZBxYMw04FiP49OnVW0KuQm0WQnUXWg7O+/nLpXdUEqRSm12L+
Y6lHEQQK+PESBIgshIdluPs5TIihjeUOvq6r2NiMNS2dcqASTJN3fA+L59lDpFxVpwbAk9BS71CC
dhZ+3XAkQPVlBcYcvZVB7yaW6363s1DqigaNfihs5yN3yO8J+2tY0+z9DiD/zAS2IMHVwUhWOO0b
woJyz7LmFGDXyPt4e9k76RCGCiCM7KkM9+6raFOaqoPiiD1nM5so2+FyJJD0mg9ubrhtNy2iHBMF
lBQgl4VYo4vhjRSEWMBhhXtJeWKUX4wagGmbTBLTRHaURa7UdUSBBHIkmhW8pZ9Rbbwa2a5O98/Z
edE+fIYKZhJVVUOO5b+7orHJSccQJ+Sz5bnnKtNz1Bzz22srOYWTltUSTtZ1CUNFbS2yppk9BZwg
LrxsKVLHkLEOcP17/j/XzfScvtE8BwmSMO4ohTjuDBorjbC6kN0yBXXR94y7xyAY6WnN6HixnEaS
39bU801nUqCJd7m8HaMMNSzuKIw5czFzvXZDe9TCU5zD6OJtbifehBzZk2gIQk3GjfzbU7KssSSL
qKuCa5zV//pGvWdWD7mVGXIsCfB3SAAH4vjaV8ND/ATpx5RGAiW9V5FRBdaAuKiTwjfL6cNE+zPM
UIbAWMFYTphOAXKFCgjNOzUCs4uu17iGPTWi7JPDJsjreYDegQ4jot/Rpjc7Q+PvlC7gMEo9Dtn+
P+ZnHHuKK/9sJm3qbn09bKDjD2bTfdbeRlTRetc400Um6VeZR1io66wlJd3WERwI5nHaWRHaJN1L
BbzkIPRma5kfWiy4Zrk8+3p+yQME6Mg6hcg7xFSReZtM0AuZJLuHVOH3o2YGh4VSVmLsJkEd+dcF
Kx/mUjh3CzBQOgEwkaZqC56pEIA138a7ECt1VdZ/brizK5H9DM+9GrRf+twr9Yxs9SdPSO1L5n7n
zYuW2DN/RWnQTzG5PKdspTVEgHLyxnRP9dGcpVzfpB9qrPJ+z1IUkX2xYFbKQHz2Z0UN02hWv/xq
Qch4aCz+TXWcx2QQFsjnPGteorBJ4PbTTwwhSuMqtlK4gEgdT3oa959xj8xhTBmakh5h/ARXVcEE
1h2sndV43kqmTN7qFPw5LEONWrR/lD8sixaqnMlxsuU3m81+oZ0ZJ5FsxkMxWT1O/XrKAeQq1rXp
SvoIqyvujAGEpMKcXLvcsBD+5ARnAxAVpdnHY+5xH7hyWi9AvTFhX1ybgHTb78SVikNsdJLGowlk
CX+ov/OujCCr3g99/vc4vl+vpbipKw5CFjVulOqJO1T03BFN6A6SWV2YIkvDGZHCOkvBsMRZaqDI
4FhiYA7wpvVcL4RUg9HJr1dTJ2vXefbYk4CeV2jqC1Uvql2nE4UpLrP8HEDXe1rnr9KwWD4rISu/
1d9PbAYZe2gsA0rzWUdvlBgR+nNQcXQGSe/QHGES1gGhQ2DJJexjfgOn737r+7QJjyY7cpLwfGsA
/ELPeCx+wXmPvZufpRF7UNsh+UkZtKpXfci2wZL111VXEuC0pPsLOe/5zHLhhscV3hKdFu8nfnyh
Zw9JGT8ChOVQklxB4tvfLHOevojzCwf+bPgMXy3UXQJgZFM/O6/GqwnDiMHn990XnD1xAtW8/myL
AWlptKUnClKt1GOEY0IQjLdzz1ECY5xrsVKfxkWm4pB7k0NeynuqyTsZFHxgvdf/11YAPTnn9eRE
rCA8Ytcpvva0/7MxhMh2hNcipqgfopFx9BEMXd+7wU9T2duOw5JVWZnZK0EytrMg+XdAtlsft4r2
3EBVXTYSyY+mnqGNcJg8IhuKAB3/+XVu6pvp4QsZ5+OMl+u8PlC2QXbXvGOBK8i5Ao4x2p3CTPhe
ngju1wwbfmV1lHiqFVYhohF9tbLoHYYKaVrrHvOmA1k1hIl5PxJGvARKsPJDUwsqHFkDwtayRn7x
qq5LQ3l+KMuZadnswTIx4A2MlSzbJ8kUdy4v4s7XyVnxKOecDU8wW4Dwrs/ML0b60jXATxXUpI3L
ry4rNi6It52G0m5oQKXwN6SLbWmRz7ZIYEapbvl5KTvK1xuroVWtYTDwQgRS8xy54t+r3VSb66KG
9iOrCZBuEsXpfwPs0bxGCPIT1hw+VpnAqrc/nE56npcYXbXL7BOvJsmsNJZos/seQLAiIyJwqyKx
NU7T5t06P/8triCkFXfTjBI1C6404Y4xKFWt7TosYUwLkwkC69mjBHbWxgFxN+9SKE0RrtjsYShg
RTRKzbGakb1UVEjIX7T8wMnASlTqLCcHY4/Hk1j4O3zTI59J9nNNV7Svi3eU97/KlZW6A8OBfu/T
U8vve/KydnQA4MprB3KppU6F6YwHjBYJVolWqCdmrMsF5cSkaZZKcDu3UhhnGRr+JVVLyHW/X3dY
4lIoPqEMNZ56k6aQ1IZA+1TDjGWmYTwek3Ol8Ah0+XT/dt98S0s7sW6y4YgkJt83z3dzy/FVKU35
uawYmdLIkkxb59C+T4qJPTskdkWT5dWIlQf2MwmzBIiRELsbrhmJJVZsxwfRRZ/dkSYMIEEmrLX0
cRluKGCNQ7xJwEefEpmfTwG2UzfOcAnjGQYp4Q5qlgnHI6vGP51jAcdoSqj5HTCeSoqDS9mTNajw
lchmptKCkpzIbMqpeM2+sBDlRvMaQ1/oaFybEzULM2lEs4gD0Y1bLJpHoSRV0a911YbBa2ebWhcl
hIjXPvGpo0oOpq9mpcRQeyge4HRkWyJJbEETDpzdFqEoSEHrf6Ojl7JwFS7tV6ZRy4nvtwx3yto/
Bj9iGspN6qI3HZub8E0fTT5yhGGDK10p0ZfoIKKTVyH/RrbsxHQfLIsvP21TkP7F0M81E/U+V/PU
+3rlzKtwPYAVzkdt9C3rVqky3evJtZhnylKfb8QjAwOduwTjEWrsq3tgHoNjZl7oucRUHZl3PlUU
05lSZdCG2AV8PY1yHrf716SFolRO4ICF22DGRwttyv+BIl+VInEb48Sr8LjrSWJGw9LrgZ8+kaal
MEvLN7/6t0MflqaZMCSC5ispnDmdfRmqlVAlKS0ZKZJ/L8ab0892WNhbOGd5LoRfu9bmV7F4FdPf
RL0XI/8ZBRuMvU62LE+Ue1TT4Y07EcpfhBDfEHR0hXlo3vfSH4MIZktc7SSWl6NQvDnXeKi9IP6/
VaORNvse0z+kkN4P0DMHhPQc6iXfURDfDnxIkkDO52zeJPoZEsO6QB+AwyPYPtOMfyAO+Mw9nflr
YPwqzc5j7GuPkQlqpTEQ2rcdPxW37kv1cwUC1FttbGWBLAu6sGSRfop/elBOLr0XwLGFNZakCG3N
frpR4CD0AhlMsLgy+EF7N3gxcuxSKgbnxsFFhOBcLd0Z+o8JodhUvnm/FOJ7p3jMmd9qkvyd+X5m
9CLSNlmJEf3qvNDzZPDfDkC507czu7nqhs26yMfyn5CrTQmtG4M4mBn7q6lJt//q7WcvkWB3X3mU
MktbSZViksy2TVY6Sxq4E2Tj9vigWxeFe1HCHVuTqNbfKTdXESTezCwskfgrvBtv6TWBUQ6/SdXV
qUDa8APpf9RZcdybnf3G6S4QB0++jW+sLA6QkdRbEl/RSHHaJA8naxUQl60G0Q9MbVQhi9V8Vv/l
UP3mJv5g89sF6fv6I5IY1JGInHrn62B6mEZ72JNDbnUESMxJAcKuuUQLtNv8M7ZGKid9HX7rXRGl
1f7MGWTxULCcvjBclFY2xyHgTNqnQCXvI9eChYDF/TdFp8WwXn+ENYmhMyRavmpQQ8/8r0MAN2Et
5DE5zkSEBn3YPVhvXazsTujCdVmLu9nPsC7XK8i8DxMLc8bj2Khxl6O2HmJuW/zbFS2gKS+qeZiR
2bMAb4kLXKrT92y5CQvYl9pPyrwWxQUX03haXUXgyIu86bBTXbdVjL0ZwWheQCVAkfMh3m6IimFU
pReTPWeTVbduJvawhYTD7bjnpnV++I3iqwhrw7AWJ6NaZEU0+F1+oqRxlN9XsbhIsksGGITli+68
UfC9qv1+1UqlxeanCle0KUlyE3OPmOcTcH8gDBSwHOytlZ5DuuYr08yoQQ5VHA44aXVK1wlX/OOL
Q6ZjbJ3gBupsS4isFUkZtQwWVoQzayfUcGoOd11CTL6bleaZ0gYueMFEx5ZfoFpjPxZLa38dcpDv
OuJS6dT7aG4xKtCLmMV/MJCHObSPttHj8YIhHjK3Qfoo6vfHGmI21aTi3Yaz/wZU901shxc6h2Zs
01/947sMlxKSQkEx2YbJIeq3oB33MSmgel1FOAN0Iri0RlLPxcYqhDSCUhAJzWQGD9GMuN5p6v5+
K6OMqyzM9f3EsZRo56tc9knWwd1oRsSH9DNwK9TzeylTXd2u2GuVomeKsOewxc1lCUGTjoPh+qlE
soEB38eLcuOp5oEs7Qh7RyqKEXrxpv02faXh1+p3rDMB18eb9MHsxIKNb/xHTXR3cBmA1ngAWaFa
ZsuK/XRbgkBDA3H8QXfxvd55dYx8wfGU+mXM4MwWBGvWmz+Jq2XY5jGghbgrhgj35yxe3Cqe2mwM
Ca0LOGivfeoDf1UxdC5JdHDbzF7OJ1CQGvPeDnTSucY512cNbS5oxclOc3mdXS0TzmQO2Q1OfgvZ
HC/Y/KC4i0VbMzGjcxiuJVfV7rWQd71N4z32s47vFnM5KdZMK6b21+uqo3yWHcoQKH4QQ/hMDCEh
64w+mR1MoNJ1c7FE5XHUIuyMqoSYn6bMgD/OYMC0zy4sthHi2emKcGpBSRYa+sVnMwCWrD2uhc3o
FX/q+FBU0G8qPV1/Fc85pguuvRSCTEoKH+qx6/uXEdw8C3ZRF9nUNGB/BYJ8zC0vDMqr/t+i2tQF
R4CajMrA8tQYUJHGke6Xj0BhX6UWPN1vLZeaiGAMCFUEMRy0ib0qCPk55G6tArHxAQvdJnvFeSsI
DF66wg56l9tw4NLqeWKDTT7q8IglNevkNfFa9P9x/XmxsT4Hd2XXd72dCoOaCQ69B9hZsO3zsq5h
nJfgmNv3ms+y64tfW0sLT6e+s2/zhvCmKEbeKY6mSTJzkOjSPl2pCHJKGDMQvldh/9COets4gPQU
Q5sIsmcOtu1Bj59BgJs+JCb7dkF+zUE9t5NJ8UWQhXtzD8YJ78u4ChLmKbEi0iRbs2TVn/5JW08i
3PsYTHciDczgLsmJggqqtmT9v2ESsP1Kl2UVm3/Q+a9wUakOnbpVua9lvctyjiIjHcyCbBn+Ln7e
XxVQel1g5N+4BIs3XI0qUvOs0gagQXbHZUb7Szd0oOszHoD6KTvHPPioJCazmnkVIPM2ntvHxV+R
B5BZqs4BmDl6uPVreh5oTW1aBiomKOSIuvT2DXbBugI3quaE6lR8rzDfgZXOfFlgBtsF9d6jggBx
U8n6r6C7d9S1Z2tqKspHRDbMQp25TK/lpk1xrpKTK/ndX2ORq+AGutg9loHmhcYOjETjnScV/ASS
/LuDBwKeMY6d4W4C5T4EnnGhxbvSh5m0s9YFTgzVOVUk2OWgnbBIRyUUVqelXGddWXkP92kzO/2F
w/cc1kf+GZQ0h8q4tMzZhfId/1YGit5QmEAxMmlW0n9l7d5RnmpiBO/0qRxVsI+zh1e1yAsXV4ny
EtoMqbLXHSYphwBt5ZL9Vf3DNf6AUNKwEFCKDD1HpuLNbPqa5Vs3sJ90avDqzrax/CXEQGqzN71K
xaqgZAQWrBsC5H0BYEUb6AH9dVhXag+bIxwANXaFcXjJWn7pQMCn6VoSixrqywgjrRqdbvrpno01
DzbLlY/rFc1XkaOrFn6ExhT2Ve5NSoju8ZN/PuXTKjRogDwGOprELHF79BWhHrWNvZE6nGzJNAaV
u2Vt3asJ+MgEfYkmfTyv+UaF7Th6cPoD9Eipir/fTKei4prcz9jAkSBdyuNe8P3PGLKrvYLMiaoa
AwZWRnPpkTVdqPcSphkFwG1DG3CGwCnqO50aPwfE6DXsfCcjQCA/LQmCVzph0yZiJ4OJoisgFCb1
xsPkR8ljY2Eiu1881BMjf6J0MNR/TNi9HhgRu0tYnpFJXR6N+f8t76aOwUZwJg4Lyfr1sG8TE/fp
20D+sVN33oF/YMl+XricyIthyjEuB8hz3e+xIzpoAUzVO2CsRojflTXA3p9m37ae0TAmr9+VDkFb
3OxCT2TfFrCo8sVFetoW0zSEV4Bj2hicjpighg4WWaOtKoHhbj+lODxKfyhGI9+i8uIRg518f8kK
H0l0H3qtbujfwS2sCy4XeRoJoZExsgssS6puguRZsKOkFe9kI9ixqv1a01D4aNz6btqluSIBjnU8
YES/IAtIBTAf0INAn+a72czsEBKleTRjmecWH0eyIucu0W/UWkKBYlrtqNwRw7DCv3JF47GKs6yI
6Hhf2rQB3y55wrRh2ur3esE+xAvmw8gF/SWY1Xd66m8B4YRD8QTrHeo4jsMoSylmEExMPkvlz3o6
KivJUDseZENc7hgDUUXR4y9cvlfR6iemOecc3AsxiamOuz/MLNcyRjwHudXgUbpBhODv2gqmCU6r
uofUfStUwmOG9vGyTCf6pv+PcNWqS3MyVsRJYJnc+Ace/jXuHcPeraVrlG+48JknsMArtTikqr7w
idz2MYFAPWez40XEU9j5F2iW9KZrp4983xbMQETxI7SDz2iu0XV+N0aCy3bhPUEvBvyMmXzJMdha
sGpwCe/I5FvUGi7wJ4Wsl0KVaffQIvgpYRct8I4DfYFB9i6ErAxJ06UGCC8Pv2ADI91YdlyIoK74
ynLFBmilXEtF6Y+RDjaOukK0+3Ip8knwCtwyxXSRoi+cMzbddr8Ex50RKDJDdaZ98GHEX5Cj9GCz
94ojRkF+S8YigGiG9TCcCSdeTAaL/nExGM3r0Mi/Ewk7CWIbZUO6MJ/rvDK6USiyKeNkjqJ9HFVp
MICkbLmsF1rO92+1jujEEKG02sGXS5a7Rqn5vxWb7A84A6RBtAhIXdWHjhHS3Nc37tm6b7ml/Isi
72hdIIwaRe+J10LUI13WyMEFVPNszetrs3hVHOSTqFhLrRS9JXPefSUbqOxr5RKKF6PLj1dw48EK
yccIXF3loLwLO4fKkR7XmHpOlV0ytpl3MkDI7JqDBj/dj5wZuE5JLMLw6ltJjps9qmpjsBSwJQT2
j42cLTiMdiLAxvlyRLhRVqmhRyaiGcyEHT7hjEr/B4+LHaQ1fVsPxGcUK7mX7hr36RHRtK7w1Nwn
r7PLZad1VsjZyfRayyBLHhvDxFG26CcKd2DP348Ac/J0wjg+zqy26nTypbta3cv3fsSWbecA953F
5DZDGL9wu7RjMLm7CCMftOi+QvyQwwdbTf3Knfnq4B4xMCQcwhPXlFSmi6B0u/ha1q8TXacw7Kh9
2UlXJqQdG2FRIER0sUdsEscxQ+zhsZIsfJOrpdyIlHQ032ZXJYQv/P84eW5V9eGiLdKOsvrpNTHL
XChBy11SAGtIhqC9ViXISdeLLHkQKZG5MahTjO+hNLMfItzsgRh9HI1Es4z15nyThK5wkZYKAnC5
EPYfHwUxO3Np75e6udu7YUu0faoO26x99Oxy9ogb1u1S478oOQbnbAEFxl5n1B7gGcSY5XKtbio6
LycMj53jm/gtly2DaqibYeOuSpwZxIPD+sRH84Pp71ba+3L159uBZ6hSwRop/ndf1PK/ePDDR3P5
AM0bwtILvQxnwi56hh62lEdoa06gbr8mzHZocfl9DnoNuwYSgoahKIeqKD63ZMRZV+s0m+FGmxnf
cbhqZz4tTojuhHeWYoshsPs5hx8MpW+UoU3med3V9B6Ic9yTApugkoVtKfgidP5nL3SAq/LGndua
O2QO2u35q+hlPiSH9UJ4wpu7QYj3YZtZUgsFhCkjEC7IFbIowopwyovqRG+zyq7Xd1nbFGHGNI80
FXL60WbA+gvAYbQYsAIUhcCZHljhSLFeQd6uIFDdimpwcMrcR40JHhOxMI8Eaf7ssbrxVkLQr5ho
rmCOLq0pk8T4G135mxZq90BdD8RYezn1yWvy5NzJ3b+EVr0kwyeLuzH+CN7xge5paCzmrif1drBm
VJi7CQJHZGpZk6Flqoh+4tG//+uMcundUJ9Ly1nD/ujTLWwjANmomoq0XFjW6/gXdqtoY8i2S9pD
T19IESl0L84inVwMWatnkyYZ+uQR7dmABoeJB63ee/Q3XFebwZ/8sJ5MtdMHByAnB7KsbVy6Mnmp
MtP2CFIQRzFNVpHmYgC/8NdAIW4J92ngxBktSh4Vkk2D/hS5wNbJEzMqmi/jdgutg3wg1tr5dkuy
4ClUHo41VnUfkEZK6NaKnXoX1KlkAvEWJvg54zyH9zWpMVcSrgTniiHE/YJu4M6VNx1Q4Jgdo4Wo
qD79gr42iUbAnLdHxIY4Igmi+OOUEYCmmNa2ZZn5ebT9eEjOGuL6WNKKbgv69tUKagEw+QZt6vBm
Hm/KMkDpw0V869tXv1d0cU93kg9k2KuwF5nZH9RqAGNB4ZvHTso2bkuKxfevgw0T4rgVlUqywhNl
KMORFACKb/gJVXEQSOGIjz/l56qK02/9sM8f3xRKxp+PWRfa/OMYY/weUs8CT0E1+eVoWGKP0Czr
RiJDgDlJlBiumtY0BS9nZiInghVS1tuoUqeYDPMlFXLKeO/OzEcr9aJLynOruZhcxqI6WSqeI88W
b3dSACsdd9eWVilIwLjrr7EtXA1/pe84Y4q2+H5UVs00r8zxgdCvTJ2aQbO1dqMMIHyGya/ZMDKF
lZOV3KrKfKFt/u8GMQepT7/nIJptqZWS6HYBGhcsRThMOE6hs1q5SWZ7ORSEk48xApwG//Gqf2UN
naSLzHMKql67Mpr5ZjHHe8qLULwDbMFseVdgUrlWpmz0i7CjEv71mJvqQdvXf1ermv+VLZkyUeyE
LGeS78VOchOay1QaCK1LEYjQTgieNxTUOOEjS756/2u4B9C2HB02u1WeX0r8OO8SAd/gQC59UGTw
7N3nsN56J7ClsmR9/6KNH0TejYDSjLDL9Hs4XExHdHqNCH8o3XA84v/IDBjDyTI+4Ma3Wp+bE+3u
HKEVs+8kCPQiGYpKxvl4AeDawHRAP6ZZY6We8siPc+Y/yuaZxJrhYkcxWxM25WoNf3y8wTyCp3ZY
4jl3mXYfQ0NMcjFGV5YIyT8P86Xs2j2x+xOQl+OXNvxCmGcnfzC+O0HNck8up47IDwfd+53RwFbs
0sYuG39Pud5ZB03kLnzMIxTO1ba6/AhF/8maTZJrjpQXGRwE0YaDjQazhamikRHg3kZuN5bWUI+h
HFnPDdx6IaGjEEPHH9g6kE/WDx15Yugq4Pj1dmXYpas0eweKzEkTgqtGd/zcbDgtO2LqSi1NRW4z
4oFnluv1Y5GssAW6nDm2bYzjkMKx5tuyK1QjPtyaX+JNeuDSAOWkAsLoFjrQflioVZ9WX6YJ3kXn
APQzkxvlc4ewReNO3qCi9lN/74LPRCMmFXsY8d/R35118NzD2PqEkZYHvvmgk6/TX3yVk8TgGasK
ZiTmtasysBzxTecAsc+xlQXNQ93S8bqzv9pu337ZgYm6j/G067OTWyrQ/8GAXEk5ThxuC9wczZpz
/E6HJ9CGfhSsUYl2v/Ah32352VUssxELzdrcszH+VeOymaNT2cMP6syZAS071AYRGqvXqXAnM1uA
eLjs4Y/c0OBdggIlfS+1GjCqW+MFUj+c1XBqpKG/0VKLCQQedYZniD8DS4ZR6A9M+b0J4VDJvIHG
GF4uBQn3AacJd/SptlNdv0HPRYCbAT/z/PCT/0MdPABAt7dRuMnd9n+WDFQjMheNdBueK/d3pyiM
/JKiG5M0ottoWOi7jm16JaW9AcegvJAF0p9oNH63Hda4hAC0DboSLfjh958RN2mL89lo6rWf/qph
3MteGgGFfzsBzHwihQZHC5eJqxqwCFEVdfOCWVrMcoDV9etBx2bIuoZ6Cmr4MS8aWMJPQCHplT+W
6YY6oz/ZlY+TOmV0IQL/PaQYMj0i+7uNelJL8jEiLVikFLluvSEZHpCHhpp8Twj3jCfHr+WiaXhf
Guycl9kj1xrzw6akh2e+7FhDHd2sR7vR50jHCfpkot0tbERAVmuB6ZcvrWy4l/Rgh4VlHZl5JhFo
EDUzUO08cTLn0d3jUl2B5zqwo5gBaT82B0BRTpOmx7YlF5DrNB7kpHJ1rF/n85B6mT+C0o3JMGTU
p9PA1V9QAWyQlo095FW0uXkIJPxoPCYRD79BqfKqh9OWvOIdGhVH4Upv1sHzuBGjxXAqaj5REPDa
SC8mq0fRCTYLm6DdQjSWZphm8uPAhjrJz5GkKVPWC0K9T9+rlZQ/Yr0qKkrACep4hTXxUmHED1Vq
t76AHUIXqleIXa4CIGqQ5J0gA2uRFmE5svefozUspVd0RT22B7rNjZbje2RiH+Iwihk5gCKWaNiA
Axc3WfWFu+eXZVoRw+Tk5h2TA2qV+Y8FoDlnDdeIfckqsbWrymwVDyJOd9oYToKdnuBKhGTN8Zzy
38uVh+syXA03D3OtN2TgX83tOS/9q4PTm3VulYHlS3l1nzryoSURxmPp6ZVpHwBvYIamMaRdCUQT
VzHVhlu/mlM/J5poSdt18SJYkbL1DA6Kd7Drl8ALprUcWW5ePWGi394JcCildKZuBxtTvOcPOsgk
PBBrIUzLlD2lbj1kp3oRxDHI3Q69bJ2166rOFv0SeL98DCqXfD+5mol8f11vAJUNrw4w/080Unhl
FamrTlWIREOIk7PTQX8jyWoNAm39yo1NuucLIl9dPn2dRU/ltkeop+w6NBfhxlDKOTbTPyuIRxmx
dDnJPYB08hNfS7AXQvQzSxWdtPGioXE1mANcgR+Yj+oNEhcUXr6ug2rbHzVb702bRR7GeNWkCIQt
RyXUAMTZYvoF1Qwm7QLiAy9xAF6GcmVPEE2jpoP3rcuos1n5pVG6O3ZUjcBgCfSlfMLeMhQ0PyHd
2/qGpqtg4kGDV1Ptz94d6+Qt3NhSnt76ieTtLAM7yKnZZ5UwSppbj/JjMS9qD+eb569PVImiDmWX
8OTAbS+0uHqLrTO96hzDdcsidjPOArP3VDH7D8L3jiaEwFQATml4h+1Ifrq/qUz6WVTMidtJZGLX
+49292tNzaJlbzEsWlBVjIeb1Y28ODaqKsF14fwPTxy5XiyAA8tDyL2rVoHcTizfTywPBiecpdOD
IylU9UvEdcTiozJCV4AxXr4BGPBOINXxTYNWW/G6vfG6DoNUJkKaGtUpQGYSgHwGr3ONmeHYfDz7
REe278snBlOf5PJZLXCd2SB9UGUwXuSfbkZqeqPtPSzWusYo+8AlOEIhSAWOK5RYbpF+fYZS79jC
nm5qBI3GpNTqtd+8urbvxxdTuBC3H7/3TcajXQLPIf0qRLGzh5/7eOn703FtRrdektSIwq97qgZ5
aOTUWk/3+pgy9NgPjKxFW3/dMvxGG5A/TXAl/3g8UPayqfxpvFHoC+h1V44mFPccq1uYmWQlEZlI
+RAaKOm3MtfYhd//ravFH6jS8pmBs+Jhs7wbLFFnLF7btLUOEhffWcjiEvY7djsRgcoKkSIZzR4/
gxRkGBswZLgiBH6BY4tuCI/0+xzt3T2hCc34XgiNfvfIdqiPk+41qQsM4V8utxYwexxN4xd0zBE0
12bwQZTMDhZ8y+NoNNOqDsdv/WXPJBWXh0arvgfiQ62I2/eCovgpKtokoFzKOtQopXiUbO4hfHGF
sm6Ax78ot7d7KfCwKOPnU5FrjnKy1jLrhFiGuFzOrgP6PP72WabSG22ZePkFvMx7CGKYLnVzSYad
NSR3+p6VCmTxfXLoqg2qTF7cAQhRvqy8QbTVUEkRZVGJ66L+cD9W/veXjsMhIB8Q10u2s9dy/9ut
3GXV0NuRzMybAx2OotCp8P+QE40VatfpqHWOt5XNJRLB3Y4AIlEevaP9T/JSpfjUsnDWp24YHyEJ
VfKgPaPwsSl8qQQZdZ5O1dPjzZlGBaZAHitLuPDpcIzzZ4r/Sc/oPdydUnKdCWT/s4BZXOgEMZPk
DfP0VkP7TSScqLYsOR1mAM3m0XLhtcuR0MqYi0xryhnOgo2I1CYOym6oFCIkq21P3dZSWRQ5nDGR
H1/9yL8Sft7VBd8wHa0i+1IsWEIcLaoi8ZG6rORLQ4iAVY2pEzQy/MZ5FGppcR8dqf9nCl5zNCtY
53572vmFThx1zl3mPeMA19p9Jm4vNvjUMCJifMMGLyC2CGCmfI/Gtcz3mzlHl3iUuIqpiKbIywij
RBn2bIAVO9EplcfvEfG63Ngtv8ve251kVZqS4AWgUuJuHNwy7sqP/guq2punhZgp64OAz1lBN/vU
Ju7TV+IBRCzxCUnUoTXyXDNVxj57iTHVW8brwRnduWa16DEMjSW6+Rti6ZdeYJPusB+wKgixEvoF
bR8y52F5sSsyhlkKZmwdISn66s1Hy+Y6+UFjs63RTUdBpt/kbiJlEMsCFYjcFKeORbmxBikyTgZf
loDXnfcLM9AyE4vB8+F9AsFqVDGkmwrXH5QfNZUiqhDwLbIEV1N8jRWzEkTU+aGf4J/BOK7Begm0
zNP6tNm3F3jh4/3S4+ECycZtvCOZf1oYKrSkIMUsVls2z9Im5lAsAJC38A/bRmlyfjQ+mHfBj9IP
d/KAqwa/kknmuaTE3Oz+Jcj2o7BXwXtiLAz5JPjW5DRn1kzd2+2J228zfOBDEeiAgsIyvs4rBNb/
0f5iLZN4Wp296iTxfK7Z4JuHLvYBBWShIWuF9orTKPldU709SJorh7PKG+krOwulMVcEqZ2waYZi
/4kc0jwA7SrAzdWtr4UifPveS0gUXeMarl9ATja+PE251vxKAe7H+w0BejeGDopJfmGw+ebHDedJ
6jFHj2l8H3zkRkiHXv5f/fOrKUwsJdreJuSRiThY8WbZoiaXrSP/N0qkze/Lf/EmPEUvUHWL+qoQ
pXI2NOBpg393wTUTRve4frzfgBH8QSybPtUY2qUHa0enWORREpgjcFstVI6ZbCcjFNHaM3kR4ZUm
6CgcvRijkqgI/0uWc55dmJkCe4Y8oVeKyu2O8bQ3/Vjz5A8zmksV1Gjy0CQDSiHS37upMFVWf0GU
/Ccwk6NaQ/7txgANeIifoKlPUu5ioUMZEaKlJGDHyr+B/Fpbx6wp/xPODcOfGzx0Wy2MRb97uCku
JZSHX9Apxs9kQQ9Zw1NVbPQ4iHjmBltMKObrdhCO+feMntbxnJoY0G1tMcjnnxCC5URlZ6t+H4PM
lewVS43KRXH9rzw/whLNuuvBGltnnnw7NKV/ZZVZRU50wk7JcYu54XSObsIP/uv09QrqaC5GPpnO
Qg/uCt/o786mUQY8IH5WMRDPWUvW8nTfA48X4mA5ZlUpINT+8/Yg7+4ZgxZN90IuVrT8677dJ2+4
5lt66YzsMUeRbzEiczt6cHIlWFskAH5G61ZrgaQN1byPf11NECjd7VSoru1saxFfq0ZDjRSsHMNP
12UCSJ579zN6YHXTUM6nVJFwMFHsUhppTL9KMxDXNU6q7V0QcUYMGwYt+qd5CjcyOs7zY93L7jdv
jIeTTC1o4yRK9QdWluU5zyM7CoazcxMRnH0q8CrNwjReJb7jgSI21nN30E9BpnlvKrdcQ1Rwi36r
wxjsut//I+KAHlv5po7c172inyG+qv+Ut+vvrORxaaeC+FRybrPYVjus3OPedPjkU6hiFX8UNZVr
UdGOcqeF0y9/Cv6r1eq1w3eBFAmZLeoFn4fkyHbW28XCSjuLu9ADDY9z9zqWIgMA5yqoLxbi1pBt
TjXEyZOs2QRf4XQFVn5jeqqY2JNtPnIqnpXT/JVJ8rUY5UuaEF7cB/k7zsFjTUz0msXm/HdkgPnC
GGJ0mRcBjnBvWnjPV15pyNeaIK7GEVnNhOuT4V9z1XRt6MXkczpW4hfYS/jvqm2XQA5CZ6o1bLem
lBxfho9TSwG3mL1mptpmhoZZf4zUqDoUGeHfTydOZADEDzkN2ld/WpAcoXxnft55KLjzIt1laeJE
Y1xkURJwl/AmRWzIVU6UQxXULIUUV9LeE6AJAB/bmzsaj4fp3nQuyUQ+6kbvnUwh6xEvoz+t24Ou
d5DMzGtxltzs0Q6wmdTVBlLKqCP5eVJ6fEjG7lEQpDVoP3hAQ1Ld9C1rpptwP9YNMlB/DnGAf1eH
qHzkkjkMPZhbO5o07aSfPmBKb4t0rnMOYKpsLP+8qbwfxnR8p+uLWknc0AyNQvfPdp4MJNwxpkw4
33yj+mTc7Klw5PsHs8hA1CO0Ba/wW1JkY6F0gPps7cNnRNUw1arPVUFvdpoUoWmsviS4mCbx3zOx
DeXoK9FXqGKZKTlwVT2olN1pGkYmW47TQmaCaqF/5zSv8wQ9IHK8QtgEXys2EL+I88htJHlZ1sQX
yU7X6W72+IuJN2tZtTzLRaK242tcThFGhi/8u53eLnR6pDnlTLpQEL+C6YeDQMf4jAHI+HUEgBuM
aIvEBBC+TOy05qjrToJ/JdJMH1t+HfKpc2ZNA2HmwowA0Dk1vkSbVwfDeAJpPGc1O31Gzir59Np4
A7AY3E0+FDBJMSUN3s/ICAQEkqnHNtiA7iFPD4jZtz6guzva0VHFUh9eWk81pCJyUdJY8WBLersf
afnLbhkV+4STrnqxFN2DoRG/MYD+gnZwD7/CCgB2vhF9dm8ButPUYsyqNuO6Jqmj7ugeW8IpQXSD
jqPlHqtfOPzcx2+MtoPFuE2+vGVYjkPiQKrYxT9Bw/Xh3DM9gKUt/Wmc0Vdg0wQUr0mvJm7cFjRL
wk5kCYdr6GZuITDzFMPJDZjLge+KlGjfqMLMmXSknYqY14xMnyIrnATslf/h7i05+k7pja7E5RfE
thA7QZNNcOeiXut7kK2k46zfAY2S7NvBrxawpQH0/uINF5UDT14nHbBkxbI9B2/FA2Acv0B8/zQP
n9cq+z1WaLQpsbDMmU4K19CLNPw3xfQXWR0cqiSR2L5Q5tDaj/skPjc6gfyKibYgKmGqQ07/ohQU
YqWnFsw26MJ75RRHQ4krlG4izYA93qxH7T0mdjCWyn8Fv6NdAn5eYuTHmE7Rd/YV39hWYlHnqAwQ
eQQZkT9WjhBwbASKx6W9ZeXRJ5qQJz7Qu7kA54xP7LxQvE6rg8IQBHayQOfkg//K7qYQzBlnJVW+
T4Jo16tZmnn+Dh8ezoRYnnqb0DQIf73vKx7t2x+ZbzI/i7nlU5vkrhAH0OPij0qoZeKa7OITqjcV
jO7mFIqQ8Q1iKNmTVxivAJBxKHL/78NYgNpv2P2Mtlc4XI3KiiLKM10i9K9OwgPS1D+4s78toPvL
gScYh5q4XYqei0x7gipBKMM51hVRaHJInIrQgNdECSiRi21vvPJnjPZ8N9rZSbexEfg2METwvmB4
OhQ77Y9I4lkaStSXCMsJoVMy4ec+PYd3J6bVMBWmFTDZ1Mjhtr0C+NrfbviN7w1NJnID4kROMdkX
85c1cx9TH3alMzUucseLyAj3oszg9B7MBO6/NIQnvz7mzZDvTpfejJ+a8mfI6410xDZOpcIjYXTx
SH9Yi1gBiLL8REu16d6CXyw04TefAVdKsUctHNsZ8iwoj+fBK4rKPHrvmblPMz7XNYw8pxG/Ecj4
EqWXiUjKDzk66S09VJxfQV8qStcIBgqJSu5eqp+w2CYs2eWXsc/Rak5fim69JbVRL6fnqd8/ihjK
CGyzF7EC+/tnGnRk6IAjqSQKzeBTdW4lIY8vPWhiL5OxYJogRnq4LrhpJM/HCU1TT/POBP+wts5A
I2VPHhGuAvXbU1huzbBS/M6MtONXZxZurSjMtcrdE34au9f/GOV7RcS6wG52ii990ybN7xVrW05H
pDzbM1TqDwbV10Q4V3hX817dZw9qGX0RYKPxLfa1zKQAxA8y1TOu4KarBGENXNL9dm0zo4myT61L
Vz+wSeurA6vNwPTN3c20kK+530ZAk7o74EvMK4GHZ5mXlFV/tVSOkbDya45rJqrbqu862i3vqvxn
04zWnsgTfLpMEa6qkQfEsqhoVNfsqhhHPs+U5Q7KTVHLRHGjRL9EzX+nLSFssGa79/Os7U9kEZ/m
QyvXunGI7uu9myEDWaMVujU8L3CjRZhZ/p+dRxxwZybaSBQXHdZTw8j/Tzn3vGqm+1OFHZ8uTVrL
Jm6f4vs+OGxhq9S2Jl5vryTTlpYa/cMlXiEc/yPLzk8Y0FsfI3F5nlJ/86hWHyLBIUaq+rlsqTKs
lj/5CsbtDG6kI0IzULVz26e+9E6BU26YoM6xlLBgjvtDkviS/2IZ1TSlbKK7HvuCWQ1x/hIKPnIM
qk5702eKsIh4w8Zh4NujLDdTtzm/mU8BkdPXm96Gacf6ydjyXEbiioKp6wA8zbZAxJlc3bkfV/Ba
DX8fLQHFElYdNObE9Iw4bwTpwKdMyqbGsVzCA69kVg192jWsMkY4uZgNC90ozpyjquLwawlLgpDs
/elKF0tmCvR13wh4D4IG+oi3ZnFms3eagNJDoQH1WGR2jr+uTVWNgOZInuXJm/VIMm8aIabvUoeB
h7SgtnBVTSKfNUmZU7v+46iceFI8mmMEKwKYoxeaZ9fSsTOGVmjxoR6tVX9Ycmj3J3a2xKuzb6QU
f4Dzqq6EfYOzce1Y8nPRWRUBszQB9xpiY0Iu6GNszDRQMbo+jRf9jW9e/sKrgGYNv+2DTQttbUDb
YebLo7WWHVBww/4QRkpSqiuBywy411rtn9jbaZFksl03Ha3S00LwNevHxrM4nxopjgvj+S+uQJBu
PyYRYv8XnlDp1ZNQToYta0KQ3RtX6EIx/LB2UNu2rBNYYjQ6mBGVp+CMzqQx9LjbKWaJ+T441r3c
uRTHFpKMBQIKk+0Wn5EcBzXcGERE/TGT61WCTuheOw45eWMtSlt1zLo1eijdGoNfm3T1HI97oPLi
WSF9G8dI1r4y4iICfILAq1deR2BKlJgluSzVaLTMO/kuxLMmbG0T5B4ZpxvvHtIBJFwADKV6tTOc
0w2k+0d4ak4F3V2ztmY+A48IVVpw3JFxSbEv2iZHSalned/UClDcVh2/jPGdQ11GlUGjHqyJfj17
QG+xygl1EZ2rkWLSlVXIajTm5glXKCeezYsvlnzxo6bKquWEk3QWIoSX97N82GBYf9BxaZXZnf3l
cfGiFCr37+Ey5b+V6zHq0wW+wVy4wrsS+9KnRovEKRsES1NYcTrtWE9d9PqdX9As1QlcClFZqXyO
smZis2+J/b77SagkMjtJIlou96Fa/a16bYH9j267V9nF4Jsa1GDW/N0GHUcdMTlzGmda3QJ350WZ
Hk2HgJ2xsp3Ojbf5n0e2gKjvYdrl7qxvMgK23robfYA+70we+VdD0sDLXAXPDevh7fLy211jTj8J
uVBeki5yGyUHU7MQv6eGpjRf/oxjag7s7aM8CCEQvF9WaSm7Re8YuaQ4hGTd+NW1u4sVf3vY6rvy
fkHxRad9RRP/1ojJLCLXhHVcWi+4Qq4B6GQHaJccKGMJjAw9TGr45HpGKw0HFU9xZfezFQxIeAyg
6hZJcotOqAkQs826PNzVhNZyW7rlWwJ5rIRReihXiugNyE7ws8ETsKupAQo8xxdg3iPhOzTVoiMa
xRurelc910f60x+yJ7yEL+oe3wVqB6TGcAT1PtVju0X6qdii41Fr32qBLJtkyRRQLY3AHqmjuctQ
n+J6E3CDfSVf35ZQtHYk495Hq5y9hiXvSCwMUw6AYuMLLVZWzm4Pccx9PXYaaBIpMtgPw4O2tpiJ
GEyghDrz6cjl0r3uvusPA3b7l5m5fwioVynoyFU/DP9MqzzIvd36eDyeCj0SdU6ZYB91fZ3Y64lo
lEvHGEHItBc7yXFjxZ5ge8OuxB8IA7TOqYCGJb6LLcLmcowDMJbglCwLU1f5G6fMpZrsb7ghNTJL
WzCY/0+shmvJz7M67Vzh3LlTKbgz5/nFbzH/9e4P0b2pYLlfKQmM8RxSXRYt6qt/pQDAH/Nfnmlb
ImrwKaegHWgV/hX0tmm3UfHf6Q/+U6v2PFGJjKEd60h6DWZSC6JMwYwA33xCkCM/0yQ6nrT/Pa5N
Q2xm9oDHCPTeuqzJbZjrmYXqfWpnz0GthEDMspbvIHFcX6G+Gs7CCTr4pIPtw8+dJy7qUgz/zwco
ogHRSEbbx/ztTpWlypTMJyYopU34p+bXly58v04PW1NrkOVhyv3/VM2OAGVRnBNxmZebZc84f6BG
kFLjMKO0becC0NJ/CqqujHcq6AyDZsPXQSSQtjD6OXqvaPWmzOCLsu8egYKDCg3CN5IUiYPcGACL
V03Lpn1QM5AmpwzLR8fvTseqfEeS+53pIfeUCoYF3rJIb08ydtoyVc+ix/N3VDccCD6MGZGq9zHl
coRWl1ZQSDzqdVZ4l4UvhBe8TPsmc7pTzUTPiCP4rT/Emqpql5AjFD3eKIf+77g41WSiUO3SFEmD
mNIeVVUZr0NX5M5PjhsfDZkMfT9V8F6aTUiZ3VIHsMnNAlpT++U+xUQiDWswHpSY4Gxy1iOBYZOj
P365kbdG5XqHH8yUscdKlrK4VvoXMgpXfvMlH/ymxi/qOtcSrwQq3TODOny+P1azoqWOGLg6jx7R
B8JhRezRlfnIB0jgqFkWxyXqvoNYnfxYKp0xzJtZo/aZFV56B/xwByO/O1rdfRYNqZGu4lyQEJzN
vXNR6yNP5TrAd6eBlcSIHOo56WYR2wN60p2UbqxSNBWyCf7vcEAM1TP9WBh1sMGBj1Kj+jsrLtV5
sEyypd4ttrxV/hs/w5ROJFZLDGdah37g+dsSirPqzIde/Bh6c7hdr/OJb78rDqmjb+tgJHrmOY6A
TKDokakXNWrVht7K8l0Q5XTvbwJFp09heM/RMrQQQ9JqYaNbRrwzo8cCkANoXjISgjxdvG0Ni/KU
FGRPyos8gyZf/S3OX2xRjrWH1OAQ3Fpb8eDQ8Ib1QzO1EvqnrGY2J3YY10lhvZVWNdm8UG52tUw3
mUIlcK+MEP1/8jEqy9eUmrMZen/nukQp9TjFH4iU21WsspfP/bo2xUNO1Qcheon3LA0noDBQshru
AQJM1FNsQ2ZstroWNaR6FHbj7wOd+bNnT/uUzxDP78JExhGcAejFj+wQmwn2dl+3Wlv6wvR3t000
JUPq5YwsW7WanY0EKbweFKlloUiTMYdpLx9UdyMI9dWmQw9TQ8axqGgeeAsubaOMRySN234Phi4V
x+fQ8JUuJnkqgwU8wHB3BXaqTkydytikp4LexfefHpMivO9TnSys6mfpbY1OsJERtNRPpQd5hy5L
muqB3Kq678BcouexLdVGf3poOigxy+CgbKJtvXP0kwP2BYrUpivsRneIl3h45YfZFpr7DRB3xVXn
XRfTl9sVVbi/QN3pAc492cycSNInhBA2+QBprrlrnPclv40Vb/V+zgqRLoWqQA8o9VRiYwelnXOu
epXKDC8kRrYWC6y8Pb8933pD3I6psQYYT1giIFlgeL3ChxINJ+npmEl2g8h9nvlKq0924m+ZObs2
7mNoLglsLAkL/hQN+BpUxy6qD32X7zmqC/J3ZvgtOQ5bPbITtptqTMpxIqBFfRs2SSEWTQ3xwZQR
4q4t99olqSiIJs+zrfIIkV/keBUdiH8uMKykLDZ6z/uhzdNueR44bybNgFMPbC39wTfRHe/LJlQ4
OyEQInCNAyqPeJp7ioQ+ra1/pepCXODIPNqWtVLDlHLPKcQVGhAw6J3szHoPlYZnu2du+0lzy5Zh
UCJ+RWuKYWumb62RVl2jNeC2MhuRZ5C7NrRNbk/BCRCmSD6wKkqmD17CQ3xrmIZhSu2m+Tf+inZ2
vDqdmEGeSytc06uVX4SxP74fxgwSEbofJBg7KAx32AI5K16EIsIaWbRLH9poEnKMT9OO12mwO70b
q88MJN6k/HJGc7jmSGp3f8TB8vTyY7mii57lWs4IvdzxaBNmvJ6LwO1OEKZCEwpiOREYT7W2KNR5
E/GbVhde2BU/l/jcHLpD88rzFKiSD9/Qi2nG8Wv8l7gqE38eMHge3LvNnsF3Bud/PohOKUu+k0uj
2H99iK6qX8GaQ0DVYKU7f3CijmQj8SqF52kMK6S9l2jSA9J7g5GFrXb7A5B57kaXEcD0VZi9Q9E7
km8DD9mHYPcQaxGB2HJA4cuTO2E32KQi3LJvPUMs6MEHkluVurCu7bC98TC/n4V+dZJyYAJj4TgZ
D5ojwopCUs7viQ3OzXpcmweXWzE4i97E1xb4kFB7h31kPL5lMK6Bzzfbr8sV4JSqdwK+QlWDwpb8
dJwbUhXEa+os8mfWAY2N5tEq7/cJMQ70oXl3VZCK2us44LnsURUWZMMw3+tm6qedbkX5aONq4dA6
NA1AoHD64CIW3j4D57a79fVlZ0t82gqRAyihy4ihocxfZJJyo1qEfOoP3JxscZJPEppoWCa42zd/
ZId19ErtfEnV5dgLUhYHstQuGMYWtZcVGpi/4ehPdR97dT1zGBS+0hnBwZe/FnIT02ddL/LHzzkg
rJfN7mgxKVrSXJs4EETa3vJCNLbL9Dkj1llQ4ntz3P+qomgHELh7nM1BUkv4GrYTpYw057HmQr2R
eQSVU0V4SJEHsbfqufd92NsQocX4qA7JZgQBEgJFrz2DBRFarJvpT2oTA6WGYBUgLycpc+S4Najx
W/1fw8k75CUC/Ker0knZnMQKuaK5oUoj+OjShSXL9Sa7y5EJIUW9k8xoMPhkv3D+X3cL1HQzrkD/
xxW26WueBwD+cAMxZke8cPtprvRjSRQ4n/vNeBCJDNveJSVkvogh6vjMWvxdYaQRg2TmweNMZNZ2
Hw7lSjuCw/QtuTYwvM7cCSpo583fjPoFRRY5SQiT5lRuPr15PzUpi7y45ypKEhRPPn/GaXOEdICe
i+7EKRapjp6EZ2wB8NEeD7vOlmdGzSAJoO8PMDRPic2oMAl6NYCgiQRJ5YsNfgS4NRv+zbORf31B
nSnD1tarn14DrDoWa8rnc2Lgsk3q6Ymik0b3LOuOP9MgYlM2UODXFFXA/JeDJtE7XQf/P5iy5rka
5lv85QeSyxI+ZvwAWq2S3QAo93O9grNML4eY3HcJWR0UBBaq/Oie9JWGWR06XQetNtHOIfUbAHbv
T5/TmBbqI85KIN+bfMFb89rprQ2Jn8Q8Zets75eJs1jbkfl7LGOJPjLB+PlZ84WIFl1XEE2avvwi
vvH4BYd28jQrlfJ/xO1bGh84GQItKn+VA84OYt0f8tkVRctBuxH9WZzUNVDAFIGc9yuLR3fKnQkk
iS2rtldGaCtJt2/Gz4WKtlNBSl41Ly8pK2IqyvvyN+iZEIC1oa3agtCwxfvBXGT0QaFnWmV4Kr41
IxeM5oNSkT/RCBXomlKoJxy6vI3tlF6z1gWB2rd7dVl42ZRVzhxdglG3aZqkK0vuS1EV1fijDbVB
ZDKiUitoGiTJlUDfLviq5Mn8JSg4hZKALyokoIewgyXAqV8COXl00FdJhgOlNDQ2p0faZV8ZrjVF
pE1aBbPGZBVDonrvP1egXUStpMexb8GYeBmoZpLxCjO7tHJ3TAxvd3IIsjFqY4QPtVX5C1/lcw06
0ALA6TypJSLfhcLW7ieNonoGBb4XsWB1V1lb4ek1onZa7lUUa/SGmwWJ9NoS/+BjlfmV6GNSBnBX
9+wpPCV92UmwU8Ug4nZquT4rMSsumuMUo9J2huyi0azRUX7BBBGOhkGCK/w558M7QnRLcqc8eI6/
kMSXIYZ7phtcH/HzTjvpADC1SsUyT05Kf9p1K7V/h+caN2Q+VCk9F0384ecU7QR8Zqc5rxSTkAco
YulVeeu1ovIyTbu3JiMydR0RlMcOHz7ReIVSzTT8AGN2mOMzdXpZdRTPS0gUMhbGZxKq8xhRHLyB
cIK+vxvn6It/OC0JHCda47Kz3PCGANtfuidpel1l5iKj22jVk6fVyymbIOzosyVjZLlwBro67PHg
wjCnOeSDOqKW+Zn4uOLS6ozSKFyfTpJr6WWWm9E9oUHzrlL6y5YtY/RzdSDLptvK2zz91CGZa8HI
rbJoKYRJeUJvqGC8d/UsJ/Xor3yxkck5ENkpsv9UqNPUzAJtsfNqH9ZmDftN1y7st/KNlCEyuNPi
wwG+y5ca0+qByw6sJ8OQH/1PEWWmOQJAcqbxxZLrszHZ/A2rH22ShNHBu3uQeiEbgT3XBIK6eOcy
wTsEESfZnXQxRf3rGQPLl4z6HjSwG26TvnSyOAz42QgLjlwl98oO8J929lJqVl9fj9XvvmhlMbME
nfRJekBdhKioNpyceTtAh9J8XNnX2xHmOa4lCAupSdTowgzxHmZH/YGHhX520+pKm4OTBvW1W07W
7rKb3hMbrAOhpTVokuP4v9Y8c92Hor0pnvaV1KJcKc0k0m1DCwfuiSAdtun1ojtovqwCLFzgEsO4
bNvb/gPCJ1Y6XXRslIfpcZRqQuYaKxoYLMdStR/FVmTRWY7uLlj0HEgt4U0LLEQBUXnUwf2bY2e2
jRWwchp0vwDP/G02fL+PeVPnEhxa1wPrDixijcx3XiEAlsM750maVbTP7M1Ct2SyNDSGnO8LANAq
jvmin9w+qlBDyNUfCdNi/zlD/cy6+uVYw4RalPUK7GhIGVcDKtJPourLbOYEINrW/EX7xKM0m+7r
L7nGJfFnSdVuFK5ZruFphmEgFw8ZpdQUMCgokkdHT5nw8p0J+tg/NnWDDmqKxSSxMvRo2Mc+nIfG
SxNPvhYqC4CyH+nOrFxd9jps8TmUVYulVaKRdbFLWwBsKXoZeFaJ+JjAquoesMwTFe03tN5xByb5
BzJC7diFA6/9P0D5iz6n/utFpDtIfoWUh6OvVihyV0vZ2P7bjccVP/Hjv2qcavI3ZYoXh4Qq82+s
a0bVI43VqRzfRawYib9/8nH9EwtTOWGVkvPLeWSLJxV+cMJ5ptmg/1n5TCmUOf5a//AdWhij6fvZ
nyKNTCEdHckafsVdFvvSU0mYwGDSFhHS0qlQlp91c27EmFAO18UxPflFcEh1y1prINVcN3vb/xHb
kkOtk+do8NRA7rdnr85ae9Q22JVF7ihoGsCg0WcMfOZkdJl6QNc3tD9IyLA8QKfS03kMALboqM7G
XrK/FS4fpv/QoMehWR/xUnqd7w5zEKBVqgGarkh5OOEaamupv5q/2vH7BrwloU9OQgH0w5OJCsel
hj4JxAi0Yfirmxh9x39CuhUwJzQjfhbjXpTuseC8TJRCFrV++k1+0MevJmSMEr0dVyi1QEIDqJrn
UZ/DOjSybh3F6ERS9k+75SiXw9lMgc2whmu/I3Y+7f59tvIW+WsdL1O3mGtfzCqNpubAA+3Rm1Cd
olieY1zMMD1QeHVYGWVsRHjJSkPQEDVXK4pG+GTBHWryqWVT2bAH7NWQ8g6qUoobDHW4tApVNgPr
27XDMoXQuRdRiw7EoN75aoo81q/b29glzvYperH0BxG7WH5ee20rKWhrAz+z0N/gYdYFA//LodwM
/SQfuI3FZyc9huSB8VKGKHejvb/G5DnRttHpaPAu9f1pn0hJwXjAfsN16tOypUQeLdW2RQ/0wyWl
C6MJFJ5mQYKRPr3+b+A/vSEDZ/OFG1fehzG6jFFQ+VvXpLks920/Za9zSrprdGD2A65vnS/LUa9n
AQlYxLZrXeC+NyQqtI+Bgk7PSTnMzpBWF1JDZsEn+m5hUlvLAVRxrSmBB892jnJnDy1BvNj4UrbR
yNB52c5idwnyVFiTSR2ObLXQu39Ls6GS9YDs+GudmX83O8J4w1BKMOkXmsUAZGHSiMT00Kq6xm0b
/HP3h5QBflqWxEXx6lSz/KGNHqLqOUcFS62yvDYHnwTKIC+4FaAqD33dgSLEtTSBX94jQ0H33z2E
TAMjS6fXNwtj6Jt3sRhAjwBx96slgLaU0lGF6bRVcgXCPk5517GWhdAyFQADUvtfTefOIxVwmEz0
tJWaPc6gQxtc59nK8TwfumQ7FFw+4VxmxvI0O/J0rbbO1Lr702zz7ne/WWoZf7J3Ga4/MDg2mE2S
SuPJymteioq8ZW+Td7EDZkkNZ9034fxbBP296Soe4bcjRf5HIM/p+aB8v6EmkErgW/EJta9vI1f/
NMP0qX2XUlcwnoLd6aADN+Z9ROpFAo0unjb7GaMPAWPJaElfoCx+8dk/MgdDOo/0wBdR28dJ/8F/
yO8iApH/w0iEcLtAWyUtbmy+7aHSxsEFLNs0wTz2WtE0qI+n2thIBKuV1boMyvz3PC5yPg+cPXhV
SLNVkaWrPvuvjX8t0acjQWeVhrHZxslIDpO4e9KzVP2BSgkviJMufTQB9iQSETEDAIRVL9OuRhgO
WY7DOPJ8KFgcjOcmfEgovrUz62UsnWSrdYZnbY84l3Jobv38WRErpATCKffSQD+PgG6fCFFPeqtW
fARt/R4qnv18+MeKWMwb+5gBmS1QxYNuYmMxu0Sx22vYG+K+ryN+Nr6zupCSjFldcOa6N0OztoYl
gIGEVrrEI0ndrWnLJxPPGGd1BLByo2410rBh/K0WWCQe9tm2UqmabCvXOJ5fSJY9eUq1plFuTkYP
9iJId/Weu/x9pZ3pJh3gRDfY7nOvXYx9LAJdsNsOyiM2zBG+o5yGnuo+KJ9odrQEgrB/l8HyOIxw
yI3qFX5R4ER/xRE7lh00127f3TJPZokrDow4iRIY5jQAhTPcvP/o1NdVYiTfAC9vXgQqIpYVzSTy
oLuDb0Nqs8ywyssz5PpeieWx4c99QZCcIBmn01egBV3OlqKyBX95GCdNb31EnWxDwgCM2yWi/Rfz
xZ02KxaHlaXTlousWRQ+TrYhUY9id7zBaTdZLfv3QtBvKP3Crtk1F/u7RYm5bUuOsyqm3e9zzq+X
MyHxTqD1ouKtUxKEJJP2INTQ7uWEfy32Iz3NFDBaxGHCnIKum7d2rYz6ZvyVxGVrUic1LRBanFbw
C6HSlOheUBmJ57tPMnfbbWR0wy5YvPTNHliSBWCQ/Ls6EaC7JuLniqXRWch+VfqDrkkGR6V/cA10
KkTNyuTx18JZOMDCf1GyuqhshrkKk+ABlpMlxqEYH3H3KPvgjKO5taa4nMnh+D3LmKOiu4E2UCwg
3qSIj2rqx6UAULru9vYwqWK+TgzeFfTjmJR/LzmGXbxTTkWVuMVH94SheJYAM1eGbASbc3YyTuzy
k4mQwytUfQZSWDD8M9ZWVqHOeZUOu/XpZ9fWMqK7nN0Z341rKozANlVsiXSsqOEhDeikic+ZjS3U
wkGsO/mvZPjJCEN27wXmTWuAFLu8pJQBzmt2d0ZTh/dDGZXoFwQi17/SMDicas38NdGcsfb9SuOl
Bentg/pqvUQZnw9pB4JM6j6hHiZqHrZ2PheSqtd6vrm52BeMbG2H581Ox+3oO4svUt4EHml7g1It
2nNjIKi1al3aSh4jmP3qH5jm3eedujR3XglRiR4HQFKb7phH/CbDx2AIM+PFDFMj0pQmvx1x6nXj
M68exa5xmbXnUqaVSXiDdS6d4ebHEx7aiuLBOHo8livqDdjEKLBQUMENJRlLlHkCG/cUfn8q2OX6
QXCK2iQM/4jugLzgxC6EXQaTrR45jcWVXreAelpxMi3hRAsCjwVITkf9iieplUTNWhcTJgyp10DR
TwPoTPUNp3vshW596T4vdlBiaRhzDXJDF78a/P1YR5NGVeWLlERe8YgJky3SX+RUGrvBsWVhC+ij
WKEpuXhtezGMvwp6sNVAPMXv73RYtJgQZDZ1gpcvz6CsfHQ0VH3pIW9UrA9oCCjaKq/u+JTD7r6z
bebsWzsmOaDPhIDKByKDY5s0nkWH6qNYyJbkhlIqKVrZUL8spV/d/G1qwLTff9Z460WzcL7etkj+
mXrkh+2TCXQFopFdZAht14Qwj+UFcSLKbHmLI1FxYmXv0/PaCjYVvcnMv1YsK3nkYVXN+1foscy2
d+WD7qG6Ubosw+887p+42GGHM6mNanUmPv5KzPfRzeqLSdKEsrenYLz+jDmfR9iJezH63CC89Ej+
BV0MxVuOqsysNTjCc3U+HR+sKVD0LIIQUPig31p8boYFo2YFjTZ11cc1j7+ZJ27mnvqXB6tRc9qb
UxE2dbVulTaE8LinpAluNeAS3UdiTTcJypSj2lPa4VYpi9z5piUeR+SW8Gz25MKjXP2PSCuvmLuz
n5J0ToHhKq62A09comD2hv0a00YWRGaWRqoVCZhYi0MXKJBHmPq5vhsgCJUa6lVF4V/3FW+CeaOw
AOsN/lMKzk5YpXzxjQ68pMZsP2P3m3lMB6y3Z4uq/2VLRx0knslB8e+5zxXAIn4tc1jybPTSnCJE
FASKZR+52msW76SFfvvAPoVWbYTag0ShrXltahbJZ0eK0iY0cV9BzKpl55PZj0aQqWkI42wL44/v
Bq8Jag91HP086ZvUanszqIyz88tdoLXCgyS/XRUl2I9cTbnHSDqjKJv6igbgBOLwqWmyKZ+yHjpG
UK1x0C6QciFFX9ARI3hVWzeugT4OMSDok2CwcpugQgO6ab9F4vXSFgz3OXfdntFnUsyDepK4WVIU
mDwHAZWF/SN48RHOZxwDnOYonJlBfd2QcYXsEKI3fFuvJeNeOtsOWFeqzf3ad26P5xorAoEEt5Hr
+NYAZnPUndWaqCXtYf3mVG0BXRhh8puCOzzVWXKBByw+ZY3yBCQIIx6Yeb3fdHuxooVgGfknG8MM
bNaeaePKZoRmKbylBbSojm75iOdUgPQGMpqOyypneIwlGyH9gsq6QkRB06e5fRVW4X6qfq/pFpLR
49KT0y2CZ9XfRS6t7szNCDy4pJLCm+VZp5TXt65IrYQBax9ZR6b2sBWde+yp/UmC/CWIWlJUY94b
OwCH092QWDIc2+Jj0LXN9cBlJ/8DogG6S3kTWE+w9GBbF80dxJQhLSBD64hh4iJybIMAPfLyYipz
BR1Z7Ty4mFw9b1brM/Z3ZnQdCJ+3aOSJ8wWFaCUKsCCWj9UOw4arpiJ/wBLSqvKW2akObDeTJuVK
Tr7nWF9ixoOB9qaqzaOBgaGwx9sCUHYSeFwV9G/1khYdkLE1Dd8nPPWHUNjaiWu9VOG8HTyf/zua
U5sWLnwqRnZ8cVl5wLgjvQlpBcBB3oya9lvBrruWvhf1lheCHzUN4SuSssiCsk48ymxfwsGwOM0E
g2H6r1ZyRza1LYafqYqDEm7eeB+VXlgMhBn0ug/Sd9Wy+JsR43z0PaMAgaHrsEmrR9gXeMn04lsu
opS7X0OwBPzKYco9RsRXUQN4NzCgDgM0WUcETcle7Lb3vjMkxSR0dUQUXH01fdrmMKgWbHLlM6iE
I3jX8vk8vApjEPo3ktnILvbzqOAQZoemj7ZnpXR6s/z52r71LWE3ZTm7VaFaon/IwgWxGUOR5MIx
knR8bSxSOSCdFtxfCZCQl13WdWShrfScz6ir6u9nT9Yzurlb0iOGZwAlq9EVlFOKvE7sdaCoyvVo
3p8joYWLJ3eNKh7Vqg/2uD+eVkuswJh/qswX05b5czZ4IA576MkrunGTI5JFGkBcHJTuiK6S7UZu
HYcSu71Ckkn/y7R+twhHQsScjpUD0DEp0DKoA4j3WKpdjAi52FACU/blgsYg9CzUNuPqYtk+n28t
/uVW1r7BWxVO5JU544hj9abxq9nGHiHVSL+5YYNZSuntHGlPWLUf55RibyUxCmF3oQmf99BYVwT8
ljNnh0XE5cbEO1PnaCz8BxtWkhDeGeSHBPt7miggaHJpuuiZ/HsgsS+AkMsVDgnq67dbW47vdcuB
TMaq/v17MFJS3XBZ8UZbyAbLMv4U4hCao/92TJnM8VN9O4HgelpPakLYLnM/9srLmxJQCoUiGGZE
LUWVHuNfOEA+zIPWw5D+/lNy58FpSeR9J1LprL0/0HpshbZYQppQuhOAxZ39Ys+ap9C3xB+nvrRt
U9jVhNr/ycpf2E3Yovdr1MNO+RRD7BXF4+zuEJDaDSJpHXdH/Ej2WSRsJXzbd3cYfQY9GnusZv+p
4whKce/hHbt1YAe+6b3NNfhlVxfG9NuwfrbOCSG2fy46PQPu572jINP7Nh62YDW4rLKv87mojlrQ
pVGT/CJa1lvvE1dVPXcbCHhlmzSiWVIfuAfktnkr5USO/o+ONbaP02qvlzp0wbQPzUB13KtG75xL
/jhpGECqI+5t32cPRxfSHQsXO/OyzDNJbCSxFyu5W9XsSB7mB3s4Bu1oIawkET+xz7f/DA5NT9HI
lSlh6xj+02B5dR+Yw+v7nDluQYN2eQvvfc1olEpfIO/5ncKDFL17XQcID+2wdUTTOWxeDT7c384n
AbQBldeZ90/epdv+/SVwUr3sJTGkXd0OxFJ0BlF3YyVoZO9jEAjHVQ/g+3bm+cOv+/QbbRZE1A/I
SkUP5ZzBWAOXAUDSMPztPx19pJ8x8QHca+f2kWg9P3TFSnu1EXdhcS5dsJksZAAEa7xD/FHpxuxi
Q8yYCGL1JW9StgjD9I/fQSlxawefX+PvVtL5h3/21y0dKQUic85FRszKLdNINIWRIyJCHUu6nvDp
+9dhD9LrXRFI5fFF+3IIEjiixn2KXR+Sg/x7UnTGNs0EtpGgUctsgYcx3xbvf5ILhJuB8/lPvkix
HXF3GmyK21kYrir0CXlqhDyAry6zS8XhhYd1MBs02rbbJS7P78aCsClN5f73o6sLRmVJXwwtyb0S
QiXYXaZJ8eXxFxatuTUt0/8aGnnqtt1S4cvJW5bP7aSPwmpakcAfs1iwiNw8aChy3IjNwlznl78f
8C+p3Rg4Ucl4W/7gmQ669kLw9fCjiXtGxgTqNyv0GpCLyBc5jkt6KAJrCwkmbCQm1E4lZjDHhsDG
c4/kFAeTy2evlFkFX7ZrUwmxdE0+jzm3R8lGbgnOMG751p/2F8LwY7qfuGWCe6E9Igt0w34ulrtB
qFQGEpZHtVmSsqFLEO/WO+QgHiHLLdbIwOVjfJRxxTtyzfks+qnZv2uDWD//tgEkni5EvncviPCR
P2mB/CtG3ngZ26fOas7NrVjELqE49bmjeawppK/Ku8yVDg+IfeR9ItVxFRT8vcZT/1RV9S2p9o5w
gYOhKozmIiKkR47LBvYrqGaFlokq+Kx55n5wjkJuPe+FwFk/1ldrljQ+vkFdhuMvYMrrBzgXX9po
Gej2NxjLqka29Ky9HYU1/HXVqN8RBltukJudv7yfp2mI3nEUcHx7PBsD/Knhd6dMTF/fbVY3pAaO
Jhb7zS3kG4KxzJnsQTr4BINj+HxspgnTPSo6SeMb9KufP07SqXAljBe1PM3gssOUgu+WRVTbYLne
6qVrTkSVesAe5r/XiBpeKYWEqKKjF/b3qZEMIqdXz020ewcdwodWxOKPhli49rgOmKFWi2rKEZGx
OfTB0eyqgttr0sm5WQHa/H/CvbAPO3/6dxIgBzAW3LfH3bCNwHP7gIQ3FpiONB8AMhDuwbNCl/ay
kJ1sdIJqRq1930fH1gmAgvizGN1saMFhUhefgb3+dKEWWsZ+/y/Y47RuIqN1kjNMs32T5Dq0GTW7
cxRox8sf2zQ3TXQurrhVNeZWYOiRz6670/7uC2qHscSTtMI37t/aSurScIKkjfKMCLyhwhKA+qS3
cihVFHixo+7snahU5Q5F+9xVv2wErA3UVtqht3QFtkS7fp0FLOVEK1eo4aH5CNfgo4QFJJo6IaZU
i5r4vXIBuea+zmW7wqooC6Y45BCi2RRRcRGx5zLQekCHFCWMN3GfgbAEqtd0/kfumwrhZjnt0Uun
dBNQJhyoz/Sdsth8rAhnHOAxG06aOY8pQNs5XyKX6uixsoqOH9hVVITuXoAxvGAUMwh+5AegFwrV
UB0uZwPMuJJ95XlqEBfQ5nTyVROZJDnKCSzDPtNerUV88RBSuFgJD73Io/KG4cIGMnEv0+qfGk9B
wSWiTtgpRtHTrqJ+zmPcmHIyv2d/xJe8auKDdzIepyJn3oxFVfB0NJG4ulQpIk1xlGGtXUUbq8Cf
rkYUOt4uUdakm//+rPYEY3HWfs/Yqh33gKsJzl1VNGNRnazpvuR3DvXAREy6wB7le7AqtEB2Y5kc
zAFuZR756m0g6bsm889soDvEjWF/4fNkAQSfVpGKlVTxU/TdKTnsGtTKdHAmz2ZCb4E0bCEmCyEK
UpHLAnv015RZZ02RYxuD0j0FG109ifRea+/e/1XcLRmxRdt+jvwyXnMZv341FIEZSSZuzHQdOi7i
uyC1w+YqPcYw2uWVPw/bqq09dvjuoCI8DH7aZowppJDwv0MU+OgKGrNFgnguV+4iHyJtKGDNNErS
VOz56s0Pbh/UhxL2+9fM7jeo+nIIk6FwKcEahn2CjY9HlwFxMdYM9RNWODjZLmbPY8EdsKJupsMj
XnMZTGzj1MuiplW4qvNXwPgJK/VWx5V/v1ZjQZVfLWZQ+RdMEGQ7MkvVhKveXKJs2wsafd/HQLIJ
TAEWsaU6rQKo1VDanwfA8qcC3yX7lAJfDvM6jTgbI5maXmcEQdaTrrSUFD600+K80KNuFXynu4mG
GuMKMQDIAMYBqL5L2g1gCPHh3+bfc3EnQZ0JZlYPe4r8urCklaxOqtRdq9P67x2sGfr2AcqWkU+1
yWlkljZJC+VwycqubAomrshma1irBqQVjFvGGBiuSrwROH3YjFEzaksepoezogm1MecUWwNXfFXh
HuuhIpVFJBmYuarQhOd7nEP/suiujArbLSxfVZCK4oAvD4XY0+rUhGcQczGgMAnj37vkfFMopXH/
Fy+s6dmyS3KEaWMkgQPuva4O8YpOsTwVLHc2bwQ0lPdNIBvroNa1llDUPB8GmLlwZR/RPaylq4ax
rvfybxOjqC7zkzukzIGlrPDvYEnQxDltqb6xwWx2VpvpcXLQsOjBXG/iFX6Sc2AQun15pUjS1hn9
uCkveDjfYtUr1cOgKqUSCpwXF4g2EnnzRPsYpcF5oXjiTLlzTCfFrhTAZDcAzjxfLbzj0jJKbiSS
0cvwy7uoK4r0vCzN/XbPFdq/TFJisAo+cobyJFZxrhRzI4LQ3fOlZYIOq0PnGkhDTU0cC75Fzuen
xi4+rtczJMIlSXYbjX1ptFAvdlDgZ8bqsp1DJdFy0ytC+MMC4cdCnmoJy5jGlWmXjszXp11BfxTN
dbwUY5aiKq7TdSfSAafri8A+u8jFCpPH6TBeJga7frxPzHjir/gMefZQjZl+HgpfwUstnIMgy6zj
1c+dAtIo5NsbeVuOqAyMkEsqBRff3QxPMaIOf4LVLIkengZhyrkSwAWAdHLtbvS0tsa1G0EhJ+ix
VMmrskfB05Wm9C9wxoVuqhdrm2WAGwO7CPjALSTW7M2efRXi5DpROHqIXPLeejcaBGlvy15Vfm3g
KqwAiXoT7aQX3MlKcWtT1AfJqgY7DJdG72QyOkPlMar/c/GeQ/BNPP7yPOO3AkSiR2FNDhjEheIK
qt6N+AjN6tA4nheKvFxmzWCuY5UFzhV4uPFFd17ePqw3r4t5kTGhrrHKqXb2f0IHWBXrLVKhmclw
Xv3TxbQvk1mlB6NfwXmOfTBS/s8WSInh6KEnsruIt+rJqPKQZaGSP/bmQLrxZpTwvT5NxNXs7X2D
rzFdTVQAb2+Zc1n0fmKngrp6ZGIy8RhEMIvrYO76ZoME1+TJ8kzh1Vax89lvyVZzXH38wMht38kz
rcorg/qM09DRXL+s45dKiaes+K9+6SCn+5t9pDOdIiicHp4GheHZVUDQSkztklSSQY1K0a1O+lwb
crn1B0fxF6wUin92l3KoM771Uw+pZ0+devcOl6bff6ZOcv8D8W++QaWwZlfBGQMcEa1f5iNMl9dn
DErEXoIqiFj+D9YO/Bm+0VE2ZFUz3fZp+lWOapBNM+2Imx4phjFaZFlluN1I+xVKqP8l5/S9caIe
QTiSMHMkgcIXpHLj/mKllWX9qfalDjO5/r6rOHzLE2yus3ec1F+xXpwBmSxCY9x9XSZMKIVuek0k
5ZKpV/41MPPtZLzMIK+RzuW55OG5xTStvg5P7D9/8XZ3UVSioi1EbN+bjKf5NLsDqORsg8lsboMi
3s36s6MU5A4L97vLAZsLqspsBU6t/glWb5ogv6OqmG9DTdS2NFDpHJaQPsJn4TeVZBH8hN1HPM6o
N+VgcTjE7wt270xYUTzHCYkJsl0GzdGPPgbfAZ9Z/jqYOcD5zYxN4e24hjP0kbNNv9a3gYhZ+Yh1
C4mYq2AKLAKtx/1u1lxCu6j4kUmf2x0/7Vl9GGL39ZZ0MLFsdKB/wUOUW7U1/cUX1R/3MxfxBaKK
bcKFWlX/wQFrf++mz2OdjTHEGO4JDEv7Sr8svjDqD+phLGxgPVsaTuOh+1CLjFTDwBfOt9eG27oI
Jkddbtpo2vW7dQ2iHtwcfawf8Ilf0xQ3QQ5kAU4Vs3y5saufdfIMHTlYoJw3QY/BEK49iTqr6HMh
8f7N6uqkDY5u9IxjoU5js7cKeZRLSxtMBMzrD2a9zxciYcHNZRr+V0yOXn99M4f7ZlUvlfvMfqqf
9a4cT8rrbrRAO798ITfLvs2sc2rj1BPi99QYSRCmNdjexHWrHl8ZMpGZWrC9guk6N9n4o31xT8t/
z0htfJQyZaLfkhocYM8eb7N+P2tzj3sG/xlqONVanGHT4/mQmY3hLupd2RV80MuIy0ucd3DkSPiA
1SO7WqhdAsTFqEOZla8XOLH8h88e8k968Is28kpg7/hjLsaIT+AuBiWPdH+aUy9fjUgBEJnbYG7Y
XCG3aob3IZW4/8g98+JJFR/eB8HWtsnow5o9KAGVtmYSZnHWvUMuIP1m6/dI+wUtPyw3nfQvRY9h
0ZL8BrcfH8Ixwk4hEv0u/L9c7ypwa6I23fWYcN+tl6Hv8N0fBmEwwkT+kZfKqGIhPajwiXTAXmom
vk8mcg3YCUzalcjiJbEDoQgGCaNAHSrMfqJXl0RLI0x7OsdUIsn7n1fa7uGbFSKsZ/VTMN8sgm+B
B7T6RoHigW8iZQb+696w8Gw9e9Z0SV8zZVCNzP6ErJunKErbB9MfqtvBC2eO1azXtNqbM5K6nrKb
C03NuVvvEMUvRvl0nuHVVgLp9uo2b1REVw8iNrvTZLhrQbs1JxbcsVGzyNwnNYFKpGCDx+quJnlB
PZI8CEmdipWwUcjafn0S/F0NTnzWHr93kfg2FCOl/rpgeQWyhYW5LgEIgCA7lxCrdhfcFWNMIDV8
CxHH7Vih6c+Q29vrZKP7ylPCCOFZwBYrY58ObEdB9ls9tqc69G1zhVrYRkrdub7/gWc12ABWTlKS
EzcmOq19zN4+nd04KHQKj8Q4r2STxkHYB8LtFNGwiOE2jmE7Juq8twrkf5SSYRHeGvNCNcOLYtJo
l3k5+y+IZDO54BmgvW9WDuELcx+tSe+2O86Xp/Z1DlYWOLVVH+a/n2qjFOtbi6wq0gXOD3/QqQDn
Mxr/9NLHolJZ6q1CoathycN7dh4yuQuLzmUyFFAm8YirBMEkV4QzNVKH18uq6W3dVjQSdJLsXHbG
XDJYjlqvTx9ZjU8w0KbQXugrhmUsf7VK+DNcir8qVuXubJ2+hWq/O+emFmCii8WNgREXUik1OSVC
lHbp4zOE68MuZ4zNqW6mjcKdybJQ5v0t92oflOH48Bu8qYSpk9bmzBqMN7H30/JAB5Ukjf2tBVps
mUkluwGdU6fHMNpv1hGvrY+o0Xn6LXHnGCM77ekoCWDX+nmsP8KpXi9BfuUBRqeCxtzukRqQwlUu
dig4X03eDOeOE+1q8S262zm0SSgeGNKoBKLfiAYep8CrmOGwUpOUd2J2G/q1ZN8o9drf6C7Rl2FX
sJlsL4v1g681c+va42csCEZd+ghhujBZtPXZvKoRep7ElvwR+K1+t4/jnwdb1MuDxSHKv/+zhMwG
Q1kMzvzVRzruAiPyVcTYgSPek44orS6cirABC9zqE76FH885nGqKipv2trDucDTGxmtOfgZQwj/c
5ndQ2b672cwm/t52HRyVFhIhS2+DTzKtqdTAAHSyQQFMeETLlA9liE/tlJFFCnVD0ytk7seszPhb
OF0840oX1PdyMGEjs+6R8PM0swDPLeAfdTNaR7KbHlBxUSHcPajzVP60GOj0YS3Y9a+CpeJ7j6ZD
wn/hK3dLKSSB2gO4hCP7cYKODnqKEyQs6EItbrriwsNhlK0mYNGRGeG8SodNJGo2t1T6kqHv0KMI
0+dXFozHM3znIkM8D3e+iUJgJKjDDixWahkbG4gBER5mH7i2f96aTUdlCt6kkFJIFFkxQrPwF2vZ
R0p/HBvRFvy92z5VZcunwaYQhbd5ES+l+24gEJqM1NuihcRWAK8cQofEuouSZIcJc6aRFj/fBJws
xWa10g6Kj71QsCbwZ8f6/YtTd2K3Zm4fifdbXnIetilNg3S2vzjfE7wKbkenJtioOVREy8VWwp6g
MWLejuN1P60UhNpwgWXgjH/LQeG+spqlcDpYmpxKr9Vce/iJDHiOtYoaKfvh9HecSb9jetTvOrB3
+2KGpmHx89zOh14isKSS89r6U9CcRd8P8F57xjBgX9sby0hPCTQeiCo79KJ7PCLdcs8jran24qYA
3rZe7oEYOF/iwlrWgNMQR3sG/M8Ssz7H5SuGDqvlytNn15F+lTxyAz/Qd9ns928l9uypYMGOdpKK
ktSSsWU3sBjzKKS3bhtBhyrUQyYXU+ZUvLb4WQHIlaVv/PWzp666RxjMuN3T1B3GC1uvh7ldrWj6
vLGJ15m1WGRIws1vh1hHzCC8yrUkYu+M4AGbipylkj2JtOu3uHhlRj0N9Qyoy2QGYPT7VcAnQZjh
r/EZVixNmSvuV1zRkhP3BN6PqauwCsKv/egtqH259UCjZXgGDoqdIqBihZBp1enjq2JHD1R3Q8ci
Oh1mMRJS/vtX4PReFjtR/wULrR55cG5vNimK5GHWGW2ZDI8w1vLh7n5n7mW2/VyzvjmhD5VUxAi0
XvcMc5iwlff+JoY0WTGjhbr8EoZdM9F2o3UjQOKpSB5s/IyoZAQo1ScI6dGRY4uFbsMvYsMumdoV
hizs6SbIOIQ2Xo8BTRNsIUS00kolaqlMAswJ1aITYXT1BXBVLsc8SLDTc0hKJNUCcA8BGyVa2kXI
vyFIyB+3OLid6LK2A3jsIUNAlAMZypH2o5HbSbBvJzTjFJlssc0KPmLFLqoNQ6sMx/e8dlbsl00s
UyCaeEpu+PzR+GKTstgBh+SOADQ0ITM8n1+Lgr4dPQfCicX9i8Aq+VhfraOl7dJDuzUOnn1ts75G
u0Ozvb+dA6cEmoPvWRlu+r2SLCfyv7pEPpeA9jp2iYvzhWPeM6R4gh9JEkdoZxQrWEsydAqAObHY
3kWCFlqDQtjMzdtxMymw4gxWA0K52NQYN9AsUTtxrnIxpTpMB2QOgepakSXdlPmR3/8iAv7iNaPg
GGEBM4TIOGq03LJZfhFUZj6VT+ZuljABdcGbVW31lTcG1CgiTYG/HqmGP1jfui8pRQup8zsINpyw
wLsreTI4oizxDej+04HF2NfJB+hpzlQdL4ibobVY2JNBwStnBHQxymqxVRCND8XvTTpL3VPfEPDs
frVYn1KELOKBP+LigKI3xbku1ptAu+iOuVfg9MYmKJOFfKKnGaNnY+3M7jpse3+jlVE/6vxibCU3
fxTFWXyZe/78Jr+sATXx4xBlICuKIJ8AQK44wDKs6M2k7O0DVYYA06pDRuFBmoaO1rmP9g/Aq13p
qA0PKHh02QG6+yjX9F+KtNqgC1PtuLVTyAgqXZV1JWI3b8ieFQnlthH8F6ryG4umP4oQCfBjDHVd
+K5r5WZk/Lzb9PZoM+2jc0CGfe7Sha18CTqZL5LzdgqwcKXBM71wGyyq4AJ8ARm5QF14p3P12Gj1
j5sT1bunvozDsTyob6Cw2HTBMgkGtqYr3jBCW7JQbEDsi3kP2m+FNeZKLOCIN00vssTX7mwhSNJh
iLS3f1pTxjvQqkvw5UW88CKGYzB4yGS7Uo9HY4nXxJGihie52rrYfpQrve3URMDd55mEaNSu8M+K
Hu6BMW/rQhffEIsq+bea4MceShbhBSAXI8Uzn92pOIjNqmR3E8YOrEwKNstlEf92jzhuM6RB5gA/
By4PH0Nzdhtyf4uN/WGCM8tKGlBAoctYIotcPxE3BbYpsdU+vPFNQp+2S8AvmdS9anuwXhkEkhcV
wW0DlLMY1imR3hXiF/kVt3qduUsc+RuxDPHkO6Y21rdAaDQayFD6PbggqMB30lMBBaNCf+wNUbQH
Y1xr15VH9+mvn72zAq64mpXoaUB851NvqZDkxJ9wsAUSVjBU5B8Ef6KaoGt9ffc5WySJcC2Yb4Gu
Yu72KUThezmxuARb9c/oRzWDb91VtyfYlimckk6Vh3xosqOYAYmRbamNXBzZSWOUDSjyBmEY9U2G
MWSgTKYsCZZRD7pF4YuOoZ8dun6oYwTiFZmAmjLmZ8QMrwsuC4nEqA1X6TOt2zeA/1IbqrAtiwi5
zsUcYtZ9VT2p+U792FfirWAAV5uHX6QfB3QPhYUvvGFD/bWjr9+5OBE8R9Vi34zmvTquJlhPrqC6
Lw+Q9JDQDUYdntYbaAbyr2Zxa34zSnhR2TkiEI3NPvBKW/XlcSFp/p5Dw+LIS67Bn+CA8WsxYUtj
Nkd3AkJqTD0zxNQU2dntKxmrLG1Q78d+5AxOzBfXlIW76L1f2o5MmGLcZOTuSRmUxmmuAi23rauD
B5teUZcW9HOW6tFuBFenCjX8vV5v2EUcpzHXt7oiKgDV9b2ySuzXdzhzGizBVgMQGxdk4bwBfv6b
zhu6WRuj794Gk5VyvlVMifGTv4AAMhMSqVAN6jXo/sz3nJrs8sKBb6N5LuKqOk76+65ZhIDNjp9c
VNk/JnVw+LBbGRLmdS7XEJM5D+JkwBUp5xDvl1DCylyJ7ME3DneZSUIWNkCg9NtReepmb7EyFVGa
tPKHTsXoM5xYUbgCwICfiFMLStXD7aPiNvbcHbYrRSc10n5wORixQaIHQQkguDs1912pAoJDn7Z3
2aNjuIW3zQKedz58XZt71qG7XFA8GiZfTL6SZIZi0BXfd+PkxlLB3blFPLeLAb4F4Fwdm53S/z57
UyKOEMQNLXVGkw8fXnUna9fIxNjkUxz0NZXItF717dF/QBFB0gRRrEwnpwaOJjj1jnuEO/u9qL2K
EDPC+mWsLRu4ld3vTkoipEehd8qFNHOSNcm3gprb/xky9boLGjTNhEVJ+KeiT7MqPz1oUKvE43qK
nKNLNkGzjRwHece6DSxBn4KaoOudE3IuqLC9+ca9WQ5waSIZJ3WTJI8US1om1wlK+By2kpto+2sq
/DoNGzDvWk5O2uIsADtp3wiq16qVow/G/5vxxkDrCMu3913wXs1/Taj4sxEN0n/WXCcH638Hkdj1
s6+HEMetdUflPyZpQcx5xwyZH1ZgQ3mBpKnmYLE/GmQEgNvtYgJrVHJn3WJOJpF9BX2wrgR+6jum
a7Dm3rPSIDRTPlEI/L8Izbb6vxcLXmtbsndmxxUUVimmZcmlCnig2NlINDa9xcJMKmrHJUJ0eVye
bTXNfgYDY1CEzrnMIen25cl2AEjXWWz0kOKvmC5WbmlvCS7EGfWudiKAAoM5qx+HVnbAjtrxjXX0
7SWWW0ZMOVdGFK4Kkd0qs0fvoajcvdsvTU2ySe1W+UcEJoZOh/aEwIs1hRtBs3TRZRuGtyjTrcuK
XdRmaj9s+rploSg8QeXqjpwZcozGtfeH560lljaWAEnnnVk5cA7UWluI5dQUi5UTTA7PlCpD61hI
cCCj1+VZGseX9tBcsY6xDLOyy3pcncytWNZ19FuyUNxryBH8CvlLkGeTNmQHtqnmSImqj/17NVGU
bAozWOnojprs9K8Qo2gYYKgoBq/PSk6ZAtpjQ/Wb/GMmtj2LGdudDaFuG/rss9wqGj+EEYQOtoSK
VSUCsnM0iGl1lOMWNYUgGhEg0kIbr6NnSzF3wvmuW+yuDAzKWUmZjAgeFKmHsO91l8yweKBku1E0
9Bi/KJmekz2MuehxlBtrnhooXCa9ZH99E7VYvnrdJ9DfF827l4pNhwmQsDkV6JJhDe0cxeGv2M8D
aylbatCvlWNTeWK6Is/EnjLH7hKGrwI4C2Zc5Jzi6gdrdxKE9YuXE5b2td8kOkxFnzzCSXlXTTuO
dTcMWXQvHhxcitSpONGAS6YSrYSECTGydrHHHkLvrR/O3f18ZY2Q1hdxtet8bVUjKZ4wqob8vkBr
Y1vIFmrKxobKPRfoTIwKZEFKzP4DrAdHaudBEbRLfIcflS2HKRerRJQzT0Ud6CAgjgBdtiRTzVTD
rFBUAndGnUOZc2nYU3GPAeoMTJO0i7WnkgiBIPiNvSNJou/IMvrREOm8OoQ2lx82urJrPKRRh0Bh
kRczCZVYbY7ymN30gr9mSuMTqk0Jf6kL8jQK6MR2m5pic1QlRiakXTTI9H2dpqW4hhlj4hOhk6l+
8ezX9iyGPZVBwods30wXawgN+EUhctatR4x7dmz1kIbgijA/EHJcglIVBaG6U1I/7EbaOxdRPHHz
Nqxtu+p5j6AyLW5bofhTx8L2dF9yAZXksTJkgAWokMLbAHaA2UPbnqYqLA6/urTAVwVZ95t5KIo8
Tcn89eDRHkIDaGzFvYfKIXFPywogm/hi4+NGS2z2BjnxL9v+tZHSuf5UHD8NbGZ5NwN4FJDhyiJE
8tKPNhYgUPKeYrnpeaU0MMm8zzsalGeGAr4M9SQ0JmnX+Cfs6XRcMU3fBsYEguB4iyyef22OW4KV
fYq/qUj1mK3k94vjZDhyJkcS/5zO4MNBzhCRTMlp7AnKzaEfQlX9snvNrMIDLkr4jSoQH7WD/75C
6GTO3WbHE0dAzdcxSHz0OYqPRsKYYo/Qv9Qxk9gOFy2C8yYoCTr2oCXHTM2qAUQkHF/x1p7g6Oyi
yT/B+GHh1CJvaWIaM3ZNnwnva+Tvy5z1mdv9/Sbi1VHEVivk/UI0pZaRmDaM9US7jZk0xga/tqQi
QUgwkEwpfZHZ9ZJZK5x23cG/dwnKgmxnToT/D3U5EndqazZzd52Uqw92bQfo72RoIFwKc8KRZgmR
4ry4eKjLFpBGACylGTitEeuKvROAO3hCyw92Z7Xc+3Xqcymq+66aDXeEzX+F28JZB9SiKjOFF1sj
r7UV+f0UhgQGByCSM4vZO9UenywTYmvJQplHpVZtZKyxmlr4XfwDr+3eaQFOLDkSsJNkAOrc2vVs
T8RHxTWE3YqOJAMWWs8L3ob23r7x9bqeXLMIxUYWlDgL0w6471nKGInu1pqpWaQxKQTlq67Q7krV
GErv/R1WrRtgumq61vS8OKaWovjNbYUGR69gG3Dtu2rzRlEcd2kvOzKzV3F8XlRfhYYNreG206j/
b9e80zjaTUepHITWKjNVDCyXp6eO0zWXctQdOVIgI1cm7Ower06weW8A2oJJMt1YSsZ/fWDNg+cR
nKPkK3D/h9K0mt4ZFk5cjao1h4Te0VTtc+gpeLIZNqStWSJ7FbxPU2p/LMB3QxdDZpnMeG0Vw1ts
Ht8jAdCuFfaW3Z20/gD9u6Zybl75x6ygQCbpt2BiqxGQdwM7xptM+YgnXpF9oSnJEwXWhaw2lncJ
uoJEY9xL37JovZQdRcQDG9szIjT0CBv/ffzm4zpW06FhcjUhkj5wsIo0IA7+GMGh0+La+z/C5Bd0
WKMFFbFfLnd/xRgwDwbGpNNIDfESW7lSFuiKpE5D5eRblaUc7AApMo/z6PUFdXipwyD+LrRl0YVy
QGAjaojHQpmJn6NLgetweGm7lqRvLtJDDkZAjv2Tbs73vI1x3j/XztzgdmeubWfAk93t9HyFoDrT
iagiCvNmu86/64otTQKrvCAQYua72aneiUVvYF9UZ5wGyozVR5cWbi+rEFFhHu4wH4bjrHda1x0H
hg1m9g1av6jBQdFHwzsTJNFjvwPPQCUSOmq62Ddzhxm2nsv/uolSvxK4YLfs+2I7ToiXjId+d8FG
+92muT7Zhw7yoFOSUcsXFciRagedxQ2KJsvzWHdio5AkFUCTvsBUNUaIru7HZ6auw2RCal04R1R9
zG+pY2m51W0F6Aaa8nuPO6ujQ+4Vlv/ucaGawVgEp+uRyhLct9Wu0AY8tPUtIKfh3+Vnt7IchCUK
5QJ47diqASrVwjDfjEhkfCKYdCM+KDrXc5txqLg/AD0w7N3+lCZNVdTe8uM/F+Nk2sNbuEmAMCaH
YpPMVNZUrDGKr+HiHSEbyVmrTm3QMGfoYo5a55KKxLZrGls47yE6trAHBgTMxanEeYW3H2aB3FgD
mIexyBOcthdqGaA0yq5FJwgUiJonWFwJSgbe0MNgQuyOh6pHYly8xV1D1wTvbnbGIEtQXqIZjcnO
aH5ujrXhAxImsTOgeYrvNnEzAn+vCt2SrBPQZ5V6yQIaHCWz4iTPyszXTq/X3akOQexYusZaxjTl
hp38Lft7MYyUDjGdAyYst4MFzswMlJeBRKxw97lhcNEgi2WUciTBDFNgF2NsAyUKylJtAiWZnQ6V
Sne98ZhaSRdgG0cnCgM3Wb9kvuZHFSnXKuWCvnj9cnZBEIRKkjly9iYhSxoH7/g6pdIoXGDwIc/h
mQfGjw3sv2eKOrWnHMFrWYmeBQhZRa3onmYniCh/1oV1nl3H+wJowHzq0nqQRvI5uuckTnjlnuX0
Dy2fzB34xpQMPBih0TBc1vHJAWvEnRMLmHVWtCjY8KiX5+IHepvUXvsqDXOMsXkQvIEjEwUnNEpO
Jia5XPadnm43QPF267mNoILWGHs235c8Mec4AJjZhIefabcpR0LkYYysegFr2yGlFE8D/0e9++Jy
gM0YoWvQcJxFGG1rhgklu4R2oVaEhoqNMrI2knOrFkQcRyDhwalJoOuJuT9TSEp/XpxdPjnUNm4C
z+4XwsuMVKBXotybtLHTOKFgsMeeUARx8dtibxpBGUB8SDQVGt+pwSKTx43UCOKlwiQoJF4hFTJY
6komZAzrcZeFGZ+XMLvBohkkzPOeRZIgQGHfHS+6JBBJs/lKMFsqmedN4373cBoqX6HOMZX9aGc6
9cIaCtIAqKpkvKfvJTPZ+iERfZBANHwp96BEDYpUwmcDNFyJAKH/UzJCr15y/LlY6BBpQ033I7We
eNZ97fLVMWCMVI1m4zLxGecuya9Zj0O3MoNhitUGEiIVoDzFrZ6oQcw6JeOlk87AvSYHKRC7csPH
1Ky6hwTKPPUprC0waQETzn8YrUGMv+wC2nXhazw88wBJhh61zEOmXKEevXfvU+4dzgsbmj31AU1p
Oq9KnTkpynZra7jkOzVbLr0jHUVgiM6smNsNaFR2dsy24olR/KyA/re9kcYV2aqrwDRoKTKR2F/H
CXrcYzfG5zazOh20zrWHn8Dqf3CEFmwq3p9o9AI0z9rr89tf6WfbujcBXZn6Ql5cavw2KE+hVTw0
DbxAZ2PPUBrfFrqk30Zdg4jnmUhkkdz3fnRnrz9MNdkZPCu9dLlqlUC4w3/uPPU/JvYpmIfC2ZjT
fxrMy4XnA9BS+Z+lEnWEM/aBeSBJByykspbmQiIzcBY3kb63kpthz6JebfyhQS0yPCEiWIU+R3VD
M2IUlr0SzXRW+bnhIKeSZLtsVJsRa3kZG4JGVu8GXltsc+4AqBDSfQO8nO59V8xZJfxnGabXusSH
flc2+3EqC8d94TqLYV8CAe0VAB4YjrM8f9RBqI0rvOPPC30zoUPFFpsU5ledxXHp59S9pi9O2RBC
Y03eODtiFjJ1+WBg9Y/V1QmrgO3ymiqmv89gqQEaisIUw9g2OCUap4TtKUoZnaeLG+u1OtY7lrl7
1bROwAXMKyZf/tV2drEYFCzsKBCajpE9K1Mz9Rxxpr2w4KD883xHeCerru/BFDf58y9fpKC8tlEF
9214idKD1D/zVqEtt03PDSY8JGochoBWUCq0NeKoZYD+7/TfgQdyTnF4ixeqDQK4rG4hMluYT6fr
jPSFvtAI4fEDbWkyzUt2Nrs49cGM5HojDRmpKvfcVj1kegS6194eXfkCx3s7l4IaIGd1N0llbQ8P
eHGsl8+BiLFaqb1wFlr/hJ6MkpUARD+zndicvvR4wxdHalvN7PhYS++4wmeuFsdBbtcA8Wf1I/Dy
63m1fjkzdR7YyjTEywx575GQZqbGmX7PX/F5mWCl70LIWxTZtpG7/c8kuEwY0vlKS7B53aQIO+wI
2um5rNocfrEMdKFviVOSBdgbWzOEY5t4VqsIsuql+2fchkTqqUJlQTDBrk36uWXhdl1StCf5WRNT
JRvqYxGOxKsI220+AhUqkgIPNgQT7KMhR+8mstj/u2eCvILuJNtyZghwZzHhFoKbESm9Le+wtGHC
Wa8yx52WzJygqtDvEjaosNPVfD6pxXaqzFAEedOXBQbCok6DpF7eYzDNRsTTVDQ+WHWGugaSFzD8
0DiSfPgG2dh8DpHwb4RQ0YkqKwpO3CZpgSS0kQKxGNIB8kVaFhfUfl0aRWVaYY9VuohLBo8sdCDM
od63g30Mmiu3b2FqZDZYO4BcpBvrqj20luJR4iFZ/6lFj+0kGRSR3e+UVELrPtpTwxJvFAm/1ZVP
7XL4qe35oEWo/91ZaD9Q+gDszXQ5n46d+lIkpvaJFfcDIt31X6gBT234fkTcrDyGozny6V/7Q4mf
aFlUT/BDS2mo6ktysZ0W2Ee5lUXga9MerxT557wzrIYkDfEU5VX9DJSzuAUFDWwjoc1Qr2GOTY1L
D6HR53MSSBDcv7/YwPlfXKpB6DR3WlCBndIbx7Yq+D9Yqx0XCOqlsHg0DqMBA1jbgIemARvPfNh8
7msPCgvPs/wylTCX6KqDQ7JtwglgdyzFNCd20BgJJUA58fwEHFBHh6LhcsRx18EYILtAY4R+xAWD
jvZb8Vhc4X28WkojuV5fMYHvCkMEfjcTVA2vZBugU08UCj1Qksll4rWYZZJcOaSJG0j5m6P8hiZ/
QEvFuEdDDJ4GHtPSBT8lIPxTmEtSPGxBNM4qmzIm2yN+xv3uKS1zRp1PWEy+SiYsPXGUkELyxdct
25KPu16ZE9ABz+aiCllIb1S+z/BfY3NVgoTzy4e0A2lPzuRkWk9BqNOkW5wIxfzSYLeXFdjdg5of
fGHI9G6iW4HnI9TgW3gzZD8VWB4/W4knsLdQTnfXoybQAkMt1R9JkAWdPv1jJhsiOtFqI40k08fk
Xk5qKHqaqwBl4TlCTXOou5aIc6jz+mSauEpyFstk3Q/VySAWMco4+3oUqvpCTEKPNmlQJxGSLQng
EKBGivHFj3E8EAvq6kFnMEE0OBsAVRdd7vfQl3jAX6rWK860lpavF3TZGEK3o2y/ikBIToS/7hwC
CSTEwI1q/v0GRknpnvlksbLVDGm3Vk+Qh9euqeFcIFRDuJgk9/5BHqWWycw0s+AKPq1kJBIvUjNm
GCR9Srv2QHUIGzW+e3A/8feT9lFvq2HDPvTxIiuLYvO+zLtLpAZc4+m/MlQVTQNr1dWGGRiofvBh
n0ND9AM/wTzSo+hrmPBzbgNQ0YJFrrVSOUzWtE1PWTnorrPA3O8rA+AX/9Fzzv203cemiZ6rP9MK
ew47fdcX3qC+oq/l3lkNpdF7TKOX3DPME8nwv+dpPx/VFQXL/PfZ2vceUbf4nfDZn6ZkvMvLZee4
I1Gc8GLfI5lmSk94HCwcRMBH93LhC4zMQPNuofZro/pWQbbOrFsvWkxtSCnCC+LC0cT4B8nI3WS1
tFqYiPmg5DxqPRsD0TPHmTS82R3XkAVObrKOSuakLgri6SN0h/FI9x5kxOjfFLWaRqVCfp6p3SHi
4nNdypLrWaSXVvxjctkMX9aVzcKo2euVk1aKgnMp8eMj+VQZkhT33H4HP212MwhJ+vN76XIE9waQ
F/rulEnt8qyjoPzObCbMIT/kpfUEvDty7phYRv+WwTMAHaMzACHTVDvZ8w8sLgjaeCB990ZtXHgF
j4XKCexNaHG94SZfhUl/u9yH9HHjeaOthIchi+FVqax80XqQDpbpx4SQgf9F1s1/yoe8Funk9fBF
4rQyibWCXWVvVLtYvZ6CcmeAlxt85/OKlYBxjaVfLm8wdl7Wj4ALMCA5nUjI9zusyN2s+ZF7Oh//
nhMof8/FSDao4Ou5RtOJBsehYYYhnzBbstPZKtKlCyGFKGIGo5lgCOyMf1CYh6RmQChJBZxIBSAn
JAeHBx50sP1tnbo1tqhzPXI/1D0Uqkfp+kt3cMRmmkxfQjSG4RDobHc8RYU06pu4LY12u2uW6LOg
Y0DWLzKKoRhDC+bWc9ZMYXlet8tcD+uRgYWcet34XtlJ1hadPdu//4M3nWhrvOqAM3zdA8wIlvxd
p4glQlT2RHiXH22Z/wfJvKYjCYYTKR34HbZMH3D/VYeq6dyFy6Z2kLg4EieqF0NgLL2LUG0kfhjM
1Q0r8jR1Hq520rRmTQjJD0x5qp70xvX3gTpLrcbzq8s1MS4zpKbfHr2WlGrfNqr+B08ZPix0I1up
e10St8GbdYTGXYO4xmVtGrZLOynuCpAFoml/z2OH34hAd1YlXI3pXnB2bA3b15FUkM/LENr4OnPk
E01bShv31fKETo99tr6KdmHTFJjQouTGYMPzgDt4XGdTT/aHyHLmjo2f7NlQnTBXMj61BIhfQ4H1
KkWrZNifeIHZi789ejoNHxcXhHMPPmuTf8sCPhDd01QwKQWNJUCb89e4zU+6K9iAsfscIaIhcJXV
5vIOUZ3QlifizCHogy5xf2EX0HsnpmNM2jKzffQxUljSTWLNlj0VW3mP9t+d/Rwnw8FYNUGUVpIh
BsLGfdZRYVKdXz2V6iZubDXCnzKGfs0yv7kEgwIBpcs07RJ0WaTlWVgpfa7PKiVvUqUw7mJkpwq4
7IhYj47OcXnNcuJcObjd8sAYjx1IIAKEOIefKJTg6c/WMiOhz7NrXeGW5IEbdafhiAZnLkqCNxvZ
nwhwmU5hggIlcDLaaR5SdxcuPP3RDTJJmUKD0zGyJ31P2fLhr02QKf6sGVA2d6kycKps+mXeuCBf
Jvi/sD70KRdj7xWEwg2Sq9pzhDxrM/dSPGRQORLm9eJa4hdlvUV7nRBm+VgEFlk3d+5lKcM8VGwc
POkxqYY5um/NyHj9STGDIyDVaWmXN4McYYRA/magOjcbM1GFUbL3HIHcop9o2SD2SgqPnhGxldYc
eZf6bJUuKA3CEV9wYRSgFSUPD9rV80eV1J8EpoplsX7wbqZbZ6IBvzsQ/OWbE0lWUROQqFCPA7pR
oQQmC9UUnmLY9kXxjgFjDxgWZAXS4Oi1nXJAaFnkPtJLwxy288LTxmJburaYrJsI3YHJ199OKRqz
DRW9GBHhhRAS2OR7cQ9KxBfFJPVX1YWN27cFt+JIrGKIWRc+vdApoXQpECIEG5RrHQwpANdqa6Nm
eMvXIEswnkMLb7rF28X6Zzb4HZe8eZ0slWHYKvw+SLQs1AKRePsLERCx6K/26Jds00qOsR4TAmND
TkL/+KrmMqqxRmg3LlSwSrPIzq4SKloM84byygzi5aeAnFC+o0q856GK4th8GvX8BdEDJprE6SKl
m/Brb+Z88Suw2JsFhKEYF6Hloy7EzNZqIo53jR6tuhFWeiFSTAhgDWmVUX0y4HOI0q8d2oBnGb7k
k2FdQJg0Xk95z/HzT8GEdpKNWqIn9x0sYeOGjWFiN3KCAG2DleQyhgV5SK+h2RpxkrKxl+04Noax
NO9727+FjyUN6TSwTUlVY+qSVDAq1K7EvGp235dDsOYGkfSg6Pw3r32ru3q7zdKdV6p+Af/zEoy+
WwqqNRUt0NwmINdLwUvwCzuZRgP1T/RPWoVkUTYtJC2pxBBiEPLJtiTeEqmWeixFeGfkvzDgL9e+
OX/ytHgAJ2oRNEXWYVXnZGcy1I8L4kZkH2f8hUfM/8rD3Gp8URzrDfK4QfrphZmTtnD5EZ7gOd8T
24GwUPgyZk1l2bbeUhC6Vukmfim0JBloHhOgG24nLd/GGufKkTuwSDrGoKSXvokfnVG1jo/p5IHK
4u7W2PydqKHbQILXJYQVUV1F+C+pg8paylZgEjSnY6O4vfngYtrosaPyqC9Wg1SsOpZ9AI6n+McO
maDiDZoliK4IFgug+DPH20W4h3e6dWED6e9zzclvA2Nscx/kMW9HN6eV63fVGPd/jkxuZZnKPd2Z
9s/bAMaz6YfAythAPwE00SXJMrvtfmn0nmBXrOZaaJl8MBIpnQG1Geshru73P13I6V/OvjqW0N30
9Ch++HUc7nJTsWkwIKzJ9yU32p8BwspwBW5mG1m9MFApVxkxP8pKAQdhWag73kPSVye7PCmSNq8v
D6x9YbEdzruH/ewnBSzvIHd0t66WTkGCCHAobFHNPgngx4c6SiGyzEjSupql+jQZNyVUcQCt7jZb
CdmK15NnNVfLluBSjGO5oDEAIhszBGDOssZ4lLy112SPev8hg3Z8beuTcQhLnsz5hSWztuj83P0V
avsb2p1OYZPErEcsLuo84vI9ohP6GzX1OJcrMCj02qwVaQ8Fsh/hKFr18HFdctyxTucAiurMAfAG
R6O00XCs2s/DeRLx2CaNFctSQwd3ecJqJ4QoKp7EEKp2WZcqSM2RiFKilz2eV3w5i7IK64nnlGAW
M4IHezHeSxKc6/B/xuRwyyo5UfeAJHASiqPrW4KkKzio8V3NQkhfqg5EkbKuFHtG9RngIhTFFVKq
7NzSbg3TVDsVlg3y14/tbWc2i0GZGtJ0Bwc3+32qFOuVCNtGQRqdsvwv7AAioUNy6lvHI62gJJST
RuZ9/8aCkEKCZ7f/WvWuQL/6hi+SZzWUQ1sxiGC9q708eh1RnlfqnjWarPTBBgOitP1Y0b4D4Kj+
O0YZwGxi7T71JCi3QFOqyVyssitiiB/4qO7Sc+6h8OM3/sPktnugUEWSIUAlAKpEeoTU4lrVMV0B
D43MJ+DIbWIVknfkW8imNmE+pIjjcso5D5Snk8qBE/VVQ7aUsQCRaz7dmMBItrQ27m2nxXOTyCe4
r1LttWiT4daoV5BLpUetoAmFL3LCPwRhb02aZ3lGTXtnMJB2yzCKjvIZTeH6e9R4ml5yWRdQvZ7W
sBZo+BHL1VvS12RjaQr/cljfuIzV5P+RoUVdzkWkrPBlUxYSvqYty67lVJltfc8rcyTev5TwjtbL
bYjvPr9iQTqOzMWZF1hNUvSE2DipjTvxxOjzTyMjtqk3x1krWTXMvDzR689mRY5jj1KrLInkvDoC
qdjAPnPLJ7+IHaJ2/JKu5Uq7IHj1brN3QHPOdN6WziBm6BImeJuSvWyrjeMEnMF2/zWX61cnxC97
Nhaj81Dkuvw90oH9911OJ7pYG0Mn2d8erRDXwXohlpGrXFQ+yuNUA+TYijMrOov6cLU73kes7F9w
PxwZWto2tkgCBAN/yQakMfxrRNA1wVzaOhLiz37tfemLRzN3nVWcwEnM9SWepBberNjo8C/S6gWQ
lehPJOjs/rvoW/Qc5Q6fhezubyxYnnCAv6W8Adyr0OALWO2mdGh37apfYp2qkhBKNIkQ2q+A2/Vb
cwAaQRBJE2bgj8e6ZXkvpxJMMiT7hzQleHt69r0TEox6tAb6tZFYF7PC9ZN4jiF9uGaeES+Qpl9W
rGBL+mSvUSC8gkFRCp0xd/fBCWKPkDB6hqK91ff4o1P907ZXPzp0ugEqmzK4oMtrFYcOZj0iwh6H
D4bYmG0jQ5lWIHnhXXJBEbYpFJKgf7RSTJmA4IeI8Srp5XpT0T47gXddZ4e3M8aHAvcfwW8apJI+
ojCJWAaXlQgqDUqgJXMbwWOwwK2Mk0li0pGtXUKWiBHteU87fsQ3Y/25DneglUMl8ttSHucpoGwV
iy3uUFs931d2AmPD/pduPKv/GRUo34UZQrgh4dcCDZQ2s02nqer2BCooCVzOe5S1F/hMiVkr7RDc
XeLIIiOrQqVHAGA6N0lcqrwBW3gYvW55+BMjARovEpP4HVObBc0vg9CsvM3KLbY4sZcVp8gUEmPX
cJ+4RjD0W4Rp2dj1VkNxNeYfsIU2Ic3kTJmWJqjDYEfN583UihQuvpEBPxozXDX/TaIqbOvB3guq
fiBj+e8Bc8lvkss3TgmNXev52Zu+7YHwLTUcJAxd/aos0m5ALNc3sz37F2zOrUMxcTNy8ICxn2V6
LaaS3AU6OCiX5Z2M50L3oECP/zyuMindKwP0qrXgeGw6qAOA1sHA8s4rs+QS/qaUOgDnYmqXahYP
WeZyuywqS/rvvmP+RHc6XRPFCp6+ovmdoaMoJUVgFbY9iVN+kwFpZwdUnl+2MfV9j/zpqcsONSrh
h1n1X7k8v3qkpJEd8O+PIzWGma8UJdjEjdp7um1SNIctaCdXh46OSwAcgPDcM/02S2s1SoHO5PfN
iF3prALJ8snDIWFPEDsSqzSeqwM4cZPo999EG+R3av1BmmSSwNzK9WRTPSK4pBTmrFZ+UtS7kje/
fQWXUzNajP2x1VAdZJL/CdN1sIuvL76emFZvt57TGn7bzSh9vJ3doIKSaHyjOUaJGEJmVcxn7s4y
iHDVWZ1P/sPVhixr2K40pohCW1rr9WR98ZLyONWnI+tbo+R/3JdxFAYGrRAoXDlRXxJ8Of+JD61T
GjwXUzsn13MSnA4JTnsanZdItbOhq/sv6t8eAoJWUQNyIkRZsYhwgn84r5xs9DO1ZFY60tWawMUs
fxUzwHA8C0JVmVnvs70ePzBzf1jt0TwjW4zEypb6gYXjae6X7Zdq2UMF0fbO2D9M5vzseQGTDEC2
0scX55f5laOcaBA3NzdASnzrR593WQhGXtg0HVZ60X1KcdbxaC+B8chTeZbJ+fbz9cLa+JEdjT0l
f8krXYxWIWYHz1VWmM1dNV20VJ0u2PQSquBa/8U5zVNQIt4X7YjUoXeSFsynidh4KUT6KTy31tG5
HKMUUH7x9HOEBfUX3V9D3oLLPNJRiBDMAyqyYaE+/1Qzsb8c03fpHhRWXze5azgx6J23MxJDSgfJ
Qx+OvyEmt6Cqnr3yZBCXU8ymIgZ/uVRWamuJU2iQYcSrUTzV6VyEzlJvrIwuv/lk4XRed+EZwi7K
6s/UwEYmalFxTyMuwSQwqO5w4jsZhmR9JsgsEVmJG6DpLffXtglQlm8rTEGr46PSSVdvHZ9FpgAQ
h8Tu7EaAlwMJty8o+wFBY+qbLLM9Hsu4Qdfzlq5o6g3JxYr3XgQhHSGmwxj18N/CP/HGiq1jYHs1
Qoumn3Dlp4tkTT59ppFHfD2UKsF72awYX/sDeo0P/NOQQQZ63LB3wYrPzrucWqgPQMpAMEfbNxN0
VkbWcst1DHk7CPrqfNeYGRfY7cpDw9nXMS68H6Q12et8XH3Qu1fZ0PQEGI/EW7257/psFR1q6IGb
qQLd56REsGzbmb8y9nGyzivOvuzv/LFN4M4aE7PQDeE1iSG8vqqA0xv2L6DziITgwjqBnwjtcTCr
mHg2It7ohXTd6w3vlAiRGzaueK6pW6RJkZXfXot8fiUboOakq4TJKY38bTPxWog2gpPLqHdNtbQI
Tu37hfELnn4k64CDMWZgEfcdwuCmRlGJ536Xc2D0vxQ08mb26HcJn8w2jzN+rJlPPAAdD55DQkSj
eKl/B8KuhpAGC1Y8MkOreZ4MhN89LYyDf2Ndy7CUDtsJ/IDayTb5tKwUwxKP3xonx3Ep5sxESEkV
U9/GGfMH5b+tykcpjWUP1i8zSr0rfxs/Ax89snTrAtHQZlnUXGG9wl0z3p4VYpX1lh6zZyfx7tCs
0Q3RUyI5ET0UyahDq8ITKzy1D7t0f2KXCOnqBcxAljJVFQcJslqdFXrG5Xjo9l+IYMJ9q4Om/Z/p
PMSeo9+kt6wsbrMT16UlPMheC3BrS7tDa1u+dBfAFPiXrsqiiCpTImUx4Wb99u0jBFqPNhN3LbFU
CuQWGfD5TiVjnrDIf5vDfWMlkio6uPyamzmDB5GAWBOy68v0p8S4l1AJ9zXthiZCjdDHStCSKLIv
9Vlw2SWs8pi7mINctpyhKAfHYfDl6KeMAMj58XhCyXM1gwsVHz+Jnb4EPfWFeEKPtMBQe+M4l+60
OMUGbfo2FvILf+ENRTOXI0tBNHFUO9ltuogH4PfwCazkMCiwks33rqkxv8RIR9sqX8HXdWWsTX+r
t3kah4yE5gHtGiMNh9fHafHqUuaGsx6epeT5C1T56iOBZO3zZlKIC/rbhhR3ySPrnjQI3XV0UO59
+iacDb7wcr1G8MC2N29FcQYA+dFf2rLRQE3Y2kd85hHNwu6kAZRI9WbiBQX2mmg/LWgBxCXtcofk
1ME3uTB2RwuSwlQodDGs4eKqjoHG/chC05fyK8fkKwQk0y2t94aez0UzjmNdmVUjJrjb6nGXEYwP
EIw3+VA7I5fmW4N7guinNVBUJWt+Z7rtU7lnIK3lGtwxdibFI2pQAbuFJx6rT0uhiYFyMf6UfJ+c
hcht6gsitX/ieTUvCT4yMaB6ateEPn/CKaxHW5K7rSdEukjrqQ8f1EPFDUAk2XBgVUksE7pmJKVO
QsZ1afHRF+AIBeNd4Ylz76AMS/zLFwJTWrxSbkkDoMsst/y8ROrior/VAiKBo2Bv+Xee99wVJaV/
ObymYZBh0SBekYNBXjmCTRxKodxJgThX+7ppBCA4CSo1TKhqDd660RXK+NJTJBTzSRXzXEvbuxNL
325VRerep3++cqHy0ggyMoPINLVE02bBbpxAS9mhthKk03d1ccbno50lhvehJj3fDSq0YJVMyHlS
c58LuKV/An1/Lzj3rqylG69+fcK8ahYbgGEg9exigN9DmBPw8bLTbbjwoncag6cOr6anrL3a8h8h
Oi02SABwch0BSlHTR3zDLf5WpbS+kSfS4Rmq0RRMuUqAyAJEnhL4JApDF7Hdb7Or+1ATTWA5KlYc
Z6993QxlBbOqNNUXC1+njpQhDaW+EyTQFyi97fftwYnyqHcb215CqD4sKsSI0grz33mx1oFruUbf
sdy5ZxHMPd406ity0eyqLZrc+2ulcCeIv49E7M+KbHRvtIHEVQf/BqBTQEFRBF8B1L8kojDHm11K
1yTj/YiELBESAEiPCq+vV4QpM+gojW4i2L9y1fG55cySLV8HniCXy8TKdVGe7kyc4KR7IwMxUAaM
dhxUr8xfX6a+x7yFOMo4rL6wErOeaprgOceSp9vda4JN2j5ATkgP0Q74e3swzsCCZmFYEJ+G7vhV
s8u4SBd9o9runFNWPFgiuTpbwgsOgDaO77GmMWLmYM34EG5B4PAAnEcA1PbCj97NpwazrfG3XC3e
QRrobuOUwMdwCO7aiXO3ixDej+POESp0gfu/bdis/3RAFXIRonLzAH/RJEXqRNnzzl9UHLgcFaPi
oO8+iTNCzGe7174iG1i7NxmHywOZUb2QZAcGFR6dLnBCrUfLjGzTRiNsmKbJ7q5MImW/A7zNtbvy
jGSeJCy1vxYl28oTefSdBayLIwDGEK/vwJy/krJN3KjJrjEdzLRST0AAcVq/rJFeH4hXS4oHcm+I
v2BUmNPkwZ9gliILDaw+13yLhpyAJzlO4brrUMSSpf1v38rWFHVBnir9eVJSBIz3xFBGYGf6q2SY
YPMxABtkjeHIYOwSe8SSh4a9qBaLt4srJTvPc8do3NoHzTjv6dfvUjY47TdF8olSZwD/WIpHv52n
qYBG6Xza7ExbOezLv/tJruAEoc8YTa6p0fq4e+P7dqpk9QvPpdMU1SI04APCuvTAUSP4qBVspIaG
wytLyeiLkGGc8YxSC1muiEDkpkozeZkuzBe6gnUxd2dBbYoIfua2xfwjxQFVj5XF0pTfKKLmgGcv
3uPO8pszOkqbaBeehHhNekSiYvi9jnFBRu6MmjztG9EJMlap5OfG/KxQS5aqSl2eM0bOfsQv65kt
ECk3Z/E8yHUFmHg/pmPJHgQIiSx54bb05ob+eZmUcxDvBRQPnp16XuHe/ARiXQ/m3GG3xnhr1dtK
UzOZ5rtdLG4aWNJMHH1J6zpVGf7LGMKYjNzO1dyldJRtMw/FU6OSluROEose9B0suNoYe4cRzaCc
voqmjcMVJAgxdIO1KfQtceNDDtj16ywuvCzGHEoTFWBrvozuNGWQcjGqsx8vVD4cCLFaR+ouwalw
JaAKaRCoKm1NapowxxQNUy3giFixaisVdLb2eYD9bJjsHEPen5ipmvvQOqCVlPAVeUT6ausQQdF8
FMqPD0S7vbpY/tQ0aXo9k9Od7Mgrj0DwfN6jjLe60mhzdAKqXV7DpoPKLOabHL0/KmCV2T1lVKOh
4+7FVS8CvVkDWxrcCVa1EnKc1rGfXbNro6gHJrToUpHipqZA74Ypny1dpIiWC/WLnHmNirjJaVx4
CtruQyeGAIFy095JFTAXCoHYRq1Gi6SwoKoD0OiNDm/Ytg1Dq8GoeqdfHzfdaeyE7FnDmQDJJlQj
9WESEsFGgCCspdUXxqsGErrtXcpwSZmJCvxDPhVd/GzhKRspAL5rnDqnFpQfouVHLrW/mXbARty+
yZAGsj/bQTwkg9hJExhWahydCX3Dyhxd8Yu4eWz8cu8pu/0+TqJ6RctYiM5vs8UEI2CnTIBf4iE/
f/5U8ikcCWzw9O36yddoLdN6ZmrsUuiatSHK11vPkq+iF957VLnzmqQotRUqDCILyzpSmG8xMmUF
m/a2TPQTpShKQ8yVDC7ZGNeBM+rDRu+nTorSEPctOFAPXqs68xS2dtPHxTe5tYTCXocp+0ZsAw+O
uo+Zjc06vVouQIs2A4v1jTNgUD+X+4X+oDx0gpTNryDi7uSNdChiHICQkdyzck5MxpmG7qpCM4MF
h+I1cf8Rr5icRb2cd52ucQmo1l3/VFuqbsxN8/PXdQs7ELnHMv64f6nweh+9mrC3xuwEqn7DZqU1
TSwCwSS/7ObDnbP5RcG5kB3LPEU/Zw4KOwLdaBMczHnmHDVTkNpu23yhiqYkaorY2h7h7EN9dO0u
gp6nz8101ayP21QFPYmolEeRxrHRr/ICSUdvvshPWF/ksEZiXmc1Wjqgflp8B+y9iWEdmL/vuqqJ
xceRblwut7ss0L1FCnxZnYnwuiS9mNAWBhsatpSQ1OEUjjG5/ib3e830rHKhvqNkZxpCVmZ6vqwe
jvmephzJg2IqrM0BcFZSrOTM/ZVvxUwjCTHzfoOH8VQnSU258kyOrJO/+Ojz6YwMfmQwk9sKiz60
w46AH2mwrIhfZAUOnQmGqDziTWfCC3Lmutp8vewiJJ4O9/ui8GuIRGmUBL/OjNoc1yFu26hbpnMJ
d4YP91sd4cjD+3M75N4lsOc21W6ZH2Iq2kY2EUbdjYkj/bbvz5wOJZxUdLaOZUdeA80cjZ3etjC3
UnjjNQcjuJFLd36UBaU4Rg+qHaZYGFwOmlSl5A3wpu2lVWBD9g/xXeJr8nZ0rDT33PoyzEcB1L4R
Jo44N9ygcdQNR+cS+azuL4ef5OaZi9A6GyEjLwjWgvkgowSzTvwZZ8IxUq9mdtM4zJ08UeFAUXsO
WzxJmbCB+48HmJ/nUhrX5yqcl39ShIq+iU340ip1T4wsNxOcdvYTLPPahpoB/W96GeOwTnHzd4kx
cdTygs8aJudZVRiw4zf6QWNeqmJ/fvCrceUBo1ANFYZMOh8Gk0TYSgdD0tsy1DGvw/Y3gVl+/l88
8HM2jCf024vuSCePauiIEzqSFRRj/E2liQ0/LRMtaOMbFv4cOoNoSy/NjsOJZSte5ktXZ0W0GbQa
3wlp/OY1C4D+tUZwQGMgP2ya3Npd4O4FUGucSXG36OVm+hK2I4mV/7LFFQqjs+rdvNOB8npZYM8D
g4jct2MJijzVs+tN8WKVv0UMvTbw83kV9V7iCvpT75skth7jWlQDJQ3IGaNF+gb4Wzvfz0y/DXel
i9nyCsPP/i5d+++9XBo4Z7/SCGxrOPsj4avnrXwWZRPVLAdWLo5m7KvmHeAwOSxrGe51ab8ziZa2
ginkFkJrkXXJg720ZGiCqfq2bpGUdJlrJXvIRS+dYhBrHvCDpFkq+DFzGacMd4Noaq8Jthyk1PGJ
eDeRvvkXGxZ/weUCyLHErfxPFkj7dy0gBg9v8q/lWnbs6H4ZbJHmSS5IL1/FshNSpY41mfd0t/uX
4hOUGrIcFVH0lvqk5s/iIUHYbEdD2afwej7rALrgblM+uBmCAloIAgmK8Zy/qwqgx7qCH7rwCcMM
6a9rUpZ2Uqxtxhc0RB2Vfhj+OGcFYY1WzlT0sj1ebyUXCJvPbzCRRUpnaikeMY+3Y6SvV8Y6Q689
Wm7mhRB+T/uMx08QHRzne5N3m3RXcKNzuFNM8pOiWYp/L7VKZHNCroiVoAk/SWJDzwQP+hEIEG2Z
oLI4tbigAOIhAj8K6gkV8qX2NfW9cCTzemBS3UfBjsDoeXpF8pgneyYcFTxdec/TwfeXyqX4+VA5
f5ddpeJVoTYM9dvhV7iLwPnUu+klZBWsboLp/U8aqc6AaTR68FS4Lf/SRIstzaRd4sb/40MiL12f
xD5tg1Rz1FZBdxSNvRZoTZ6CJfR2davcuiQvD1FBz/hwxskuk2QCGd0albH1D19ptVDvhsVcm++7
kCZZrdInni81Rj7fy4vVgipB3P59gjfIVLkVKXu+BcS+UJZieIv0/PQevx8VmnC0cQuJ3U1Ej8Hz
+4o8x+BOv1UsuEIry1gF1T6HMlVMxbxlOppocGkuYDRS1U6a/I+pGXlMud8ORU+bZGisW8PDwZY/
JF/Fz4wAB9kEmbOF2BPvOEKVphET6bgytxixMYxMNNTL/L3FBdHoLx6iaRwE5KyrKZ2Dd1eLv76i
qEB+gI56IdzM5kvKdc/W8+Adasjf9WrxilEhDppoaqvO9zbkrPiD2PeBKMbAoOJAQZV97fKuflYc
X3sHSrF07kwUitQnFn7y/exQ1J+toaxj6+PV9/AO7ap89S9Hn8BVJeJkGfeRwSaCrKw+SQvkD334
6itc3p4lE0EvbFTM6zMWtnnhXRyChBNUaluCE/bbORO0AjTixfU7ht0Kcfg52Qauj2tVm6sfd0Nz
dtOt0/T+o5cNiBjmY+v3jUZa+ULOBmgcae+3/Q6Mz4gI/TFbp/L9kJCYp03276xECRAK9KbOyOx6
GUQ1/ut788SHXUmNKC1y6rI7vqpWLg0j17CCgUyxaf3DRWR9yYvfUHgq3KV5iHL+jY8Q8Dk06eAM
G2lZlBtgcCCRMtN+qaeeOKCGfqB+lXJjgfg+E9AtQE1Xxk7okJ62c4jEwEoNVJorp6yS8rR7JGKO
+8OzFcqUSlHCxfpvRKSw6q7VLdQ+P8E+0lpzWHh277yH+LiGBoJk7smzUQTqactKMcijDa9F2KZL
MM//yU9q8FxDTn2s9qntjqrqbPw8UvM2wRDP/Wl/GPLV/RWOb4w/TINsVgFPsQpfE9YmLZVFpU55
CKZqRdRRp+7N57lcaKkvP1MXCu8sUcFA1Yc2RWfEyYb1gG3bn8eYh5HQ/knPnCt2gAm0L4Xv66qk
v7vu3Z9UvZjMkiU9/25qOgK9N8XeV5zf+t3pFMeUEYa8NTADDndz5gZB6uV0c6MUAvoez4HbtgsU
40EucaBJIYaHybM5T2IZbnSIvsnAe4Ax+q7ujkFIW+2oIPtiqRhhIEWnx5vk8H+JTU+4tVFL+z58
VMaDH2JwdnY50h1WQQqIGyQeE31S6ZohaUtmpMUTANwD+mQSe7gKkj3pvpVogjvShG+gVE7MdlVn
lW6rWp5+mnNoi/svTXd6OXWKazL0Xn1A3ByMYSMd8Co7Bz4qMdcr/AvpAef5ANSeF5SngkMkjJT8
1x3w5DGHlElPXdXfZzO24IQRd9xMKuoGyA4mr1cySpUnZh9vUn3uSYxGyHByEPbBbw8OmkBWwWId
HktHajAWb+mFczaphSpg94MbhyGChpQ2zxpNFlvFhPFW92p0yfU4N68m0WybaJiMuw5U0eZuM3Cb
8KqXl01ZgYH1algQ+cLtSEb0uCmsZWVCMb4s2Gcd0Fp1uu7i7/12Lywg1GSXeYYFbEMwYR0N2/c9
MmK3ER8i5VvKVZitEFsYTVelho/vcTHm5GwFn7yaSoZ8vVu/8DZOrz1AaGokSFbucTxA+Js8ZK9V
yvtrDZV89gOfVFE3amoKLJXzHshC4+zo8J+0nwePnnnp25JuNuxMqMPlAt/hwI5qCctfJ5h0bG/v
11Kj70OwUAHUTRSqt7hWrDYIgMFjXtd/BxQSld3asi7Cj0GkIFHZcLnUAvmVT8VCXxzWF5j8WDyF
AjjZYGnA29l4z6/08p76+IXgpk50CdLpdY/w6YhG9zVNmNUFM6xNj+x9GxF9M0wzRgoEQw5sfZHl
N7JVNNqOsiMokWfjvZWJY4pKWOw/goCOAHPJLfqBcQl+PbL4K0/Vz8DTwKX7QS5C81CbZA4kP14F
dUk4D0WmFcwx/6V9F6Mt2jngFNFG2A7hgGWns6FqblBeNFRj8u//uvkged7nQ7+++vZrF2O8nDbk
/jOzMX9UKQT8gi+tl5z9N+zmt1LpD6bXgCtw7YF+QZ0J96KGlMWorG1Gz5VGi5zvCizwoKWNIaCR
XQOW5FRvVnFiofHzUB2goaQdF1dlffOlA7f8zpzRt5ACuwLTWQ0FAMUcN/G2vrvJpMDTP+7OuiRL
jkKB6SL7ZtGneu+9A5Ys0rPeVXk3oBQBf8UXl2l6GYDVjHSNYQDowstEr/F7PTbRKvX/cdX4oEnN
KGDGyApvAU70seTNnx19v0XhmfGuOZTIBP8xDkcScAfuf6EYN7Vtsf5QfL773yYnAv5Dl3idmj26
oyEzIzNs/vDTdVYU3tJEQS+IlqgWiItvoXeqaTogtwh2EPi2FGmYgn6bQHh+TbRBqkpCPhGx+fGg
/3Cg4AYOJKTbXtB+j0fFQdR6nS6NB/plU+zBSblJHPMV3J9GZTkDjagQE4xeMs8BSLE8hEFmxejM
VWRiY5AyoF+Kjqj4PtWT9Z29c96Z3U/jPkWqqMn7G83c1tGsN8HkNtUS6YxDFS6JyJpMGr4hmqjR
nJgGaZfdXs43rNUEnL+OcVLCF/TwhFTXcOe+/LJbHL+s9CNsEnLFEG4nEmsfp06mmZV0d7cgKPMQ
U9uPsG2it/D4bUHMn83KP6mQz3gPx6bC1jwNJfafOSXm7qF6oVYLanfJClb5r0jHMbe7R2QdmjrR
L2yOKJG3q8UsHeC5BGR8QiNyaUkVA1ihIcETc4OAe+1p9YnElE+oQTWeBC87d3FRnZN/SJM6RWLq
EJtxww1KEFUo4LhDnH4Lv6ilSIuY4r2PUYLOeH1YXXMRv8fvwFZdP/TTWC8+vJO72JxO/2vqXo8U
4OjBb+/R/ITQpFWf9H9FyIDyPEr2tRBArrArrgL4FyCecMxKHSj2XlxUBU/8leetl/vPaW5L/Rgp
d7VChcw6tukCSSmvmhXVPu8qMZLq5I3sVqWYEzsoGHh7md9k1vCfq9rh//OZt62xULCgHum8jeEg
JUjDmKYdgRmwXZo0kQVbQxLgj0LAdcqYcJ+/lRP/5W0vhUL8qpy6fZuBt0k2n3rpMeTN2E06PVRw
opKQP2Ckt/tsDHWadbai/c8GIVNd/1XcSdmBtBHxA4OxsW2vYSWdJDRAs6FERlhFG97UNLiU87/I
AKosJcFHyuu5YMTGEo3simh+ARM2k5SMsjW0+T1nKI1QEzfbW8q3EYCOo8TtQE2e5RE0pGYK4aDH
qaWx6VrKaosBsGMJScniEgqmfoKTfgB8ERXU/liaa+g3gXflXeuiamIgx12Gt2lZgGOAfJW/d2/z
kvbkZb7lHGsCBKl+KGgyk7eM5w8h3LpJAuzL8CzEEnaouVbusidxIG9x6wtpOMm49ppNH9gHqb4k
jKt7uPT/CrQD2k/v0Ram97ImzpeFSJKyHjiPZv8tcu5Ts3M6XnqYgkDX8tfnQ1v3uZE8obT27TbV
O+mODnLivJ6ul7G61JgTB6c1RL7gaLdFwvnmaC0pmqao6eEXINzGdDZMdBjC7XXocpGmcxvIPTQ4
4UmLv07P8MKVLk86Etgm1YF/lIodJWauuMYE3rH6yLT2bBW1hkJaXGhaFgbOtnBfxX88x5Wrclbt
Llg/aR5KWrKG8T1aZWew7xrNXtq0G9UtsLu4a0RE1ulSqlyjwjXRhg1LSfoYghVEbgwH5a1417LM
p7txNzGBzfv5tlHdNms1aaies6jvDnPc8CJWZXLyNFNtAA9X32+jUXbQ9FbOLPHjxflNl8+ssC3M
XsVaEdT1N2EdYStXzb9tPdUnd1vtJw0ecF9bWqM390EwWNTUFT4Hbze/R6QcxqO+uZUkdL7S5kPz
vgHU+TaKmMbaewzpS/ynTD1EGTlWptf6SJJnsekXiskeQXAH2pPqwVYEH66CChXRAOlXTjU17cd4
YVRgiUj0iPQUHXCJ95dOvADUHyDcYwkUH5PqJq01SdkYYtjhhV1GNCvND+Xmn+Icfh0W4YAL2r/x
m3vRsAReQuwXDva+XdYD8KlJSIwfWjQi6G27fE4i5nKWm6TBMkY62bF18jWfM3vSL8eIeMhnTH5C
xFxSK3/ffZCJBMQemtRCuNyZvZ/RdP/vbOS0KNiVvx8SqGcnJzeQOtEzzf5WO75EmdrveL++xJvU
DwfYO9osNaTX77RMr3+++W5SqNZhrBzr9QVp4kdV+K0rPmuZoFJixHKznKtAYbTQ4OSATZm4mK9E
tPcIRlKRgy7XhQULtB2Xn8erVsHItzfIE5RYyTlVm2lT0Qa4uwk2vlpxDEULvVsddGBmh+I16y1E
Wcpyn4RIptN8ePrTuB2wp1vDu7nE9WXqT+QP2BNvkbOVsdnR2mUDmituscUwZFamGJTZlmbBgBbQ
lwiCwN0ho8m6z2JGWD/6q2vYMhIYnmq26LdTdG6LmarwLtp39WWVyAeCfJisk/kI9/QLzJvFJ0vu
MWFSfVDJlb2Bkxh47ChUSSX0/V9UC282QFmMNTAeU+C5yY3Wy86JSnDZqUSTFmb2A20OibwaIzTB
ikswGnx0hfEl8QhNt0KWyoblDSirpVPmfDNn69LNs1WRvHogqHe5/d02ZOCD1LKyQWf2QsyHYRCu
7icHsfuPhL0+pIGh1bZ8+addcmaJEmq6ycH4IvN/If9zdl7w+2WLL9ELnAJr5DtocwvOHSR0M1WX
wJKyxrihHHHj8SVZX83x4/F4XKMpg3Ys47QbwrgvTwdXHIEqMxA2OaymeA57kmImMphERgTH6F8h
WVHNLZxfoE70lrY02JWtGo5vru1DQcgzPLJ288pjNGFbpppdi5h/U2Rt4PSK1B9o2MmopubV0YGf
ZCixyRWZ6JqrmNqTzDWp6J779cZAHZMems4knkb7Y4qeAusDRsSMium3RohDIol+8wnGpw+J7hiw
C4G9nO2KBYL37amPYaD1c/Y9JqFVQI1y05B2fCj+ttzFM/CdZZZn6FuoBFgNpBdTuI8aB6HbcQEM
C8u13FgsqeYOXNjIHlmUlCCnnxAzt729jXGqpl4eWZBw3rJt0OV31HI4oh/K+DiL/E1MsOIljDJ5
1yj2/kUCfZE8pFSa2WVQqkbaRHor+zclrRJTY62ApuFqLTsYawrcJKADiY1VZT6xG2Kk2UKKfmDD
xVJNzrsmpUjJXpt798O8eDNY8JIPKIxGzskSeujVwhb2Rzz/IpvgBbZqdsXeGKoprkcVIqueSCo1
6lopYr1zG4DeoRlm2dYpdQ8lsYcxQubM7fPGjaEJXdhIDuFcFtCJvOnfVDa8nDbYGqcFdlvKTfdh
1jg5tX3DytIusOGRWX7nU9+eJH6mSKDi/TwsqIh3ryGGIwaMb09xj86DkRnpxLevu2XVltP4gjP1
h1m8NYzRh5qkxnJzeObT1AJPIgLzwtV37ZcpU2U8pqyxQs2PEhRmZH5R5n+KbNfK/fru0wIhaBSB
Rhd5JGpTjvloO6cW4pQfX+wdBHtvlGevRLppDTJt6Djq5rpoLxqZRWcn3qiDTW9lz5QolpFOc8zx
qs4HJ888v1IK53zY37vkCZQfEG3BYT3NebxaZbBjbq5aJBxFaLKLY442XQTisWi4jyobyql0KC1E
IrlZBtJ1pXIisH48gWbygVS7pwHHZrgony8kmv+d95MI6UtbO8Q86UjgsGzzpbQVtdiNLU0l2fdD
pMx0dSmMtifrOeeMvyU1mbHKrxnOjc50OAw9OtPsQjMMAayVd8SAuPRfFJKRVPhV00oEhw9pmv/C
mr5U9oFgjSiiyh6xouUh33nHtWdIblgATzzLj3asxfce0gcg6jr86xtcFMggBgOp2KqLc7ZAh50g
J6fl9dSaliI91nGgN1NOityVhljU12Voa+N2Ram6Lj5EoYonm7ejYOw/YrtuFk3aIRjzLlNUPV1v
p6FXkrorcqWWGGC5FCJxpSzqRkE21ZQMbodQudB74CviOCzCcTSsl/ue0ZMJ1o3NBxUU1Zb4SuYF
lsfxFezjJmtOmeTfSr+8zUox0pw8FGbcWYh8yxeZddQyNp7yUDH3f1aiAuM/W0MhT3NZQdV4G77c
Sn16jy3LZ4N051mrBzmvfcXItMy0uDZexibyvhcNTAtsvFTBSCP8LiGGuvsXQXUv8MtSDsWWVDjP
OiAwbJAPRunJk9JCrpTVZPTKf9J/PeGxpSWXdTaVfbGgJUkVc4sBQOaTl+i6pVmRuJ9wbmKzoPvr
x+fJUpc6Nkqp2ib+aYqQRgaE4S+R85YtL/rcuOtA0D2HnINkzC4F3iNa+pdq3fI2xCcWKHWgSQVj
C60DgGZf96rg3Hc2YEYCjAibXGodTu+vFpfn9NkMzBKPdx2daKh8ht8NG0Crl9FGwydxFUO//S8p
pFQCPoAwQEfx/3oIL0FizTVXRldAT0nWdrlIPdEDl3H9BzNfUcyxvdFbNXnhcDVLSBdFJJFIBJap
YF4xhDF064AeD/A+/lLYA6gR1Ip+0krwerdOiMoXQl6WwSvFK+lHchxqxSuH2NGUJYO78ju1eLKS
f96KTw5pIIATUBCNYer2DcQ6G7+3IahaHXwiv2sA0vtMfw4t1J8Alz+hbLEUAxneRyAOeIr8/2ns
rS7sIHHfISJHnraTMK3opJPZPnefvRZv7a/ZNLuYJawKptCY55RB/dJTpKcU9s6pSjFFoyDezrUp
Gv0/nb11mJoRAEWiygtmQgdDj9cV/RiwDYGG85JRRboF/G9bcS/EbIe0tvGLxqI9rKro6r0XEgHo
/xaOQQO7sEhDwR0Hja4R1Nbi9//3eonsZ9A9hfL8uEQQt205PRsm2rTSgcFIoSHQfGFMAeKWKUAZ
9HopIE4tZBcPR4I+HyByaGu0AdgY8nX/Lq61bq7iS6aXfSa9zShng+hi9XhTWbQExlYhOwDZOIlJ
1tN7kZz2d5hAUX3xFXD9v4qCF6IeXwWsn4ptjioMfpivD0gfomTL/bF5hLpOUs6YoKwXODqTDoTC
e9lSi1QDdSuOfc8su5XTWmOs6mZgiGbEBCdbM5/4SNT0tEA2LamZfNF3G5rLQsbjkQWYEBFZsk9M
C0/iT2u7HFB+mELcPxVxdniSTeQlrpbDag/czZ8mEEal85vYGF+tijrxxqwmM6oGc6lp2VZ3qfTX
nVJ3JzsgJy4RuYvbDTbIcjiOToVfsNRaPFgdNep079DKhAcOPkqu0ts4Se6DREMxbbj/Sf0UGXRb
vckh6PwpCmvy3jhdThWxvIidMdb6F6Qji0+Zpv7CSWnLmz2W3yZVLCjRDt/ynguVA+8e5npFtaQH
0oGP6PIDVPSwAAAi3ww0dXCjf16Oscf/XU2gShv9KhxbTvsnVdolVv/SrPpqeHeaaHMVrRt+Ybgs
yTbP5jLjdgSuDt4clP02H9rAyDY0UbvTSEIYyhBR+o2g10zkOxOXK1xBJLEHIlIOlUUHzhzfY2lF
3zpzf2l/I9OpZUosQVqfRzRSWhROjzcRKUYjYqwyrugbVXG+RMvoSmmLpldQxgmrlBM3C0RFtBZi
6E2We7pfY9lakaxDgCDQFabesNWJtL490MFcjcRx2GIZMpxPZ9E6hrngi8RtJIV8i1G2u7cPs1bX
biZwmxgIyYkXkmxjHi7eXZJ34Mos3q1W1vbbRh/9OL6iIICi6U3XP3fzZhWIXW6/yw1CNamrm5ja
GPs2ujZF3eQ9iUmuwU4+fvZDAIgQTGUEHyjEfjQPoUYkrDhbSiprIgvAivB5eePPeXx6pcEnWAvH
jt9WucDKAD61qmTHh+yCJXaAN+gSNY2G/BEiJtv3eNpxAXrACuscFMSzwN9yHfBqsRPdsKK7UQJQ
Ai3iskwT8sO0lxcnN9XiOm0orE4ePn1qB/q3xbD+Owd8u6WDGGYyV2sAIUiyObBM0dyRhXPAOT31
Ld3ThV28CqnSRUaB5Uig7/kX5PQDG/4YZx5PWlLPE9Zw+yXxM/AlByjNl3xftwmQDQisW9khqX8b
YNMleCInnz2PQb06dR0XcBUafQPej3BOT34GxlXkrt9gq5GRxcARPthLiQNhaocupF6dv2+icRHG
U4AYs2ZJf+dgvyZfZnBFILIWA9vRm10MtsTir/Yqon7VgHR6DPHRvJrEFm/tV5xKS6okFFXJGH2w
RapUxN5OqWslXzoCI1rNgYjFOMu7wRr2J4yJ+UYYe5podlTpdMHQm0UBy4tn7RhVW+0DP/DPFXlO
lblT6cG5Ruvicor0GjNlTab5DO6GQI9vRfx9fAIrNCyaqkrJj6ia5720+GuJ60r1ib+L4FftDegw
VfYDpiSgo8FZPnIwIRbI6+azdIuHGIawyt4SDFohGBRv1RzbUZ/ffN65TNH/3kUnb9C64mNXc6IG
WlOaw/vpOhUhe6aIfTQFzVwtCs3d4g4M+FrkCWjLGOJYGuHJaWsbDKbPZyvigGS8qX308pb04IrV
j4O30cDUP3nTXs37uoTWdJDJ4x7DiArfge+3wdERA+ZgNHuHvX9eBWokepoWqfo41K5y+5W41Mku
7oVldjJhstI38B+wOhzQOVsS5PlQPQ6jJx9s7tzupxIP9Mb1dc5be+M0vlU+4/U0m2jmDCrOZEzq
nrxZCrEfEMsBpx7s/CVWLN5560otr23tm4PZRnAnO1frHugZe+z7y+qVBjf7HtVtcjsLqqWA5yZz
Wb135D4z96PkNuuSeA0BI6IhxRRPmdKG7AyYJrrPAg5GrD9sIrZYhRxoBaxUuBVK6UfG56D5EFHf
iPgUbTaOQeYH0z6CUVqvB77yzwIcfgkPULp8g7SnHrwdYmZxE/Ei+mad9q6uO6rFBb2tmYCFRz30
Czln5/+DZTuHUYJGMVEGCn+jH41qOgcfBLPB62JtKfI/wLhiMijUz2Z6iPlhnwyuQukWmQQB8ARZ
CbgkHdrXKD+PpQu3R71cn+nTLLBc1shVi8wDG6AEdKN99E8NVf0wAyKbfrtmyQnQHn2BItW0WqW7
L4zxN59Wc1dXNjuEDVIOhDkRPe5lKuCK4y8Xby2QLZxyt+amGkL5IzsV67G1WORVeTd6kuwTm9mJ
zKwp6U618VKceaECOhZ80GFF/1KUDVR4R/FMUteefL08fLrEy12g+44GTiQ0qGw+gTQS6aEhhqvm
ZgociZNbkhLVwWPP+iEkVIX/O6ZsmRj+fQSYbvIxjKRtXqhYPPtnJ1jLBHeayba5friHxJbFXYvB
mQBtr4+wG6NrJJKbvS72Q1fuJk4GLOafdxro0HV4CPwkzih/Yd9IPZa6mRfuyCfM0n2l6vfC3yrv
nqWRXEjFYt8cwP+hOATu0lmPkdH3nFzxoFdv8KG0b+aCOqh2IZvJWdoXnszxJlVdIHyqiziNuYB6
KhxbcUXzThZvPcH2yT1a1M9xtbQOde3XXLZv2myRrmxDsIs5YEJSl4fj/Kn90wg68kl2zLZJRSNH
4Z9TDpsV8ZValPqMtDa0NKm8Qx+s+cxrmw7vK2JnFMHnUXv9tbciB7QkRSoCphBjQVMyL2TBL2Br
YAqOkX9fVSG1SK/xDZOhYjV7LMiBIJt6ebV5KfxS9y/p4CRzB0uXj6aFRjqpD8Mf9+0EMKGhf7qC
yJHAJRJmd45nMqrIJLUnSQv1qtib/x55WKAtSxqSee9KgZ0yKDwZ81CD5rQ53GHOUYTbaxy54scM
bmT5rMLVaqgvEuf59R2EA+Kh/aIpZl3vuOqGWdt3rFMH9yMyh4gZ/Q+w4ejU4EI9zeB3xd/5Swcp
kDMp5zZu00xaOd8VAMAahFEotEFPl0+zaMTk6IBXp0hYYzjuQuGVChfW8f64a0rqcj1pk0Xe9sJa
XpsdsellFxlBbwQGuLbxbIkP5XpRFmPEoo/TqVuqPFVqnfWfBogyJUQ0RWwL89QEFB5h/esIwupQ
DF7jqUdOvBmHKKj57qOj4Kx6uUjF2MGncYOYJXHgxoY25K6LBxGK51sLmj+m60xIuSCOnZhCAccA
le0ifhM6ckDD2jqejsZ09C6YMrLllctDLr4a4rFKGB0rVb4nHR2UrxSKwZU1FbWRr0GpznG46f+u
od4IK3TVE2oOgqKdYp8L8CyrRV/Lyew9EhyUIF8N0VKjZCUF061Z6vdVn5sbScbxj68J94Ph62GK
S/p5gkFlnmpp0JeQR07ioEd8550B3tum6wbcR9Fyr404Cfz0KT8NrjoWXfGOXatj1tTP7+62yO4Y
VnIfjR5WOjMDDw0jqd5wJDWTn5iSukyB/pdS7noLZB+57/hmwLFWH42Nc6jOv2UMWSP7mu7xgglM
rLNXkdkX6F4yL0BcT0mjJdo04rSv2eHfFWLhEnIfwUP8a9AM9DwpjxiKQ547B8OU1YxhDXQ1DBLo
TA4GAN8FxQKI1T4ziVZcPduiVSnyHT9D64gvMWJIweQbSmp+9AIe2wPBP2eyL+jxDJVCsf9lGjah
TYPHijEzR47ZUGdbBcYd1drn5chgr9H0veC37VgD0oKOZVTcNyxYM+UKGRqrj7BqeiaNH2qzMzlS
vuvc5tZ2/H3TmXE5BOZw2uTX+56FlfnyxMFOGWyCoyhoEfz8gH0yqdWX6VY8o4ZFpm4NPRIymtwg
XP1WP/JOo8Tq6gVmqrjdwNot2/o136WG0/n8OsTViGuG41LpoFavlo6V+tJdbOyqT3V/ciZr4hD5
CA80sUIjTzo4Ruxq8zIyhs0oXOSB/YeeTUYDT0BuYzAiXBPsHbQlpvZaN0qhXTRlk6L1BrTV0857
WBbyAnXkOnQb1KyTaWj090l9xsi9gnMK59lys+1k1anuOY59IThmTSw7U5QD+iKWOhQhIvLbwnsd
lM5tM8jE3ln/t6BDmVEWWTajVoFV5toGizRIyC/9X6rc0X+mce/VC5rNl6KD4zTZWIE+irS8wRtE
MTZlBxjQFB6W2MBs4RPqqLNeTLuKVlSDPHp54vRDzjQXpcb0NjwUceMyjSAA0AkO5w90YQ5myahW
WsfuPaIp1V6VkKdVaKiwloZ5m4tQ6g7a44EryM1W7rbgzzoT4t83sGyQOWPvVd3fFG4SFPtbrjvW
6dcynthucHYInXdljep7DD7G3o/mdl7+PfcjiGrH1+rV6iGCLuWhb4qqWI81GkO/OfwWB7J4/R/K
d7WGx1ke5eVv29mJFZk/O81IEyJXFUIZzfOwoHcdnPmW9PIguhTV2wwPKajtXGOkNu8DwmXkVQi2
5mV6azglJXGmSf9SREuVx0q1hLoSHdm/NqvDV7GxIIv2Lb6Yr+MxsVONuP5bvU/Z56xes/7aHUcz
fL2XVbARPEB6Q7kIpreh6fbz5mMD3sPrhmEeeYDR1GIbnw0+7Uh3bYhkeyNuZvNKsriaigSCl90R
1SCPrf7N1rv9pYRrpZjFZ8axcwe9JCPlYuLCYFhtKkeuMbCoMyn6nS+JPeyKxD9iIzsqvtGaBx2/
N8LmYQA28YkDxeQlO9kzLVWh0UbohulbPUBZecKqnnA0TPWCmsA+KbiUqA1HtJ1g2KKx2R5N+DkE
6r7vK5kFFsHj3FqYibj30EeD8lKI6QbYaFlZ7K4xHmDGmXBtsoBJkM9eJ/pJbkq+/hE64ev2JkzK
npFXgKibURLTuXELuJaj09cPMgLPpV1I4mxjSaJNR7MrhdXQbDZSGCNruPl5apm2oFwx1rtILxzE
arg+U3+UFwt39CMmWfvnMolTiArAddQEdh/hiAjRnRpZwqmJCKfBvIHumgsseVUKOmwL8OGm5egq
Mc7HT0cVjEb6XSolHb5bzloAYc2hUiJhsUnZZfRVJ2pxEveSbQMp/Rof98TD1Lp8wTM27OJAwJSM
hWKuQROisssAxewEWdEW7S5JvKPJrhT55vz6spkEyhq8ps3lP4WlWFn5qw5M17ac6m2nFryG2rwq
Ljf6hauqUT6GRMcfQ1FNPThg/UXWIAJhuHnR3Jw4RMe195TYrMd1+TpSzA3bAYWK/bIovFT/CuBB
w/4+lzvU1/duA+oMSafpOr51TxnSxS4bJzTGCm00UiwrJTGINQEQo/aHNKt1BuiiHOkkzDwW6mIJ
w1M2Zt2j0cXNEhFRTgDMRVOl//fWGxw0WOHj11d7e5pstk6JLh4y7CzZt2DP4J9HNDq8FUUIxL/+
EICH8fZL6d1O8AipA5hrKT0lSxybHVrMZ3+mPjOJB61ckPG0hiVvbgYSVA/GWwLmkT/+UmvyuE6E
olxa3ZP0MQ8qP8pxUdRjHPF9Iz+cgnfrtwPmXZGdpFgB9qOCL0eOZ2VnxPHu0znEehO/sLtgElUx
vUVxOfSDZeZnR25zMwFORJRsLVkDovFv3kErowh01S3Mex/w6Htuc4uzVfqV6c3pM7YxW6X59zZL
IQI2s70EicQoWN5z6HaCE8i/GV0nSzRzvjkEG3k7maVIKAtC0t9SLv9aIBXqZwjVOvW1GVzuQrn8
AVrps2TFy7MoSsZe26dVA6DPNfqLWC2w5LnmxmZMV74yH21FP2C0afhpVtCJAvgLTtEKAVqqxCLn
2ELjA5Yl10YGZDCoH8mhrlXJw60NKZqnnWU5cClgAb1vEkzwCwab3whohJIoBYBuFiR4jyYLI7qv
Mkoeku34rghukFoxV1yaXjsrbgwyB6pDL/8a1Q6i/G8lCnAZKrDE73YpDv8OEgbW54TWEcxbz9/z
1Wkp3faS+YDMH1UtANImN6nEimv5td8i1ySddigLVVT/tF5yw2TLdncYN+zhcHgGKa5ZNAtz1UIU
WzeGBdWg8pkVHnPNRmDt/VMxr2fM8IheYszEt6OPqCBOhVdRuqsos6WBSbNippqKVzyNO1n5Yq6S
vq/1IaigMNuRRASus3bmxOoeaEQCdfct6A7GuDnmrrV2ppna+/rg7UEA2T014ZnWxhh/IaTyZ8ek
CXAcwD9xITcgUtxsaBKPqteMi6i5t7nApYeKupSlB8NOFoNYkUYBIISJrj37nBOu3d0lJ0tWIJbv
1mZf5v9MM793oyf4HWRedE18tvNXaOg3V7aCAp4aJ352bVP3lfBaQNtcax4swn/rfktRWWBJFwK4
J6mPXVtIsY8dbYvOnCrM3o7srbIT04jdkX90R5o48D+urHgZwO2dFQgEHK74YD7WqiOlOeH4Gyrj
v+fc13UjuyBuCR9rsIVDB2qx9SQoIPjbHcFiBPZ9Jzm5EvYNXQ2TYvGyHTK1y8qOgjCyg9vXlFlf
/VzRHTErLzXyiq5KqOvSzEZWfkx/wsBeWzmvc+Jyg4Q4m51/aDOluq1QXaGZv+PJxM2R2fmvM5BA
IKtyuujLYP6xf05vFgITCo2TNEN/QxpLAluug/SvS3z4FBFa9wt5LjZ/0XjQegvlGtTxK+/kgyH0
2aNKxzJAkaYHky4HNwpHwyLSJnI7GBQt3xh/Kz1z/7ngUnbOrP5vpp84FTtVdJh4N7uF0frvL0wD
5o1aMSwqVsgjKlzCmYLBN72rZoOXbga3wtezdj+2WFYFbCHjNo9pEmZEQOjF4V8X4nWu4fr51yAW
gfV/30OdJ3frOnXWjo47sbfoP5+bQe7LSJB7Er4olx/sKT6aN82nfmd+FKp3Ukpd1y7Ul2nzJUh1
Bb8lenvS9BkoBGYOcIhoe5hnkcOkhGEMMm0YyYYBFCwVPuJOHPD2AVHZvDHsBvGNUzj84QNLYhvK
ROp6VBoE+Eb3IzKMcFzRwgOYIEWi0FEiBsPdJEbiPMBnA9OGpbw4m3a/2T5w2iUSiGec2xq8g94A
ZEm8OPonEPZu4rBjJpp6XWGK+KnK/DaZ5vlKUZ1delDG3p0ODpaTBYSfZMkF48/b73Sl/SQsgitk
nG2WerlzHOZjzy8CoK83D9IAt2FH13487odhcH1QAQQfNpR1OvYJ+0HVc0Jr37gEgbQ8NW5jPbE3
TVKFvfwDmwIjlEt2ecgJTRY1WKfDfbLDA4t35SFe0v8UCygxp8Z4vGUmLiN8hpQjGgEVUD82UhW4
1KGCyIfMEcijuo959I+zSJBf6GtmRi2Mqhe17GS9NSxms+tXYlG0vZ7BRnOKHSFp/0DS0ofLbKw7
9onbY2KHMStD6/GWZ0E5NLl04VfG+sKwq7iw2OJTWf0NxmpIdrbz+0gZ8WqFMHZk6qOIaw2Mmdn1
gIfRd6EgZ/Avj+dLLvLDTPjSKrSIz9k++2VtmSoGTgwknfiD+xrQYGGCSklYFL2dIeMu7skTGTOg
KoO1vVqt8RX9JQEOfs3SFNHlK6TDKB4BYGtkmIgOV+UkmwN2RfkShARk241e7qBjTrKwzC/7m3oF
V51N4otgefVEbQkvOaUSuT6w3ykFaeMxmILH6BKaPwRo6+izCWpqz56513kzx7NRDmEXxfIzvBaq
fQjnPtXRMYsF/94mUFah1S5QkMY5weJN4VLf4+hhAJntqJrIsA16qMPTQlxsC3ii7sE3J8huFcEi
qEdLreCuy3TI7vGtTwLuWYJhdgjTE7RiB3mcZCLHI0SX+yX9biZuzWMg70fFdLTfowYoV0mhInyK
iBfAFPC4xdk8IEWp1f7/GjMEGiSEq2aJcf0muqKNgQQpq0xS6eL3YXQnZUEgH69bD9ePUQb7eI9q
iuLiTGBCPdk30Df1BedlyOXebuuOO5Byv7GvrWCdNVeFvDhQxo6ZkwZ2Nh1MZ2kRsG4qsIKFLjsG
LFQ4N0NYE0DlPWQgIXvQVcOSfLptBPEgwOP/8Up1N9Bd96nsWB9y4/rk5u4f72ij2DOX8KLA1DZm
wdiNHPZsbjcj0vCZ1edGFV5Jzimwr3XL7Ck1OJw0Exx0NsW44Aye4K3GwPM8bTuGa6vKy2Bu1xF4
gQDAqzQSt7DmcvF1c5aXuC//avHggxlUjRmaB+U3TLPIGVs7UxwuaMJS/dBAn7D9az98RcJTowMw
XvaGjfLaT73CSefYpq70A00HpDU7THYbHJU6Zlj37dxPC2PNqHn/inYZ0/D3U/nfBgaVN61gkoam
F5l1DdNLf0CU1y1oRK4KjWsb7r088SEXdlCDYCD9em7nGPRwe6/b83AGx0/Bquk+zCgDK+ktHbbw
t0No4G8uA9uphdx2kuNS5sgM5Iz+qHUhuihTaOWmIZ++VwD0v4T4AX1DCsiIpHwkjwGpXngtYX+s
DEdZ/OrFXsaVdC8RFKu1D6tct7cFw852OkvX4HVwLn06sPl91OTjq8lhlgXSALNvUQU5vDUsUfUQ
JSZXZipwLSqbOfDE13PFBuzDAye8cYXeNyTnc4bUomNOJFR4YG3ve1e6TYvH8OfPoP8wD+71f4qV
BN4M1mdi+wzWy/218MOQCjF76jL2Hm5m6hByyDyt4GE123SFwfw0GxCD6Xy9luVSZKSOrWpccFKo
3Thm8gSqnbxh33L8yNr5BtRJ7E+RdZVPupFjt1bu0oBJeVOC7CcXanYut9h7fYobl5a0e4lQV9tF
SVGnddjQnNiGJwIY22qBLAsZhMH+RcRqn9DtuffKTCnl8/fAyR27JxQMjS1bVcpmG/wDMiyuIn7D
/EUIDtZwsujy9wbK0MP+ikMPnzSPo61TdICN9mmxplxEablB/hrPPEHp2tzveTSfBLXuUhAKTn7M
qnJYsRQ+en6uscC6g1WJUYQfdn8kA7gsiPCIy4UxOZ0Z5HyUjQy96de2CL3yq+9b9ThLxcxuTvtO
ak6uWy7TNBpxJYTbKiBMyoQ2BmI7xSOQHIhOy0P0ix6VzPeCoPC5LnbnAhi8hTwHSZPlvWXoCoyD
BFEayMoms5LOcRKsKoqf10dlO/5knUsG3FNygOQxkMetHxq3tFXgcS+VW0mJ/RyJ/fDwPBi5k7bm
1tyZwB6RXZRd+F/1FF0hZsXyLYQUMko3xEtOW2/bbFSyeJ29EaxL48EYx4bO3rFGygs39TEEk9N4
s2TjamqbEd7hYDwOgDL1LvajwxXrFhVVTaEIu4GZO0Q5ZuIADjV412UN08kuU3mgYrnKPfQv9L0T
HhiRE6zvTCfvggjfslm4CPJaj+X/5mT2+n/zfisypxJB87EjZ9na9ZS3fzTWYqW9L9GmqTXq5kQl
bc9BCWtNg+59kwG9ogm0O5dz/lKDOMqhf67+qnB1dzZBYciYBErY5+LLnkqsmcQK25hYY6duDiOK
Pr/zwUhia7TelS7310zth9Ol4g8HO3OCVwAVqnpDTL7VNGsg0frJGTbzmsnaYPLdFRKrKLDHPwz4
XTtO/sBBedNcfbxLrIhuquVF7l7yrFk6JMLqrRS6LnouKO4IHB9fkXupm/Ef7Z+jw6CIuinCoISb
eLvySSe638nf/lHGzaR5JTru1iM4OuoWnRUr5LzBdWYKlWo8yf9oxujmFBwOwvWq+tBCCo4tOBaj
RUAnDZnxLFkN2jB3NdpjcYQzhgivhJ5OMWj+KbIkbcvQbC28XNcw75YkT92m7Ii0GUMism3mcEIs
C5njkBJ0MI8WCO00qma54/igfEUtgqybJiKkx6O1PfQT9XE18K5uoICNjnO3Bnd2Lut+iQuMF2gi
sYmnywQD8b2vb0ZSP55BoTnUtEzHI1/eu8rsin8KAIuHpyfk6g82f/G0fWfuBP8Zj94K0H8BHRMU
IPG7FyVGetps3DRGkbe/z7O+zRrFHMi9pXdS7voEVfEW2FZ+jzNHpdfBmmywzbG/dcDTcw/Xs1UX
egF2CB7F89bFv3HxSLStS9owwaVpGckRqY8fohiP34kIAHzNcvoOQuZqD0pT4TYW4LhnM7/06ue8
n6BjIFGJqSgTPFNzJjN5BGSLlluDncWy9d2CegvwPZ36bXdCIg7ZAhPBxsZ+UnxtrvWcLcFryUKm
6R0I0LQj7wjW2xLDsn7cm6aF3l6g4TEEjcQ2y/gpyQVJ2jqivqP2o1QL72BTrkhx3ZjRu6UNObV+
qXJ/OK9NGM2X5w7gjdZ8dqQviYW7zqG244RCcKrKoLl+p7qBOyWJ+rZfx3HdBqKfZuVnSjiJkt1A
Q9QVx2mUh+3yFFBL30OGIGWdafOmQrJ1B0B/zqV5MyrWVJwzqFD4g0ipjsKTmZPmyabcW55gUW3n
1582bvA9OHSAwFN2OJbkZ4Md74tguUXDONJUrkQ/yUafJmAWzeuxoQuDt5ctKiM2HBAj04TOeHTj
wrkufszUJ1B19VDhdKDlCNtVCZW/aD4PuXYEsayXi/XFDDsuSv8XzJ1pDARKpznXpjCFyhthx6Ib
Slz99cDU77mFE6tSYCAw2cdRntPK8IThiETP4QNLRkxZPyjgBQ5N6eBWsantqqjNByKFsFAPOo+B
Jiu0RZdJJ2Q3rKv45adM5NBkFqd5cDRzouJP54uLJ+Iu3TCX5aEEdi56SlaRvx1ryR8R3yGG5ibv
3HWPmRxjTz7UNLU5kyjSqFlZP5cSNlZgNsz+3eKEtLF0ZWaIwWKFqUW/LHH+SsAurw2BoCxG7jQS
YIfnCXB365mbTubmjTSDJUndJJLNtUPpvXVkG7T7o9wy4LEYPqkls/PLXgL0KP7PFvHXkJ+87mAQ
UN977MIEXEAdhGXry52+zHpZW1QCF+jpfhmQH0ZL//WIAGQCSzeY9BdAO6qaKV1hMKpA2ACDfZs0
Pbg8A1UXllyU8G0SDH5HdgFLZVFQo+NvtwVWdTA83uhx7DswgalLOx8ZWKnL1Cv5D2o/8CEyh6dG
+MVSOoq+vohq9OvPrti+nTkxZ2jd90D7u/YPSuvleahhJqz5TZ4SIEcSDfq+R3TKWWaBN6MXoAUj
HPbjb27fRF8NxVlEx/Gyt4Y7fQl9DqVeCSj8zdZ1GHv0kAtuTYLaAPBNn3inO3X9S/iDbE6ET4nS
M37WqI6x3oQ5YEdlKwJyYjzHfCJZtAwkhD84Fd32UuKoYaoFEqwTytEumxWIKWlPcw1DlXotyw6y
BwDRRkXkTtet+NR0EmXRhX7KPeC8B1kB5Db4uFUj47llZb9RAeL3AVKgtQMsh/LRe3IkAiJTXIMo
//MW1OWXcBlclBtVxv6tAW2zMb4yX4nWrx4BGV5kixMU7v3qdMSk/5oV1TltcBQbjUa+LT5reXYl
5/u0GRbmR1RKHbRkDEdBD4HB+7y8YaKgETWo6Z+1mV/hXF/b6KKw4WBHLRierHdaAGIHopRWnIUy
ArxW7BW8nUPEkvRJHrFle4kSUb4VvhYQaR8mSZgeLw2mqy1C8cPg1lbNYuZCatYVJJlV/rRyhNoE
UBJNnDnqXvlG2VxGOw1IWlnDJ11+GEw7rgYACB1F9sMV26Q1rgQyYnG13Vz3ZTk3xAQ5VRNgksB1
LcaUWubIWttlLu3VBWXU/F4uNZhB79aqn0Og6bdDLy4q9vivaDPO5wjKx4Xtu8TjDFePPiuFXRpd
JFHavQ4/CtRexVq48h2fpMX5IZfVB3Est++zgKo6GPFJ4YEppVECpJu699TNFmoimWX61UfBRm4+
Tadsu+jSGaLmNP6mgMTlAp7o78CE/LUZ0FfYyASTHkYnptsHs+3BP1IN7IfPRhGUQ3SUKwH+IMTl
fBju/0+JPFfw9v09Vo+YGJqw5mwV8OUY+xG4SQVKDHCeaOJKAQZOZkw7SH6S27DuKWFqfj1pzOTk
TSLpzjDjsGA23obp/1Dnsoq+nQeHUZfcL4tk+0jH8WJykCJbUyFN1DfZuk6UzwSLColG/gQQQULm
n5EBMwXclkMMNUCY6h8PaUcUVBjSABIxCBmIeZIzDLQ/jVZIVPSsMZk9oDAE8/3pjQ+tqIrZg3Fa
dOSXcpNCH6KkLZ7UnumByHByzMjjIA8V6i3LnF5AHb0LHMnO8RFiZq1Ei77pUHu6jUWlOGGiH3Ue
lLJLrVBUianF5P375l6Bq+OsrxAV5bm2Eb2cKNRJe3fKCKcCnxANt0MCHo+WuVRB/3GvLwyTkUPA
E8YA2yl4yv17puBQhOM0GfQsuRThoe590jiAbvqzN4fb9/fxH6nH6nlZy7qUi4sAp3K4tHGSGkTz
11d/ODKrxraR/Um9TDBrYl4qrawBoD8MrNJR6gC7bHojhMYYoYb14Ir3NRclwcnihYDN5ScPiCcr
3R0xLLIje5oHZBaL+VQ7c6/QfBjA4Hlp3WiiqmmmM2bI5l8ksCBxl86a8mkVq8dKgTVUKiy5xO8q
P/9Kkz5/7NuYGwlFcVrEE6qdMqnwp/NYIOnKkDjkSYb1RnJOVZGTNO+bklfN389s/9guyjm2B+w7
rHtPtpRQyP0kPstRumEo1E1ZIcnqNnn3JqgTCw99aP94Lj6FlBQwePBuN+RGUcnzl/AlvM7zdYPm
fhsY2mqAb2eRMO2YWPMEKo5PzlnYZ7A2b4pt2+MNhJJWNru/Fudq2V3n1dNOlJOO3ptlzdpgEQlK
7VNZprhAP3QVwNuy3o1AbvWbV67Hj1qX7em4QBDWTEQg3hBLDiuqXi3OASrau8HGra3Nqnk8mT7q
mXJG+DDEKucCwuW+YEoDV00xhho0xGUO0kJfzDwF/z2nlmQ1hij1kEbPCgUX0PT/+uIeoBH5UPS0
5nc8tZ7H1qW6gc5qbSBnBIz9nKeVj1atHHB9qfh6DxnO6av9eIIUrOnR5k++oeTSKURJ76fHAE0E
ImLA9B4yA2grF4etuhUMRoMXBcN1QEePbke5CDQeCgjUVzXIUXRGXIj4EXu8KczxRxqjnn6lEqXE
QId2WWU2nAJc4n+CrU4fxqTlIV3LKjEdBVTg7iizlcJyutXudJ7YnLG26lspGiX3jLKJZVXqeqSu
NIsu8wMP0YKN48wZJ+uCzFf7rG12NrLGWrIdaZ+qX1YQWKeX5dIFBmGqnYpqqMD+kEWqY92oEulW
EfcmfEhwp+ciS6OS+rpNtF0ZHwLlIldTv8BJAYNBleWaSi7R1MKE6KJyt8V/Mh6jAmArtVIeHZsB
CSjq4YAgGoyKyTA=
`protect end_protected
