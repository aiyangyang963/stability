
module ddr_ads_contol (
	source,
	source_ena,
	source_clk);	

	output	[3:0]	source;
	input		source_ena;
	input		source_clk;
endmodule
