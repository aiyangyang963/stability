-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vx3wXRBN0btT/ZR8OgDJfR/HaTWJfxaaK/6ip79LT1NJ+3KrtFk/iYDxtdh1YV5hwLMC87uAij6g
4xLUglhTcPWjjsXMF2153yxfgxRevZTzrR02RZwIL9tiuDrv028cxW2MPCQ14C07k2IOZbsjkvN2
p/bs5p2sV3SXGoJUUmOWRYM7nymUPDIS6QLCMoTGS7CwGp9c4l8NKZBKYkPQycIMb2bS1AO2wQDb
tjm2cseKJLgV3pDIn3kSPJyHymJq7Fgqt3KO8GdEIoedHXIhq2S4oUeAtaq3Ik/4XkVbfiN4f8ib
4iyB0Xyq/WJSvJ6swwxcPh+sxeu/ozMnJT8GRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
uD9w1Ur93JFy+/k5w52tZ42OryT2KB2xxGulU0Dw0qij3wS7SMTHBr6mNaG15qdKy0MoTbH0ATBd
LNHv/TXis0+G3S5QgOAOvpy6ePf5BgtX/XIUb1TXFT0PFCcA/rTKv5I9DaTl5jDfjQGWNkHgJcs1
hBRCgQJKzk4Lj8lD3mmnvVgrJ6W7kOWJcF4pFtiqsHXq8RN5RHMBFNkTshPY8JlWAYsLdfVUddfP
rRLLrLTH7QFP0Za7LN7jIPkksRkh0yhnwQftqO3EuWIDmTKkXftvNafYFgIPOVDe7SxIUU5qBu4j
tEmU7M1XLneBCKj4GsEH9WSWMPegp9tVZZ2YczrDsVDnw1Rnr5kTP+/G0+uUZypF6b8Fc3TlIL2z
GxTxKowW3hgPz6R4diQ8guQ1Q5PnKxnAOm8hzQZzWluUV3XGpgdckBBFBu8jE+id3CCAEpvnoCCM
dk3zRoiYqmrVotvVXa6PLbrEnb5eJsTRqHE51nSfLQjRozPSd8wW5EP/B4JxeDY1PfB4BtnjNJRr
ZZ3zKjhiHiiuQaLSAow01FVpPyAN3gn01kWX7V+OFON3UfAHr6xpXC8hkgIGgZVU1tUPIvW/7x49
lspSpy5tWIPfbH7XFcazwqzrn11Yx4fKY3Iwlw3r8jnw3ZYpBvgfc07XkthD2goFwufUFXsz1wOg
S3Clb00HDVBc8Ig4s51iD9YCMcKZnp9Y26LoWh3ggLPezbw9eO2b3lri9llF3BX5CMWNfM0KeZci
j2J6tnuq60hdBHTie3Tvt288eunWSMecKDNWufb+kiHerky0kD/jQ6WB5rGKan1GJbXLWOAmM2bR
CDr+OOmLLu5TnDOGEtWEUEjVQIE+L/Ho/7wGWwvUcRDJxmLw2qZVKEjEcQ90MXryzi+VEF4TN9Xk
7LSrSbOvHuEU8QWEGNe/LVVQdqJJnmdUfOQ7S/52Z1r9NWvrSMaDn9IEjGbxPzuZ8x+fvX6coRB5
gSQJEPBYWaSao0+cP2c4iTASlGXkjfzlK8X2INnB/KTlUPl9s8wwRfT2VxqUvDq4bp6bLS3Kk8Mr
8DMEBxfwwibRluRBn/9Q7HRnsQkeT4M7yCHUTbih0VLM6vh6OnZfowTzvQFnqnTDrIGjq47RUP7A
q4tVmsUpFinogev7BYyVUspbTUFgnbGV+uQpfilsYnmdRAmnfrm8P3W2IAfyINAeiqxBKGYbMFVR
k+hvxRhuZ01fi0oZ/Lzf+tG0B6XlMZ7NRzg8W/0BhEVLaEb1x2e6ERwWsERgrSlD1VQa/X6t9zfm
2GWsLZpdJqyJdWv0S5s/jY49fBohl6FEih6pi8P3SbaXeQgrjntuOiW6VDxAl7dvZKN6s/gpI51g
xKWB/gmV2tTWgBVKuOFV7j7g7LS8whrzfRIAGuUwQWdJcb2UVR0pkgyh9tC/LZJ/0BnOw93ej7GM
GdBr/YCmdFwfJAQQl1jT9zpaFiLkbiqV2i96iOVtHspHo48RljWfq+F/PaIY9zIFxc5OsekF/QJl
VKwHKZFuzIdJIFYoRu1/9rlcXcJq1/JtA4xjdjRvFOGkB+GB0HBhWFQ0EAx38zkor9TQzaacgQjs
aAEGYUCHbxWu0jNZ4D/8miP9eUy2VCWefNgPxzEW1w2lAQ4I5qa9s8aMeDZY3k4w3JaBwNgSFQGx
5kgsj6+6uRLUAThauL0Tr3F9HERXJfskYaeRva/hkiVlxoU0ptsTPW6s37CBXchIwFqcSVX8b+6W
1ncEUs0gmMLCfgrf9mprNZumHCqXIc/8f5xwMd9+8CGlA3wBCS71Gyljd5zT2/fT4ooT+kNrBJnh
dDnQv8gmXWdYstA//bvl8FZIgFFSHEdiELJiUBMs40obDZ3TL2LxBUTV2xW2jRKZ68dEqleNuwoA
qepauFPyaQSpZGZlLkslD9rFQHTkZvyS9PeGQPbsJz1/u5yeyFijV5M+OHXGMLaVZTpsCQWb5Bdn
bmF96BmY+lXCtEfl2I7dGS3Ax3Wnp+ydQknSmhtVDLjmRPR4VD6CBgbnP1coTBp5dyyBPRERhVSe
MsV+zRcPCGBafVfG3/kQ+4gHobKbM0VS18As7POpqmIeFr1gRQUj6e7ZXP/qFEjJznPoLUhpUeA7
1Nd0sh0A3an1dDtfQkiAdkfo6M5+e60BX8Q4DPGjDcluNp+7tP2xphbJMBUm/7FVKLRCZGHi2HLT
Qxx+I4/RcVzvC5ueJzGEUMfWgq/gN8FyPW4DVKxhjfDY0sXopek7sUCEsWmbOWwhloBHSi8J8uPx
ol0LWfa9iQBYD0hraPPOLzj7NE1I2duDRy9lrdJda6w4lkw9cPhSOykOdcpGF2cokSZe3bF4XN7D
wO+rAGQT6ZaFm+7o2zgt1fu+5CSFPgbhDePics5Tzj1TwLNadffXtfw/gjkZN9ZKdCt7ythPxzU3
gJBXyjI/ACK8WwxFm+GMSYZJZiE+vyPd0UV8Y4jfq9msd7eWgvXn5zSoI+R8fhtdTcgLOQc/eCkq
EiBsmVJiU6ZBBaYlzIBpx/tcNvRdSGXrbnNjF/LEIQJSl5ZXD70fJkcG3mVqGFemwhJWfBc2RRdM
NL3FsKs3+2V0yKsNj2SUwUuuAXgIQ4COO45wR7lVIS8HUZTXyep2nph+aUVSqn1vPx3rzg8EUMJ3
yr16TnLOACNyW4FwrghF9X6+syHAQk+bGvjggAcTRrB6+B2U3kgnRgKVdNAyoUS7pyomJkPgBYqL
FP/GANhHvXfRcBQkqnKj2eZAyHqY/e5bpM+3LKqQ52GzUHUquVuE9iT+WKJ73haDm3I29yoPgMoX
tNob6g99e4EbzD4QCrhG90BKn0St55gr4VOHNC9bcSk319V60+p9Ta8KJmycxafy0TCQsaQaBkgl
QerGlfIRGmGvsWjxCETJu0FTZkc7UrvYdiC/aD+P/ymnzoMnvL0PpylN5ACT9PvmfLa5oQ9R7GSY
DcAlZu3KWULfIwC4rjxbpMhlWR+s3qAnFULX4+9qOHx36qgg9tJIeOZlX8kF4eN7D7NONmbffWhH
WtkWoiSFAjXwCEM1SZnuc0lrt8V9VWuka9u3jt6YhEDtBjER00On9/tGFUyEdg9FLbPMOhsMdzCn
/dzV507gJsN1H5umkXs3wHI7pr5cUkMBBCJXE5XIgwfkShmPzq2LU6RKV32tRJx8CGWtqQLUpRmr
nRPd2xqpyXY4FjGolM9QfjBGKrlHoQByrKXiGXOCn/HQ/hA/Hfvs5soY2FdIrPKMEx0pV759gKZ8
owTskfjUkbtgSqSJ9hK++sTAVR4wNjEyUacEYROQnQrTBrocvBBHvImXY5D2sTlUgTq+X+atgAL1
GlxkH78YB0AGwClZdekpZ5S5yZAEn+CxfX2Pm61Ylwdul5PvJSPHP16xlEGtMCaH1nA0hn+UXciK
QVLTozIoA7FbjVoyW7gmNfrpu1Y3DqYETOdxunT10dbfM23P5YK+NOjr6qUZQUxUuAEegsBmCQsh
+bYDzT6JPFO4+IFEjZU6I8jvI4Tf1iZeUP9A/+L7L299liO1TDCI89b7Z4cM8kMagpMpA0xxtL34
dGNYzB+N3jMXaPhiNd4/dtXTCd3fz6uVO9GZQWrNK5d28MJZ16GXK817/y7U+kkJLP4OgEa6dyq7
JkgTzZcEhRReYVVKZDCekbSdami7H4Aa5z56PoFoSHeKtd+Qh9ucA1rE0hh6OevmiyGVIMxxiMJK
l50+aD8CJH/7TP0XHybpaJvxHJBTQTEqaOlL9CDZNoQZ2M37/yv0+a6LeFIWBvqpz9l+b32CVUm+
v4siBtPQxEHTqVNHvXbGpg5kFD6GZsRXbi4aop/wYmU9s3YHVmmNjqp1T2kf29JXtAeuLneu3v6/
7X0Ci1XkvIYQv3lm3XAIkxulHy6fXeasUOx6NncQGKZsr/sCDSxMxWh2TkpyBgFTYE+GNbyf8kdj
3/fNq6c72nj/d3Y1hbRzDRcs47bSmbs0bqCoxxKP+3s6z5BZ1WipBESxskt0RMUBmMwPgAmg+nQr
7ZPp93uet0FItqdS1i0T0nb/b85KZcWWd+IP47Cg10HwS6doJ5vnvN1bOjWpeD2QvEc/VLEtGqGL
Hty+T4i7Js+EwmK5bk+WCq8SUAQpgsGSFVMqthWKWPES8RSJ0Vk7n8wGCREkhREfzCY7sZEHhnYg
Gxdn/ZHCFWD8c4VPQI/KAw4LuuCMu8vRrgI775/eeYaqyXEISOMtXj1neWTWye/6uaBwtsHNdwGM
It1c8OC+Od1hdoev0hHBXo+4T+OB5IBd68JgMGFj4Zuiaz3ykFPiytxoPto7dx7naz+AvM59dTWS
loBiB+54YHO527Uoudhmf+/S0gcqAdWVpDaDPUQC6LLojVPei+b1lFu6txalzoe37GryBp/CqByD
pFY6/9/bCeiJtG13wxNus5mb+z+pfqvK/HHmjh+UK0Z2ctZAF+odinYbobT7l3sgVS+tDt8O2R3m
iQxiWug2wzfACWEVCSWPaS1TWPnjVw/baR5521EQZlwUS8jFKSuTXOu2J7h+KlV2IoHMuXsjY74y
kQNBsptGaYPvdSMLnpXMpQ5HySmGL6+taKOWp4yJ3M9Vpz8mYCD6lCHZZHz8RBJWbzAUfimEsBBU
vGk25vvDMSJnnvZxwyKKgl4OIYeQ+VU0u0ELgiR6wwLoa5DHhXFDb8p3Go6UlozB8iTW7TJy0cRn
JU6xkZHqPyxym7lHFAC/+Nbw6DvuW31adiF5PODzj5UaJ3/N1X+3mUNhMBFkyubFFfj1YfLsGgNk
xYmRoMQxIk9DqmnvJPPbg9xeqOFT9dU0731zcfwm1UdMDM3H0C6QpO37mCxtZWAcIfEfEIHI4r3P
qloeKc//XYv7jLwOYjswzhFI1SmmdFkNzFz6wMPQUvREsqUnEZWN/IoNMN1Bh6j/l6vN+AT4tQth
iAPbJvJbyZBaCODCQXRI/RaVY410B6vUCk1Cvu0vZ5gUN9aehjHShYW7Af5PrdmY0C9SN7bEI4yj
nln5r2tvPCjBp4FpKukE9VYFHnEMUFdKqBi//reFx24asX5NyJPoqB1kHIY+BvWGQE4o3e5KamOU
XscQl5AvIInugQpagA2d+BSYMzswcobAx73x9McXxriD5GR4ZPUQsLNmUtdZMsvrOvrltoUaq3tO
xIeRnbec6E64HiUWzfDtoh0ZXCh8g+zAcxBDRC0toEC+R1B94LXqU9WfSMMJTnu4z304hQIt41nt
c9SaLpD39dpB5Gk4fD8dIYWQdTYeGiZg+nXL9CV5+0U5llRqsALabOu0dFe3ebgDHc9CjMu8wsYT
56JFXHCfqoIepEPHCY7qSVx03TkIVkbjsGO5n+NPq8GcbRssFr2CddtC4aTdP7pJ8clmW0QzbbXD
g3D+kfFON+D8BeXODKVNs5r7I8oiQtg3+148H/foB4dKF27qafS+FBaRg6xUV86tJ3GF096fn+xF
KR5UxowKBkduqxKKyEqdcOG81RdbCZW2jeXxZE1yaXITMfbkoPAWOUGbCDby/omLw6WA5XpuIgZV
FlwYrgTVjSCi+l0v0MY803ERIISgLl2hJdo6fP5L0WYtdyQzJUQ/+e2w60XrG91DCrIfBZ85b2VH
wLZzGKDfNtuGvGLe4ALFUC9p9IWWXZ5jWcq0E4cGqy+tBT0evZD5GKTM4PF16aWfLkqsb6a1Iy87
0HbZN3X/sEC2RTwbZo31y8AYmxJCuKUJsejlXOSN7byAuXmVIh9dWyHJ+p9w5r0ikcwWYEPm3oyE
OcvGBnX2YMYekAVr06aHuBD1r7KBbf6ElLC2D7BUswiJ6TF8vHmPqWICCL0Uqrt4Fp0dNqGI+7tJ
yxBRcBgZfo33tMlEIuZXKfBh+swwr32BmXj/PLhWpFZqxhtNuCV5x8yK8XRA68jBV2ZgGBJUC4OE
rQasbNjEG/i0Pj+wni69Juy39v20gFtUGja1Q+6P9gyWQnx9exDLT47Wvv1ch9Oc5HPyZks7j+6x
Gtsoq4gh/DOWahfcO/pm1Mx2+0XEyKdBJsz1mjPvwz1ZOZwpuPsnVvp8HwFHgwLpv3A5A3REBg10
kg8XsPJPCLtMRLL1VrU5HVYiefRXMR6iuyrGPCqAuNF3SdDr9JXIwePe3YO1BgRU4NUXOZEUPyBa
BlF1uijXrzarIic8frESemu8s+CBFzitWoQ5Q6VE8fuSLamnfW+Z6CpxCogCDY45kam+I310Bstn
R2ca4fXOcPpDFf9H6MwqqAD7J93qSeKwgtomUlpDxpkkHu/CyCTdLpgzc+erCD+JEjcBP22zhlqA
P0Ius63oy+J8sDdHZ0AMehlWZ46sGoPeQhYq1MHe07BPN5eDgOp17OoImx90GsPIUvtafdp5VMPd
5JMgNe4snWwXXgouOQmtxMz2TLkmF8Gkpa5vwVqhusfQ6Z33ykvNt85C57e+6kNogiHrHwx3eYnt
AVKn3rU7B7Sw2Orsson8lS43AL8VfPh7X0NX1zFbHzJp/gtKUfapTysyvoL54LSI+mGAskSZBlzP
ksLr13Fk+vtodnLXVA/FJZmvc+u9V3vHBNVFZJvHUD9C/4+UB+SyZdL3az0C7Xa1pxMUCtDTTJ6I
c8fS6nACCCkQWOY+Va0w8xBkFG4dYgxcKBFmpwgcIvPngpgYoG7agLAQ9AFV3knnKVROeL9Jgb+m
3Fy42XTkP2wBZIeCGHpCRvMDg/nhLwVTh6meZQKxvGfT7V6crFT8Jp4vYTJgrg7W2rHR0aacOxHC
vGsjFC3Q0rUTr+esEWzN6xV863PEzr3vyXAaEFrvkX8H+peBjWlZ6spJQ9MNF9tSqEiMB3pdRLWg
IlDiS7EAcy7XoiOz72F8eAPEPUxhTs28q/W/usprxLfsTBaheMfff0IMS16788Z0V4bXggcy9aVe
eb/CUg4ddxJiWhf2JD/lfxj6JhFn/rKdfIeULMNrkB2QkZrD0jmyepBm251Od72RPferGcMWvtgm
rcQsK01ZfhNVxhgQq3Ll+3kuy0GA63ki6sK9fzElxOg9p7Xz1+LPMkQDWxMwObW8Se8vtIgJbRMK
t8nICXqmPG32JQ8BPTCZcoGBIPGyDFOHknSxPd9rmloTuB0mhrhU7JTMbE1lbCKoOiyU+pa63cXF
OaagdCfWfw/LuAc+mXGcV/rxrw0DJh0ijXaVV2xL49uGPIyllT0EQ7uyAQazy1cXwZMYMioqtTAm
x+sfOOt2FeO/8ieknhh6JNNO/OoBHD1gFvqnMI8dOb/f5apz7jEdQdBPEvC8o0/0YjMXXbmWuoiI
O8A8IpOfoG/6nKjnVLEi34Fx9I8n5CPCE+O05HGE50g9qrc0MwNjtYMZ/naFOgQT4+MX1e4C3+TZ
G3npt3wZ66HU+ClX19P6pELMkE6zx7Q10ti/XlWslcd0xcj51B5z/2oPTQxqBSUrn/sdvcghfNdw
8d4l1enC4XJ0uIEkbcvw5AOYvvwHnlmkFQzYdVAsd92Z3lwfITwHoZyZNGtmHpENkBybUp1jjrLU
ogrwvWdHHMSORH6UxfIuNDE71i1r3UV3e4udDfELovjSfJnK5UeFGaJSTi/O0KCVOmrTa1nPUxRU
m4tPyjoufR39faQZc02U3oTLq7vWY+craAOE789oX+L6fckc9I7BtFWr/k0=
`protect end_protected
