-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i1AWJ/iroj4WVrKHrTzHrQf4yGKH6HCBrbrpv4oFKUzjwG+1NUm03Uoxa133yMMQS+R4P8lZJ199
40ZeZ4yGaasjFDojnjBVOlFPdJ6X1o1CxT84Scfq8RlReXTQKjhAa0CkqCAO6Ctj2x/h7ThkYWhb
+udOY2AC1YtDhHMiHMXNo9T7sSmZ3AVsaHL8J0F/xaSUOnqmK58kvFlC2ZMo4l0ypmdmn96POZwS
B3tYU/2y40G5FAd8cNWmP7NNt+O0RFg+fWG2JpJ6qXpPjKRyUxgjDeIW/JTF8TJqtTJ9e4+yOhPA
43CcWvVTp5NpNwoaeaw6RvLu/JxP2r5/KIB2mA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14544)
`protect data_block
ZZgMtM3lgfmKrh6EtiyVu5YzU4aI8rbEnxRTt+ecRufIajIjxneVy6iuWmJIjSvZJ11HXFsKXiEX
i8bepcG3N5/eaPLnzyuuNwpfyvMDqB6LZgwDYwwcz3okyLOGuk/32wcG0wSL3ludzP2sdRmyxKOq
oUyS5AesFQfc1U5CJYPhPFU29BzDsNyfgzqdvlUNytiYz5PPx+D3/3ue/zLR2dZ/PY1nz23S+/lx
cN4rf/8J084KvA+dC/w9v9EXu4Sv02wz2BAOSCkNJdtXjGMxBGmhfXPx83MVrVNqZ0CaG4zg2JhX
Lu7LlKgFdNcdwEZQcyKKr4QXJS1ajgT+Q8tVUwlQa1LS/r2596OJqWxN7FOJprfoqYZvM6OKF8au
LUOmAuY9GK8a2SKNP9GTgB4zTWUnNmB0pIlNghye5t8tFK5sdHkyO9KsGgVzp+Jz5ibGqMBJTgaf
/Zzlrgq+/gqAmAL7rg0IjfypsUyCevlUNQ3i3i6h54D9rofRNv+qJkbfolqo1Wk8GyaKaOJ+UZNc
ihCad+i9JPRNyLYY6Ma58lhxqTfN97SeIx7xnl59yviU+vr2fT54HGvd5DDaEDn1F/TtIYTB+YhG
XBGEpdnVbgLDbJtlNh4+X9XMHBlgSqt/e3ST/i2G4Ew0HWEBHM30GGM3OBrfPuk1K8tSFa7MUNjp
m38sIvhM+mxbr2I0LQV/YBBdIVl2plI3djMKDn7GV8d30bOmfc9jKj4y+G0cDOEg0yVhgb44tK1i
Lfxs7eKe5+8EHk2bYgthCd/ZH8hVzuOceLkK+a1mqYo3ZRAlMfMfTeivSevsgAmovinerV/JJeli
GIvcFDBA+ZFOdsm+Wrdf/sIHrjYtvbjjuMJ6lJx7dnYpE/KnYscoSp8afyJq8o0RpqH159VzUCHz
CC6DSSpmxjhM+4/pADAYIy3Efk7056ELB3ugez0ysNUs04DrkqTKBFIPi0STkMdd5nCB3fhrxb4D
7Rgw0rEQ//XiEkQ1MYc4v2soTdS8Qx85cRfqcfrEUMWPgPdK+wap3iyIp+tjVcpqgBwiUTyvCYXV
A6xKSIvH3so28IRB+ivVGDv97J5sChY7Ygw5Y9gxAJjOLjkb/hCtlNu2Q7McSy8Ocs+rPrXjX1u7
lYDQ9wyuRqKkv85ZGc+y+07M4gTFfJdazV02wg4fVC7+paniI/Jxy7NE4KpOCxpfOhXglkE+PpiS
Y5R/iHnH0kHmhKJ56U+MmUj30JhdzXIvcyZgLrZTah7H9cJsyBEsfz2MW/55SVxw1QSc0OkBBFSD
erEViapfj903gJ6QDShoNJI1kpvujVUV4YnniYCsMi6D/rEl3+5jNGVVXm4affKXHfSO/9Kc0uwP
7qHj/7pAWzphzKWZtFFvylsWy4fHk5bMSb1BHAcaOEqwgpOcXGXntxCty+p6Wi5JkcE2qnnsLfzJ
tw8QCUEsxXhDswVtEK8+dXt2Wz+RdvV9gbiuwJeHbM3USUxiI3JFmRs6sSnNIz3qAfreBL+bYdEF
Nr+A0/bJ6RI/qsA8vuah7bwiHJOqKOQbreKI5xoBPTNu/aFl64o+FA4VvUp4HX2cP/Vo+wAtB5U5
FL5k3OU56eDvKn+sXD9wnLjSL8xlSoOI+nrDpWj+adeCVw7RjPfEz86Bj+y5cd8BPoi/rAVirv61
PmggVs5WnBpi9oKkwkJWSh0PxgZnlPvceRZ678oEr8NzuNtwfpnIVV08e58z/jVA7m9o4wYgVvcu
fWbvbUcdd4RMn2ao5vPIXz3gDZNapfNFKX2fuk4PbCTrtl6h+hbNN6fWARA1tkyZa+rDlRcl7AG1
eghpkNZuUyGkr4nnifiq+NWyiNADO+UbdgkT40/44ej6Kh1wVVDVmETJiCtGDeWnGaEBOwHwn5O7
3lFXGfmahzUEWju5EkOXtPGizJ2FYVoI+ZyMGs+eeGBEjoY3pmSBHXwY4FljU7sSV56wOvDTK9Pa
mkiLD8FsvcXNSFWB9tzL63l+wG7LXQK9IKXNDOD7YqTj8HmLuqBnnT08tADa5CuX7z2/T7TSIhV5
egnqHSnNQdz4R7hYki6mSYEnlyTPFOD25mncZNk3iTqv1omk0WHbIewbr8pk5a8pFlXE6GW9nfe8
L+dXF1Wpg4LmbSaEYKQlm2/LWFm6+bRFf1eS/CSm+tfn7RcsTcPr/+spolyfSBsfer6R8wG2mQsx
1lAIJ1+MYf0xwhrn8+d/v7szxMIQdQaLmhBEEAK/a0jfq3TqifmH6EHcf2dz91PvefqzCP0waobu
So3EW4vMPU83dQ8hgcpH0+WTX/RBloWdIyvfE6ScUIWtjdJAJI2WGDLEiLUTunh/ljPhok+yZpRg
YjaKI+IoLKVUqtiGaf6HjZnwJf+FIuR9MOz70zAY1HFLuhznCQfr4JlT1y0iqQkyURBNI5Wvl8Lj
mmjKAS4jBbvYyk/n31Y0X6gqFFgxqb/saEyMWgdXo/IEg/KLQMgSbZ71kbcoRb+yPatgnralVHqL
aLFEspPspHSczC3YzM74JESq5t/B7PxtGVM+yiykbF27s4okebQhlq+b7wqjBD/Fsiea9zpYzxCc
eAIPwOA+ZsVicDeD4/ASeyXai+uqY0EIYL3auU341f/nZKaZpRfyOYP59a03jvMvIVoxkw9elSKH
2TQEjuOKy/D3BwdjYmdsVgh817jvlmVTIjO/SHGw5uHPyzfWNbMBai2ZKvvW1v0GwVUEMlj/di40
C2kZjugBJXFJfhydQ0kwTMZKvApGhdqmX9WgvBnZnLdnOLXHpS4rnA6PD+hQf0qlyuPQJXAv7fwR
5+54sET+jbu4rjleimMEIGlKj8dhMwme2eh6K7GCYDVa215waStslaK705DQh/YxK5i7ADNKXwHD
L5TIZATWIqkF48Fo4K/moz5dwcqo29QEydSrOnv2pxpwCM/Ej27Yo/I3uxt4JGMfT4VI3URfjLkT
2hu62mRzjFDgZfDwA9LG63UaBj55bZxO/gfLYQ2T7AUVL7ZdYRQh/gEVHEiK5nQbTTgHZyp/IAyL
tAC3nJF7C7hOeU0c1PtvEQ6+EISDsc2CwwUwx2sgnGIwsKHUp06IgOnkTEOxw+uy0v3gAM5c6c8n
ivsmNNKu89zE3nzvIZXEtTqubFZK2Ms79bcxcp77C9B65JL/OVEXSARJ9LlqjYgCay4zD+rEWKB9
YfRAN/gHGkqRNfZLkfCEQzeW1WiO7gwPCjq6FjAPRgiFxTnVdOeVkSFKYLVp6JULvk8lfyD0u/1M
vnq11j6G2/LYaNhwKK9VXmGaWg0n6npXi8IxsD6b4k4L/pshF9B1pCvk/PqLy0wT3LR00VKteaBT
n0BErZgSejQLudZrtaZ1r61xZQEismx46crknABhsphEzca+hdEHCZbFm2DFtm0TxTFwPPyQJsbT
JQn+ta8EDdXl1u6ASolMgtD6zq3S11jPUr5Bimqfw3k+BWcUvfFiBx9K5EszAJYBMJ3BgYpdlqdf
MamHwsXlyomu6AUMV5gA5HynEFtMXoZ4n8kg/zqKWvtyZXYHg8TWRfpdguK6npA46QBN7GHsocmg
8Ae6bss1y7xguo2e3ECZa8F5pcpUGQbgTMavZsLl34aqpDdlJMaQbVZ6jZwS5Fo8u5FCFFFz/XA4
vm/qM34ow74heOMqRaUPIf0ycFgwyg2NRq6/kqUMq/1M03VrWFWQpg1EKEcB3aZ39X/k7PfNXikf
x1eu7Qy/iLnjFlgURuy/IhlmrHXl+mGb6oRcZQKE3AmsyOksTjs+V7upO2NUrccinBH7MZtZA6IU
3z8G8BXBW/ODpvTtJES0OKoBb8xP89jkjEZR9pNtDeoGpiTkJ79Ps4W61iAz6X78N6WHGhUleJPD
jTMaYHPhSTV9dOi2/V58nXE9MvCBBdrIrcpsllflBOnFUqsNTKuEEWLJ2esYpFxKRh6l3z/QsKog
g4AoieXZYPhkWO4ltfzxgwcom673ehaobOz9lToOjBaXQbHEm6p6vkaUwQtygGqMftkg5bzJZbVp
vvBjDVJYCk6lLs0XwNdC63Br74HRULBEjzWpedjyhCmZv8zKpfZ4MuwTAajtSDOzE4P73xbl5n+K
ODNQlPftrI+u8B+K2w0HQ4vorp29yvHyoz8GxewbId7n1fZKl21aA5t1bSZa/VyIqlrFcLrgQh7P
em+IQPxNukLsW5G6clb4DQOZjeqDXlkJ6b1wNabyry3KIrKwg5MXPxQZRlWor5JzfRtTSDR9yarG
qACvlQJcz04VU4LJ0j5BgW5L/a+yQBYq4O/XW7OKoaMgLbLPG/jRTyFVwARkL6yNFBd7l32Usz/c
pFlo4ecaSTZef27tZJ+1n/f26KnIK0u8PlFDqol1a88kUbhSqFK5ky6fKLZGyyt3fw/texRYNYRd
CMna6f64hMnD69GikLu/2DYc0Ype8ZGs3SBX7/WQbYB4ox5yzD849S6GoqqhMzW0cSkxIWKxyAqk
Z/FZzxPsXWpvVG71KD8cLUQFxG1SerKIxjaxPhtOIUC2iB8wFfebO7R8fLzcclEMMlOV8NfoKk8x
lc/1n/sIQHQ/Jyr8IM+tR7pAbJFOpCK7/HgsUocvEHux0haAEoV16/35foRB7KlJRmCfSplKxB/i
MD2bqVNkIXuMGMiTMGqDZcsMlptyBfcop4gP9sYDCVRR04UNZGJ7h14GrwE8qGWv/0Gi/IcJxiz/
5cFaVwT3fMTUoFpgdVKDMhp3RBcRJEipv9Y4Imm63FfE1AVbWfRNmAxBYc+Q6aa6W1BEmWd9SDs7
uD4i/dquOE2F6z8X42UBIJmWtatkA9CGN2HuXkZXQl08G6CDdg0L4o4U5Q+uEGzOJMcIi8PVF/Pn
KiBDaDCKAwn8Jfyq36DWf99I3TiBsHG1+Xv8UmTj+Sd57jbVuvD/qBV5CHjIonAw4PHytD1NDBH9
6YvEQk0lCLBVrTUGo/rueDOCuGHSSoH7RbMQdaoqJYxtqFv5hzYRuEfwSbi+rCvhy+gABCZ7N2MY
lFHrImWOwKEeLffXjdDyeoXsnOr/ngiRIQFzfIEmWXGHzZGmJXYJyKGwJIrgnw8yeqqkQibM2BZp
/9YDl6eIvTVgh2fQ1dmI3rh6+bdS/vY8w4mKjIe7MXUU2idcPbBn5fztKlHJMg4vzY9KoEVTgDXV
BQJ66UQt68N0OrHti3GgucqIjvsxODQazzenrODTLGlEzrgztzVamRTKnUze9gGT9qCyYzNnig5t
FRoNx1tPHgWCijpIjBEKYAO/8SB1AF8Z+Mbk8G3pb7DptNleevaHzprPnO2s0Kw2O0RU0qXJnwKT
I/JEwsfNbVvjwBAbFTDhgnA8hRohbXnCz4EWB3c3/OUngyBSqXksLYMSd5LutoTIq/N5FP1JEBu/
GEmx6CX1k4ixXHe7L7OwNhZwrbbdpwGH0IV6UX3/qErFiL6DAcWyzZr3z04RkdqqTGwseHQnh17j
9yiXmFH55ji3SPrST8TH9YEqSznF58px2VBj7bLeH0SmPNuTQ8peCVT132iXV3+rBJLzzDJbk3Ts
HOFLtL4LA2GphOC+cfoFXUlZnanl39FLCfRSKzPYfm6OhgLgwSo/6iKPXixjlteK9D6L5Pr4IjND
adF54ss0zh82GcYzQpKO3f90h/N+LzKpjv1CETDMbthVLxFoWi5poloh7XEwQVqoV5mfpcEfCgmb
fsT/NpVpgUHWeCwhV1An5HLk/Yb8oB5iSgXfpyYHB+G9uNtHQQUSGGf3M1mf085hF7WgrE7WnQLv
VGTAfHj0b9xerHqhe1ITShjRpB8N0rfYkRzT2T2sW4zGAsQQO869o023c9P6YSCzDgCf5YG2hL/W
YCrqG5Dp3nfqJfFWVFxptyRkwtiqYMZjwGm4xUBY1U/XIZ2I/be6LwBaXiOhJYEw00jWfhVf/8Rj
yQmHIHZEFLbWBUT72Ja76mxfJKiwYw03TlYhSsMl5ZJoT7ZGW+7/+ktNWMAesJQyqHCemLZDsZW+
ADyTrfKzoECQkYsSb/S3Y6hlo1HBPW16F1MvdI7KHzvJQMYxCRnBr7WNEZokZ3EQyQgPA4HoCwyi
OS1ShWglk8O/0RXhtlSZSOqzMabHApoTfkZkAqlDKMACzPE6Uv4BI+03Qd+prynYPcI9mRcvNDyJ
wJ2Pgdn/f2GXzT++GKH7yfhbvwDUsWiF6yFj+jwOMmdc2fmeRCLqVYOHpJuUmPS3n+Zpu2roDvfR
8NRoyQ9EgyEBwbHGaGqWQ0btTyS4MteDZDjUgpWqMEve/DjslnDs7koXqT3gEY0T5QXCnszgWVBl
cgak9enNIDl2a4gUns6/bkfQEqDtX0FTFB15Vgq2FqVaP7GaenW6KiIC8ICE4p2nV0XnU+HIvDMk
QKHglsXUrm2OAS2LXP6Us7JXFF+6zJhX3oQT2fCYN3zv1v+oJmBhCWb7B2CfOQVYQDsr44xVsxb8
uL3oDo1T04sVAeJ7VH3MdZEJepoYr2Wp2yHC8/1Zyx8mXrmhaDH7MtxgqJ/sJtyVCxhx8l+QeczR
67D+VNn/dWSu4LUE5Qm8ERWBkvu9WCd0YiU1h0dwiRMBFZwGmeDpdp+pcEz4QmAjeOmHHaW492rl
ufx+3w+crhJ3/+CZpRfYzPKmcNE9dM4XI/ZBbAJUY07bdql2FrgLXAmi66Td8aLM3qpMru5e6YVk
N99+Dtkni4YmLes84u1DPm3mefsAxtGD3O3mpYudfZvlC/iDlegbRPtW9nt2rrMEXhep5NnLg3NT
p+OPsDUc5jGtPu61vgA4g+9SGsFj5Pq8hVFI3EQyXzlQnt68LdLHguiudXK7gtQ20QNLaCFPgQPF
1Kq6mv38Gm7POibyPX9T8fgixm3UiGgVDqEkylnVBHJah8JQkeGreOG6dBCglN8Yn9sua3oAZopo
NYp/hBVnySdOh6dbkNy+ripvpPCFO6eU1HUuFNPukQ0q7BEQZnGuEsVs1NzFb8YspY/fPOFWq53d
UQ54JcNJBSkxivWYLmG2EXhAP5Xd5ozeVqkDUmu5wy9MPMGW0P6lk940cy9Ou6oYBxXF7IjjnxXf
YENqYCvEkR+SgaydiV21JzMLhtA31aDhtkIZ2fd/b3BnI5reOM19C15v19x3M6m+355dMCCTDFlV
Wkr8DjpJkc1rpdX5GX/WIuDTeDBSFqzdC+1lxSAUzcwN6k0yGn0h7nbI0DpyqBbY/nOiDnSanLb0
3r9DMMgEYuXrD1AuE8tybV3ZGUBqdA2M0SuUwzjIvB8fVOROdaEhWbj916iIQ2t+nSoQjcN9QqKA
vdtHRd9Bdn8acfZUJGiTL6JpcnM5jYWjcF39rVXntk4yeQFBhLwIsuR7eoOwZn687AK5wVpgF4BG
VoFT2NS1ujRS8e9qn6z6Ufx2vkwBF3qfWzCiEPDhc/5AhsusgQbnnsXInkljere6CUwAdNajJ+pt
1wFl/5U2MYdaFjPPDBAFKozbL+W8y9EgwmPAhdtS5DPiG+i19a4iBCjMjTkGbZRFtSedZ9LRSvi/
tC1Pr07WQlrbJ3DZ+w10bybt5MmvrDpSRQcNmOhxa/N6gGzTKPO6ZNk9x0omcmisK5yJOGrKW9IO
w6OeJwTPL7vWzzEWq9he2P/bIr0PkXvCkZt/lKQh2j8ncsivaia/k2jeyOsOOlm6w4yonCxFsliv
odJCjsLs73/qJshu5re6tug9TXS0Vu5L/aSGEUuvGtuu0xnhaMxx77h2HgPMo8kng+dhWBY8vKuS
uBd7EuzkO6QmEBdfyFS5W0d2ZE3U6sh3lYi/EwxASmKWb2Z2ap36DC04iVnHbba9drVepDeR/R27
tOvB/GHBdKENAL+AFXBSgJGdI9WjZbmUv/5HFeHx3O3IexDSSqOuOmLeC5PEoBBLmTxZTo8/hdyq
hi81AHp3PdERXvb/DVyM8nC6ttGH6EnDKchEak3nK/sYMv800XKj4Rg/6SrGXnBuY31I+brdc7il
t59fozpbm4LuWTS2uE/8fGRgk6pVP8sQH6KpGzuJhP/pcQTbOGaau6ckeknW++BRXfx4zntnud5Z
2uU4eL3DNh+xfgCK7xQjenlJA5qg5U5rDu9O++ShhgndioY2WGRdw/7YoM43nWuts5SrdWr4wxNE
qtzJAMWWIntLA6pPPnNTBIrghb4G481/V0/MBbnYLDigdsSoyf367GsHTCCFJFDhplY7uJP2k1bv
o/2GNH/1RQ7uuWIdWsXseTaCb1DdkdXc3X+rfNh0WwsZxxiOtKmmzm53beDAm8GXscYmspFBcCRr
ym6v0D+mRusjPjnmjPctMDMd9LMUPg4x2sYepWy1cUn65SuFpRCPcc1B8Ghft51hByAHdhEfQRyx
yxMdGMU7Cl8AfzruoWiFKnW4moJKPk3+UpqjfLkP1iSFzFnF29qv5naQX/DRCR7UNy70vIiikdup
dZrCpLYbZMczIihHogcG7tKPmAaKuOTwMSSb0J3ozETnwQrBCelkYT9SSYDIjNgz/twDYgNl7lf8
vOGOvLMst5AgRnXMTpW4QLJeyD3Tz+tS5YEaRdmeAiYCz4aOlffzSYxo+mTHt54VXFO04vnGoDeP
4NttE9KYWYhcVChLYLUdyizr3KvSxPPmFvQkMLaNI+pQJwGWM8X021FggSeYiCbhrqKgZ24OWqYS
UCqu5rmZDNbGXAu2dcemWRtqBaXIVUlrky6uL81N+lI1qsM9PfeZqnCZAM/URyueiTCGagMPZGuC
e9z3x03a2FEIngMu+67OU4C7TzDjbLZyX0MX+u1SWBSj/NW1bRpRF1lnXlStpeuAubymFC5pGosl
LS45VrfOSqMr9p/FLxMkawaeBOf53T84hainuv50QAfk/njlSwCCzpUUZiAPQ9h05NjkXMza2KWO
rR82pwb/7d2nsLx4Kl95V48/c4NuyN5ZxkeyGKp5a+P7wXztdFy+j5Gy44puP2+LBsXmve5jAQOk
nyy2m/5rESMLt0xFw/7OijD3Dy8j1Qo2q33P2WsJV47OIa2WZP32Cj3Wl6JsjR0M/cjpjz6NX00p
FjMLUgcL1OvMaX86zlTcmYg3Kxnm3y5e8oexb7dSHGHO3i75VhQemVJiyOAPFs65YhlFKGfKr2Th
a5Ptl+Stvs/7+fGAi12t9Y/SNyMhatUYUEjHmZ+ECfkZp1wvp8bd0Y/cvLLSP/yYADmNVpRhgrwn
THSg6Q5pXIjxfU9nb/+jPbjNpV0AGOo6LjBKKh+qqh27sE7BApDv692lRghgvwSbGMApmiZnimET
khBbi2iv8v5Ld5mLEadnL6cIDU3o4nR+xMlLocBEwdk3NOBV/1k5LaQEIn4h4D1g6BEQWzM5gTat
XGj5/hk8E4tBQHI/Jv0tbnTyTeMlaZ03zHVVJl+5x3gpTWs2l2/uLLNUGr8YS08omkWXJP/G7s0T
S8nv+E1qVUTfdspJNsxQsqCZXyG338fCWm4i4Ac3KP8cjNm95r1uDH0ffaL4xeyGNYe4EPmPyu/O
UtubA482rbZt2/tIqqdKRIq5dc+/KFbmyraVybsUqOzuqzMHWy+F5a7DOAQHJAvczNz6XmYxm7mz
j//sPAJuZA0mVkhE128bf5Q78umQ29qrBXX9BKy7rqWhU2AqjaVHqt51mMOOu+hxtU2zHh9taZb0
TuM5S+VfCay1E2cOmKcJ1urMZZy6njrKt15zuRXzd112RkDJ5bbmMDe/NpZ248NJwTXT8XndeVTG
Ln5zUzhpDoW4PPCjE7VeWXUld1Chly9JTCZXwgC7ixBQLbBLXsO7H34XEIkilPw0AGTTb6RQKvlu
4npuFKgtXzLRCS8dC56QI+UgL61RVXX9v2rx7AfyfEzYNYhvqLDIGGyatHchBhGzD2zv0/4OdWSc
/BFD9GRrnprdQiE66ItvvUPBasZGnpyRSn6OvIYusC+ATBXKLmKDC9QP8LPXbF25EYkXHsnNk9CY
3M/JTD55oQnDnZoml83GRyGyQunBAw/jTvZ9OT4hvERp6oVyY3fw1aF/VkHssc9erl3+I4CPkOd/
iorV4Bu68LQDpvn7ykHn736wQMfQAccJMWeknAGpoLae04XAh9pzBvSUU73DfPfXaUGscP6BMjuD
wcQkDGGUMcLMS4ltMmdQgRNpngfH+PIRum+0rTAxOGlOp950Z4tPzsX3nFkdYnqkKYOUXuzU6QCO
I1YXt8HInf1x9yaT0aZH4VXojx9T/1bgN9YYWML7KyZeSE+UoqaPgUcjqDfwAAOkaX72HOPQTqYm
7j53bKYVjCnyqqEOdkp3N301YheXjSTeA3cMtPqvcggccL3hAdq+zEYP5mFLU0S0G8/MdgV5Y2SY
wAUb3UmFM5pMujclGI4BVsIE7zbaE8DfelRzvhfsaMojF3EwqhJfLyPYJMnyxafF/GlyQzVIKlvC
MLort2i6YuVYv7knW7Qtkoc9v3whq8kKWaXepW/AseFH4BLrk94t/eJSt/eN1KPQw4NtVjuJnlOE
WzrW9HBOnLGt5rcKYwhHLOLaL7nwy+Lenu7qUtLNSeRCq7Flz1w9wV6cfZUWLlgovERXAFAZWuuh
oFvN4fHtRy6jeqyMw5jh7tplY4kKbZQhfwY0jRZ3Ov6WJ5roB4XLiKYUHe1Elal+yZV8xj5Gp1wH
6bhFRw8dAZa9c3ilx0vn7prA6utAY9ZwcXHgtyxV2wLSiiGdp22lCgbYZAt29moO9VfLrYlcQiX6
4RN9VePAlL6HviO7ASl6hGgIGWRCv+yQb25XZ3VxGvpgF5RaNOtWsJ2iAYAOjhfvvSH6gSoOXmKR
g2ROyw99PQlK6BZiLZSQt9YDLNUsfaX5CAj8EYthuYytMUwTwOxSYfWdD98V4mC7YJfrBNMxmhTd
x+3uO6U6soF4P5vEqyx4yRMQc4tBgH7dDUWAqPkcHJ7EyxU9E59G1q/+j5Tdaaj7WzCUOUmeFgcz
zIcxvYPi/QIrYNf8p/gqQx9+v5tJSS7FrIMyor4BVRdsI7pXyBzZj1GpRIgQ/p/+bmn//nGKQoD2
toHO68ltL5g52byCvNEUdNUj3Bsq3GnVsQbRxDxoO5vV12HGH8pRu9bQluNxjPzREU5vjsqvdcuI
aGbvz9ZyYEa7OryCUxZYCCuD8hGedjghEaDT1/7oVvx5f/+eFdWUEq2OQWTRR5Br5RSgXp6DNtOa
sdPI6o31meBsJt3Mlz2Ac097UZ0hG/d6bM6baEbqFIy4vZac5mlGDIm8cP2vTC+GKBKsSeGT8gYJ
SLLtii/cnDu3YuaqW7+sDqLzonTQphWrLfdtZO/N9bsHVn2z4OaYLZM0A5Si7uriCC/HI+UqeKjH
GTKzBX9Gtvs0r8FrVMvK/A9DTpQW6gB0VmoGLmSsA/K6jN+vEkIFpDkUeB+Db5d1F9aj4W+jiFGi
flEV+hP8fF+HWMp32iVy1lB4JE1BSPJ+uXlF7EJPWhJfCnOW/jTpgcZBA7j8eEB4hPKPFkpu0WCu
SKUJ/VpqupunEMHSOUuYfILQFHSdNam8ZgI6cl44e9vK4TdG+h8UzfbrxlFrwnWu7Bm1Gl913Mb9
oOd9YQ3vcqGIOqNub0sMi8A6NHow1k3ovEDY6+pFNEb2hYOogW9dp8WTZ2QadCk1gv5ZY3SvNO1V
7mE7byc69EdHheGrpx1E1KA5h/dKxF3UQk6vbC49aYrPOW+bCenL4OUdYoAS8UNHYPnJkei6+I9P
llIrOGaYeh8sa5SUbElp0t48H8b7XBWHlA7s52KXKTmhYfvBHphoTeLqYWX/JnvCNudWRLkP89BR
MO/yG7b6Tn7cBpvFHj3ht+oK3yYaoDFWkpC0mqQg8QwGaThv35+u4LrJuRxJpsbaYXAyCnWHobEO
2lD2PTe2B5jOCjtytFomqwprG7hurqwjADaDRZXSJoZerTskgBCarMVm15Wp1YHNzNwlMeI/8hp6
E9yXRAQfxznNbH7kLUV9GqnaCOmrdggYZ/FicbWmIQfg7JHKVRBM6rZ00EAuNBCrlIxB0icvZJEl
GXiQN2e2e7UBI6Hg7XOKz/w7BdUOfH4o1zMQVPbEnnHyxsonads/t83cjHEwxusnsStEt4zfgmc6
VvSmLJkPeHYMnZE+uipXcR4C8TY9wnAjnOcEqxEWgGgEIetvekdXRIlNnJBQJDvjUKAFUizduXp/
4lx29NEgA8t2F+Aggvp+8VHPhMaGVdLqTBQloWAK87QsL8d4BeXJhxG3BaelqGY+lOI50vMEkbzw
eVBzh3I820Zf1SDgYhVIy+e2M04jn/4zIOJAz33LkdXjWQP7MypTj5/PuxJK7EYNPPqWJWZPaD+/
N111FdlyHzAvsqeLImNf8c+sKyxu0Ol6gTgaouqV91fV7Jp5LbmamzLaVM63Q5Us2uvCiYz+SrSC
tdxkoaAELqO4Vt2eGnnfdo5n+NFiRzbZ3INJj4kMnsO1SOAtulUIc20kN4qWeuYrLZFHx1i63Rd6
3ZUreJ2jndVdAHyCzO+gN8cxaVNDNFE2wyTZUo7MUonJlq1r2X0rwSvOgtq+utw235B+tv84itAO
y1MOkcFc9fSAv2RU+wrDdF9ihuYImEj7W4TFG4c2D3GHf0k0M7U6GgZkWJ3DMfQnIf8EMQlgFoDE
yqIvzFRG6ITv3JJQVzynKrDzCLwyfCdU9/Kg7jJhUE7+vTzicLTGdA9pVF8Q4/rvoQcRmxD9FZkY
kZbKuxJ2s+utMG/T+NLhbNiR6j81U4DoQTz41oLQbsDWP2i32BwHNpztkkLfBCJuPNuhrgbwqTCe
/ZBlF8MF/ou+1D8FlPBSLrNHW6UokLODBRjrunXZ8qWsASxgxXYrKWbSTRyEdLQkzWzeDgYNLcrR
sY3g33GY6RGd2vxm4id+mKPpHyfWa6VSYMA69DwVE2fDPj6eFsiWA9TI92I/tgyo7MiU55NveljI
rDkooJWm+ERML0C48mW8PCUXTliM70snRDFglNFkg5Z/u+tm5/BOmxgclX7vavHAUczyoGD8ejav
A5UR5HRBi0p5AGYjWbu5RqlIkueN34tE/a+/Co3UTWlH5N/awNMqbA1L7MrRoF0zEQSa5fT1O1N/
nDrSTuRhFyQYVr2wbZuSo1OopZopygAh5cSPy1Xih6+R/iVzfswkzjO9Kz4yzp6nlGS5Br0XPsFC
uzbod6jmIPZci8mGkSr7518r71SnKpCWFcKr0+WQUnRD6SamU9nrBrQ0jpt8mwqiLqEB0DB0BSWs
lB0rUIIk/i6bxyMQqZe1MzQn13urZYrkRw6FQA3Sk69E0zYm/SZh7gY/ksOqLqxBRi/ePzr4wvgQ
mxXaln+vJmHyKQcG3yYF2reol3w5HGwE75aUf4cFFNGlDTCCDJKi/qodBaYeTyHpsyBnSUsg8Svf
tJei6dSZdClSNMqDEXS4Pjzs/ETAPdUWV1BjDtCk40ZJtalw0WRuR9nmVw4MRjNYShVkZYGDImvh
jEg5Krz2L53AI8AUyUy3fhySO8Y9SQGC7Vrn9/c5ve3xLlLOqMCkjP/h+W3hqGKoPg6DgPgP+idu
mu5cm6quzfsBs47F8XjJ/x1IO+pNgXzKuMdOTvged2fSwpdh7Ma5NF5jYTw/Efc0GFxhugFgJ6jd
5n8bDRYx4TtKBwVJziEEoXTey/8HWqwUlekbskNy56wmC/2d+LsSMy5Kon6PL3561WmRPXw1cUgy
+zpws6vO2NosmOWM8krKE4zhikSymLZwuU1bx/DG0dW5emvZzmJzNggB9OOSoLG9M5UOVSp+g9DJ
LWIpJ7SMWqo8X2gnOjlDkzJCLqdRw8wrXZ6MXuoTayNbM0yf9I4u/f23CDLXjtPSY4YxCtLPs1Gw
DmRjpO4yq/rwfG21S0c8urzQJxDwt/TxU0bkbcin1NA5xmYcCUoVME0upXBmQVwGzTxUn2LkFpGh
xmUIqPhXQZswtLh3mGHe5KMfNBG6btu4l/G0RUh9WanDxi1spnJte/zIpOf5jvi+eB5dXBZz+xbN
RojWULi4ZjJtKPqVpD4kwekMMFAFipIwtOzjCs5r4QHYUlXmlja11f43ZxFWA7ouucweWXC+qWH0
LHR7dN8iYeRYXLrYjfkivY2vWQ0N3Rux+5QK7wCjAlG7/9bfSKIrIvhfzTG4Uu1j2SpbGBKFvitg
S8oiKZanBQ+7133ZY5GLTvdL7kvaF+8s1G+oiRlzhKRhVV+q0NtSg10K0DVwtaMhRZfgBx3Y2bFh
HSiObwg4aBluycuKYEF5x4wmB+5hT1BFIgXijhDqVD7jz2kuq6OcDba/N2Qre0Opd5EktM5sN5zv
+ZGP1wKzJCpQXJgNui1kVCKHqIZ9IY4WxZE2t49e4PrIDLQTpwLR+7oudUkEZR63QBlRMS/4tFO/
jcEqZc9UQIb/NjRj+3Spe53Co580vlRfd/6czB9aBtk+YXOakXBlSLXoL0471siojUDVIIX0q9Fk
IgA3TG5dEF4vmZKs66nU03mgp9+CRVahIZ2KKK/le67Wm5y0lYe09a7bNZd/T3zFi4gDVXJYZG07
V7DlCKjhGa+6R0OkcqML/j86k/vQYSPu0P5v0IZXiaXZuejdv2VK0UxvHFYRqoa+1A/ALc/cTY8i
zfAzT8uo00igiwsx5Ur3GDZE86AGY95sZAhOHXcv1bRr6ZjANdnyzP8kTz5O3zMfGLchtP/TdkNi
TWHBuCvMRxkNThs/Cwr8KQF5JickNIhPkCuOLXJRZ0kB/vm5OJu5iqqWeWuymeiGradt6Qdd8UYK
WpE/KXTUNTcWHAvoVOFiyXmw2kaxYtaaFO1pfS0/U/3me1U0gcM396hNnydQK1YB5Ugfgl8ncku2
P9Y0jXDZCsnV5sLTh6MTfmPbaltC3vOvYnmdH+eAqHFnapktTMEnhr6m8vZcAEW1lp0Z94RW67pL
w6ZWasOh39bU1j1jssnGrseYMEdSl9R77bhxnLhWQpuv3tvJLIvArtxnQl0T3bhkigcdEL7W8CrD
F9q99f59DPIE6usBQZjS6H5Y3zVC1/ODJgOjBTEiYViGYaT4v97rV5mzieVnGt6q1+Vtcl0wBef2
V331zYLJBAFZR3Vtlsefp0/Bt6nTkfGW+k6PLUScWvyIptfNfoVnKXvISZIiiZ2lcVQbbcBpuXA2
fZgfsb0LNAf8mEM1p5WhqnfjezJoGLRZZSJMW5is8xGD0zDfQro6GX33jFoMvxCCD/VHYXFVeMbO
WA8JQoNxSpC6oC92LEbYNDJvT/dZnQ/1NtVOCwmP2EKD+vH3dQ4/+ylKTdgBfECzSeVzam/ZB1LR
M89fzrCNxv6S+Nke4JktUkR92z/eXh8wzdvDy8J9ZmkAAUqzBzY5y7BNfJKrBHjYnATI4MHwt+Nv
O/q3z7UnNdn5vOyGIgxETmDN0PvdbO8GMlkydi6bXDsrs3xj/+0IfOhT0Wca7Yjr/GCXO/CeP6l3
WJO2fKzur7yAwF8pJU/nmfNruHdWFMP3QRWMsmjtPaQGdDoM/3d2Nj5Kbjppbw3u+kvY91ZtlL3q
k1wAskAA0KPjLYwDMUAL0S/7EVbT0DttWmLg+grCQiojXeu6zjf5KH9bvXH+9TGcn2oSjWQa/o36
IDTMpE+q6qt/G5KR1GPHdUqjA2UZLLCIxGgEbJKcn2F+CvoOBOIagAIkhk8xw3IhY1Kw5hLmHsyW
Zym749v9YhA+mVyqxvL4k0e4fdCQIduRZsTV9B7wObWZhYXbt+kNvH8NUseok9RiAqJWAYWIxqRo
AXWM+pyEGNvOjgzpL+jEtZQwYHHIpbCBIihP91KJhbMSBjs86dq1TIBSn3F7x5sZXdtOACRoBAYV
hxtf9cQv3aRgRLAd4H+hbP+ndXpikuBhUEJOLG5dKaJmE2U3Qw5id2L0Pa7Y+IXRJ3C6g9H6l6VT
ntwk4AbYxdpJJlMS8Sacb3vdolFNcSTG4ClwdOk7YdOlCck7yseO3wCFiM0kdfJWNk5av4xXVHx4
JOFp6r93tkfO+p0N9ZCLuYGUghOVHYtANfn3XUyL/5ePe05dO6QrN15GVFucq3zSVivgRlvyxCUb
YZ/X4EI3UviCDdKEyE/DGwB+y0Y4+oyJKTTRvOZfWFM39OsrqPSWFe9AtkDz2+71+zMycCwiTC1e
haItOrj6S0HybtFfcTTkh53bx7C3Yohgexw7goVnQ+M+OSPqpKCJ5Bxi+h6X8ueoXa+0o6KPy5He
JJNjZgpQSJZSmJn3wp44M2/mQXKgBgFr+JtJXLODx/bPUySAFq7RGaY0/xefbYLq9vWE6IJR/OcQ
snszswJBkwGSfPVYIdY7BoxnbBXynbLQJ6m2tTDFSvcY97uBscO7Es6XlThMg55oZuzLCm6rYMO7
4echb+Jx+e4jmMjQRnxvEZpLDtpYwaUnwchYpq8nBB/KgVtYe2y/riz03gefTSyNowcF47l0UT2u
dw1ZmgGmo2/obEqkGhUq6eDQaahLMTT84ZoAFEi2wKvndNHo8N1bmGPt6t82L4jJCiGFiD70GoIN
b6yv9KlLWt+PcNHdEfqAK+MFlsGVOyg2rIVbicFv6X/0OsUvCQrEo+Yo7N/NyOkXHpybnWMkzbDK
H7fIv8f9d3Mvcb13JRMIzigvbeFKx0IfCLQbJemYvtqLBNWfllDF+8WajZafbfudzWfcdgAg5OzJ
M+qzXHRLPlVFcWWf1+/+Q3MwHjLZyAF696IaA9xQ2ExlTWEgbG9x93uriXvPElqXxSVTXhCd+z2Y
kSMkwVr2GIImCuNmAzVJ8/HCKmDpR14utFV6hGujY3EQaaEfI/0enkNaVPRdKBfd8C9lGQS6vnoq
e8xwNNYPJaWQlaFxqgdlgkwPZHoQ1KNDBBVLR+8eOkm9EV+HIfYKABV+46gd+39+ZYC+MrJNhXJA
BiYykpTnnif5OmVRTeitOSqhF6T6OjUlpXYugwN1LA8fvT/XzxOUt2yVzNqthtGQR9Mmz3C00J1y
WL8d0zTNkTW+6BWvvOnylfu2Z6LPkXJU3X6uqQN0KBD9GbXQe31C0ajhlVfkHcOIm3Z1pOoafxZL
/4bUvXgg/wPG2T24seEaVbuWnLLvfL6hpfR9l4V7ts27oJJ5hZ3k2ZgV1I6rla/zrNEL5qZ5/cku
Fam2x2xcccgkBnmuCaEEE22/wWc0GmDZ6eZR0Fy6r3wXClWUJUa065V2m0XC6dKDwt+3tXoB5bGM
9n50+lrdK94bAGo7LAOW+fc2CVWRqZxVHUVSzG/roFUmYreEuIdq4KL/d6tXiNzaLX4Ld54fvXjZ
3SypIxRggs/hdPRzz84BCm/uEOorjsD3LdFfQO03hFAl0pYIz6VZo+9wInUbDbT6rlWRCcwp2CQy
ejTzTY3Y0/CmcsfEh5nKREAMZJ+zPb00Ihi+Kp+1mhUn2QzGq0d8B5ZYB/TBD0VNwMc4Oo9Mpxi9
SYhR5ivyHrx98GBCTdR9aRZN60fiukJ0TAYo1FcMDCvbIeZeC2cRZDtJvO7Um2t3YyqelcszaK8U
UAHcVgppMA9CNBIKNddBQGqSNpYaowKLaDMj1Et1N4XTv0uu+zlkAF/WXy+Im25GBesISa+IJf6S
GCrMFbHpigx3T/8+d7eYJ/Ck6s7q6iN0MG4rPElKjIWzZB+VRYCP1IvWScUK9a0ZueNH3MphX8xW
mQthp5hYqPatDVkm4XXu7Mqaq7G/wASNKi5cgJiCw1DaYeGqP4ypmZ0/Y9X1mPBWJzf5tK7iT2rx
iVC477dvJdK125olLyaZ+Dk5iZApIiYUMz9rAMattoRfk9kc58KALGiI5LjYnTrlNLo/VzHuZyST
oRGdMHSu7jPbzIGl64U3RamCl85Uq2yVvMFN6WwjjqCzoShoW9plaamEAUatmn3fb0Et55gyrg6X
90thVTt9fe1+R3jjaTWCTP74o7isGxmgtNJb6eqtEV8k7RCogG1r35593CJceMEUN71Vwj/TaPFr
dcclt9x77JxegvjBrLjDqgnRFvJuvezNZeTXVL2NQySwRSUDAz/knt6F80NpMHY6JLgVQbZqAvKe
tXTJ8ZydMhlw4aKU0AaKrb2N30vFK4wbQHTIlTnj/awa6kGEozUA2jFFYvAulOhiMB81RNMlO8G5
h0aqN/f4q041UsIrQ5H4oeTd40gtgz10F54tnrDTCQEtcMEI8hh8MVhCsJUygt7fU3UhMR0cNOXU
AENeDoHRm+2Oinzuwt/F7o/ecfj+pbHl4QKCU7ZBES/m9yflhsHbGRyUson3gbR9BB9dlbzTCy8R
6sIRw/pHm9wDFpq9iLDBg2FWcNzZrz/4V9W5wgIjivwyHhhudFDo1KFGLZ3WAk5zdSGTYJF4FmJv
DUQouImgr8AJOwpgC4l93Uurvq1qhD2dqxvFMi7007LImw6HGYTJYTWrTdxfrOrDnvBIoTuEyHI3
d8TuYC26wcLhvITgFNwg9lmOkHMls5ycsReBpDM5kBKkCspiyxUxs+WyPL3QVbwnpYfl/wdm8Sqo
LD1zppQB/igAYWCMlNaRH8dTFoNW0vrC6XxemgukqLvWAfZ1WNHQyXAdYPSc8MrtkGXZfg0Bo6Uq
TXYeMoE1XKqHl5W5wdzhu1KfysYPd9OBSbjG5/TgRVatBO9+qebOL6gN1cYIxc4fKurecLx1rGYt
P/pQw8HAz2BfYQWkLd4TvJVrt4nw0ndD0DQSIFz67Dz+T35h51BI7ZkXkUh6S5XhRNcHueWUn+7J
ZxNE8qJwy2YGFicrCQwFXBSVGiwr64vlEyp7S73HyGB0mHX2IF8nBAMqFeK+08BMY5phEXPCPC4t
Xm8srqcGwXk9nWV9RfSShUQ6eRlRs1S+sc0nCCnbkQETln1rgza7WZ0teQWA+rnJ8vSRVs6fqJRX
OAq8Trj4iUUF0KNbGhhiHY1mVL8fJbJwPmySNaG6vHaCDzfE3j8XD+oHIB3D/btqx7q9G85X3Acg
cuMMm+C1i8YwUQmxb9txlGMFGewjpa5IyukldojW5xB0qvNa/mfSJ6Z97Ck8yCwoplhNlxXY0P5L
8Rc7eqHYKkgzkgUu/nGtUrEEmLzxlBUqwR9b4jRhzfE3w23b8X3sVKcNC2Dy5+ItizSsmUP0YgRT
CcUA83KD+ub3BWxEO9b5QwCMgWIfQskof79xs+Px99rYumVI0P8KX7JLWmOmnL0HG7Kc9jw7QLk9
BhMYe/FEjYB/uhosbXR5GgEKkOqyg+WBQtHztctqj7xiIxwE1ashQuQJiVY4BR55XpAMGZlI7zWU
PckAPUlHrSSeg5RZ5QI7wSSSDaNdsuS0E4dyqrlcBmoHqIMBMr/Vr+rENXfE/l18MOid2rUAjj+P
VfL2vLxI2uLTg67YKiJJ/Bdt+PlQWARFuVSaAN2KUxrKtY401Zj2HsKrpkIcuOvBy8GxLuGuxf3u
NG5lA31KhOcw
`protect end_protected
