// megafunction wizard: %FIR II v17.0%
// GENERATION: XML
// fir_2_10hz.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module fir_2_10hz (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [12:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [47:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_2_10hz_0002 fir_2_10hz_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="17.0" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="nsym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="50" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="0.00025" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
// Retrieval info: 	<generic name="speedGrade" value="medium" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="frac" />
// Retrieval info: 	<generic name="inputBitWidth" value="13" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="7.772445678710938E-5,5.2809715270996094E-5,6.842613220214844E-5,8.511543273925781E-5,1.024007797241211E-4,1.1944770812988281E-4,1.354217529296875E-4,1.4972686767578125E-4,1.6117095947265625E-4,1.6891956329345703E-4,1.722574234008789E-4,1.704692840576172E-4,1.6295909881591797E-4,1.4960765838623047E-4,1.2993812561035156E-4,1.043081283569336E-4,7.30752944946289E-5,3.707408905029297E-5,-2.9802322387695312E-6,-4.589557647705078E-5,-9.02414321899414E-5,-1.347064971923828E-4,-1.7786026000976562E-4,-2.180337905883789E-4,-2.5403499603271484E-4,-2.846717834472656E-4,-3.091096878051758E-4,-3.2639503479003906E-4,-3.3652782440185547E-4,-3.39508056640625E-4,-3.355741500854492E-4,-3.2579898834228516E-4,-3.110170364379883E-4,-2.9277801513671875E-4,-2.7251243591308594E-4,-2.5177001953125E-4,-2.3233890533447266E-4,-2.1564960479736328E-4,-2.028942108154297E-4,-1.9502639770507812E-4,-1.926422119140625E-4,-1.957416534423828E-4,-2.040863037109375E-4,-2.1660327911376953E-4,-2.3186206817626953E-4,-2.4819374084472656E-4,-2.633333206176758E-4,-2.7489662170410156E-4,-2.802610397338867E-4,-2.770423889160156E-4,-2.6285648345947266E-4,-2.3603439331054688E-4,-1.9490718841552734E-4,-1.386404037475586E-4,-6.73532485961914E-5,1.8358230590820312E-5,1.169443130493164E-4,2.2614002227783203E-4,3.427267074584961E-4,4.6312808990478516E-4,5.830526351928711E-4,6.979703903198242E-4,8.033514022827148E-4,8.945465087890625E-4,9.675025939941406E-4,0.0010184049606323242,0.0010443925857543945,0.001043558120727539,0.0010149478912353516,9.588003158569336E-4,8.764266967773438E-4,7.704496383666992E-4,6.444454193115234E-4,5.029439926147461E-4,3.510713577270508E-4,1.94549560546875E-4,3.9577484130859375E-5,-1.081228256225586E-4,-2.429485321044922E-4,-3.5965442657470703E-4,-4.5430660247802734E-4,-5.234479904174805E-4,-5.651712417602539E-4,-5.788803100585938E-4,-5.649328231811523E-4,-5.252361297607422E-4,-4.627704620361328E-4,-3.8170814514160156E-4,-2.866983413696289E-4,-1.8334388732910156E-4,-7.712841033935547E-5,2.6226043701171875E-5,1.2135505676269531E-4,2.034902572631836E-4,2.6869773864746094E-4,3.1375885009765625E-4,3.371238708496094E-4,3.3783912658691406E-4,3.167390823364258E-4,2.752542495727539E-4,2.162456512451172E-4,1.4328956604003906E-4,6.0439109802246094E-5,-2.7418136596679688E-5,-1.1599063873291016E-4,-2.0039081573486328E-4,-2.7680397033691406E-4,-3.414154052734375E-4,-3.9184093475341797E-4,-4.2617321014404297E-4,-4.438161849975586E-4,-4.450082778930664E-4,-4.309415817260742E-4,-4.0400028228759766E-4,-3.669261932373047E-4,-3.230571746826172E-4,-2.759695053100586E-4,-2.294778823852539E-4,-1.8680095672607422E-4,-1.512765884399414E-4,-1.2505054473876953E-4,-1.0991096496582031E-4,-1.0657310485839844E-4,-1.1491775512695312E-4,-1.3399124145507812E-4,-1.6200542449951172E-4,-1.964569091796875E-4,-2.3448467254638672E-4,-2.726316452026367E-4,-3.077983856201172E-4,-3.3676624298095703E-4,-3.566741943359375E-4,-3.6537647247314453E-4,-3.6156177520751953E-4,-3.4439563751220703E-4,-3.142356872558594E-4,-2.722740173339844E-4,-2.2041797637939453E-4,-1.6129016876220703E-4,-9.810924530029297E-5,-3.457069396972656E-5,2.5987625122070312E-5,7.987022399902344E-5,1.239776611328125E-4,1.5592575073242188E-4,1.7368793487548828E-4,1.7654895782470703E-4,1.646280288696289E-4,1.386404037475586E-4,1.0073184967041016E-4,5.364418029785156E-5,5.960464477539062E-7,-5.447864532470703E-5,-1.0764598846435547E-4,-1.5485286712646484E-4,-1.9252300262451172E-4,-2.17437744140625E-4,-2.2745132446289062E-4,-2.2101402282714844E-4,-1.9752979278564453E-4,-1.5783309936523438E-4,-1.0335445404052734E-4,-3.6835670471191406E-5,3.8623809814453125E-5,1.188516616821289E-4,1.996755599975586E-4,2.7692317962646484E-4,3.4618377685546875E-4,4.038810729980469E-4,4.470348358154297E-4,4.734992980957031E-4,4.820823669433594E-4,4.729032516479492E-4,4.470348358154297E-4,4.063844680786133E-4,3.542900085449219E-4,2.942085266113281E-4,2.3055076599121094E-4,1.6760826110839844E-4,1.0991096496582031E-4,6.127357482910156E-5,2.5153160095214844E-5,4.291534423828125E-6,0.0,1.2993812561035156E-5,4.2319297790527344E-5,8.654594421386719E-5,1.4257431030273438E-4,2.0706653594970703E-4,2.7561187744140625E-4,3.437995910644531E-4,4.069805145263672E-4,4.609823226928711E-4,5.019903182983398E-4,5.270242691040039E-4,5.341768264770508E-4,5.223751068115234E-4,4.92095947265625E-4,4.4476985931396484E-4,3.8313865661621094E-4,3.104209899902344E-4,2.3114681243896484E-4,1.4984607696533203E-4,7.11679458618164E-5,0.0,-5.9604644775390625E-5,-1.043081283569336E-4,-1.3148784637451172E-4,-1.4007091522216797E-4,-1.2981891632080078E-4,-1.0216236114501953E-4,-5.91278076171875E-5,-4.5299530029296875E-6,5.7578086853027344E-5,1.2242794036865234E-4,1.8489360809326172E-4,2.4008750915527344E-4,2.8324127197265625E-4,3.1065940856933594E-4,3.192424774169922E-4,3.075599670410156E-4,2.7501583099365234E-4,2.224445343017578E-4,1.5223026275634766E-4,6.771087646484375E-5,-2.6941299438476562E-5,-1.264810562133789E-4,-2.2554397583007812E-4,-3.186464309692383E-4,-4.0078163146972656E-4,-4.674196243286133E-4,-5.148649215698242E-4,-5.409717559814453E-4,-5.44428825378418E-4,-5.259513854980469E-4,-4.8732757568359375E-4,-4.3141841888427734E-4,-3.6275386810302734E-4,-2.8634071350097656E-4,-2.0766258239746094E-4,-1.3267993927001953E-4,-6.67572021484375E-5,-1.5139579772949219E-5,1.823902130126953E-5,3.039836883544922E-5,1.990795135498047E-5,-1.33514404296875E-5,-6.794929504394531E-5,-1.4090538024902344E-4,-2.2804737091064453E-4,-3.241300582885742E-4,-4.233121871948242E-4,-5.195140838623047E-4,-6.06536865234375E-4,-6.787776947021484E-4,-7.315874099731445E-4,-7.612705230712891E-4,-7.65681266784668E-4,-7.442235946655273E-4,-6.978511810302734E-4,-6.291866302490234E-4,-5.422830581665039E-4,-4.4226646423339844E-4,-3.349781036376953E-4,-2.2721290588378906E-4,-1.2540817260742188E-4,-3.5643577575683594E-5,3.6716461181640625E-5,8.726119995117188E-5,1.1324882507324219E-4,1.1336803436279297E-4,8.821487426757812E-5,3.993511199951172E-5,-2.765655517578125E-5,-1.0943412780761719E-4,-1.9943714141845703E-4,-2.9075145721435547E-4,-3.764629364013672E-4,-4.4989585876464844E-4,-5.049705505371094E-4,-5.36799430847168E-4,-5.420446395874023E-4,-5.186796188354492E-4,-4.667043685913086E-4,-3.8814544677734375E-4,-2.8634071350097656E-4,-1.6641616821289062E-4,-3.4809112548828125E-5,1.0144710540771484E-4,2.3496150970458984E-4,3.5834312438964844E-4,4.647970199584961E-4,5.484819412231445E-4,6.052255630493164E-4,6.322860717773438E-4,6.289482116699219E-4,5.965232849121094E-4,5.381107330322266E-4,4.584789276123047E-4,3.638267517089844E-4,2.6154518127441406E-4,1.5938282012939453E-4,6.520748138427734E-5,-1.3589859008789062E-5,-7.069110870361328E-5,-1.0085105895996094E-4,-1.0097026824951172E-4,-6.949901580810547E-5,-7.271766662597656E-6,8.296966552734375E-5,1.9657611846923828E-4,3.2711029052734375E-4,4.671812057495117E-4,6.084442138671875E-4,7.424354553222656E-4,8.609294891357422E-4,9.565353393554688E-4,0.0010235309600830078,0.0010575056076049805,0.0010561943054199219,0.001019597053527832,9.500980377197266E-4,8.518695831298828E-4,7.311105728149414E-4,5.953311920166016E-4,4.532337188720703E-4,3.1375885009765625E-4,1.857280731201172E-4,7.736682891845703E-5,-4.5299530029296875E-6,-5.4836273193359375E-5,-7.045269012451172E-5,-5.066394805908203E-5,2.86102294921875E-6,8.64267349243164E-5,1.938343048095703E-4,3.1745433807373047E-4,4.4858455657958984E-4,5.776882171630859E-4,6.949901580810547E-4,7.917881011962891E-4,8.602142333984375E-4,8.943080902099609E-4,8.89897346496582E-4,8.456707000732422E-4,7.624626159667969E-4,6.437301635742188E-4,4.953145980834961E-4,3.248453140258789E-4,1.4162063598632812E-4,-4.4465065002441406E-5,-2.2280216217041016E-4,-3.8373470306396484E-4,-5.184412002563477E-4,-6.195306777954102E-4,-6.819963455200195E-4,-7.033348083496094E-4,-6.835460662841797E-4,-6.254911422729492E-4,-5.342960357666016E-4,-4.1747093200683594E-4,-2.8443336486816406E-4,-1.4543533325195312E-4,-1.1324882507324219E-5,1.0704994201660156E-4,2.0015239715576172E-4,2.5975704193115234E-4,2.796649932861328E-4,2.5665760040283203E-4,1.8978118896484375E-4,8.14199447631836E-5,-6.35385513305664E-5,-2.377033233642578E-4,-4.316568374633789E-4,-6.34312629699707E-4,-8.341073989868164E-4,-0.0010192394256591797,-0.0011790990829467773,-0.0013039112091064453,-0.0013866424560546875,-0.001422286033630371,-0.0014090538024902344,-0.001348257064819336,-0.0012443065643310547,-0.0011039972305297852,-9.367465972900391E-4,-7.538795471191406E-4,-5.674362182617188E-4,-3.9005279541015625E-4,-2.332925796508789E-4,-1.081228256225586E-4,-2.276897430419922E-5,1.6689300537109375E-5,7.3909759521484375E-6,-5.030632019042969E-5,-1.5270709991455078E-4,-2.932548522949219E-4,-4.6253204345703125E-4,-6.492137908935547E-4,-8.404254913330078E-4,-0.0010228157043457031,-0.0011833906173706055,-0.0013103485107421875,-0.0013937950134277344,-0.0014265775680541992,-0.001404404640197754,-0.0013267993927001953,-0.0011963844299316406,-0.0010194778442382812,-8.052587509155273E-4,-5.652904510498047E-4,-3.1304359436035156E-4,-6.270408630371094E-5,1.7154216766357422E-4,3.764629364013672E-4,5.407333374023438E-4,6.554126739501953E-4,7.150173187255859E-4,7.175207138061523E-4,6.645917892456055E-4,5.617141723632812E-4,4.177093505859375E-4,2.4402141571044922E-4,5.424022674560547E-5,-1.3649463653564453E-4,-3.1304359436035156E-4,-4.6122074127197266E-4,-5.682706832885742E-4,-6.238222122192383E-4,-6.209611892700195E-4,-5.567073822021484E-4,-4.316568374633789E-4,-2.505779266357422E-4,-2.205371856689453E-5,2.4235248565673828E-4,5.282163619995117E-4,8.196830749511719E-4,0.0011005401611328125,0.0013545751571655273,0.0015674829483032227,0.0017271041870117188,0.0018246173858642578,0.0018552541732788086,0.0018182992935180664,0.001717209815979004,0.0015599727630615234,0.0013576745986938477,0.0011249780654907227,8.779764175415039E-4,6.341934204101562E-4,4.1091442108154297E-4,2.2399425506591797E-4,8.71419906616211E-5,1.0967254638671875E-5,1.6689300537109375E-6,6.139278411865234E-5,1.876354217529297E-4,3.732442855834961E-4,6.070137023925781E-4,8.742809295654297E-4,0.001157999038696289,0.0014395713806152344,0.001700282096862793,0.0019222497940063477,0.002089858055114746,0.002190709114074707,0.0022162199020385742,0.002162933349609375,0.0020318031311035156,0.0018291473388671875,0.0015655755996704102,0.0012557506561279297,9.174346923828125E-4,5.701780319213867E-4,2.3436546325683594E-4,-7.045269012451172E-5,-3.2639503479003906E-4,-5.189180374145508E-4,-6.374120712280273E-4,-6.76274299621582E-4,-6.349086761474609E-4,-5.182027816772461E-4,-3.361701965332031E-4,-1.0323524475097656E-4,1.6260147094726562E-4,4.4083595275878906E-4,7.097721099853516E-4,9.480714797973633E-4,0.0011360645294189453,0.0012568235397338867,0.0012977123260498047,0.001251220703125,0.0011150836944580078,8.932352066040039E-4,5.947351455688477E-4,2.340078353881836E-4,-1.7011165618896484E-4,-5.96165657043457E-4,-0.0010205507278442383,-0.001419663429260254,-0.0017712116241455078,-0.0020557641983032227,-0.002257704734802246,-0.002366781234741211,-0.0023785829544067383,-0.002294778823852539,-0.0021233558654785156,-0.001877903938293457,-0.0015770196914672852,-0.0012432336807250977,-9.008646011352539E-4,-5.756616592407227E-4,-2.9206275939941406E-4,-7.200241088867188E-5,6.651878356933594E-5,1.10626220703125E-4,5.3882598876953125E-5,-1.0395050048828125E-4,-3.5572052001953125E-4,-6.885528564453125E-4,-0.0010832548141479492,-0.0015166997909545898,-0.0019621849060058594,-0.0023921728134155273,-0.0027790069580078125,-0.0030976533889770508,-0.0033267736434936523,-0.0034503936767578125,-0.003458738327026367,-0.0033495426177978516,-0.0031276941299438477,-0.002805352210998535,-0.0024012327194213867,-0.0019391775131225586,-0.0014470815658569336,-9.549856185913086E-4,-4.93168830871582E-4,-9.000301361083984E-5,2.2971630096435547E-4,4.4667720794677734E-4,5.478858947753906E-4,5.282163619995117E-4,3.904104232788086E-4,1.4543533325195312E-4,-1.8846988677978516E-4,-5.869865417480469E-4,-0.0010205507278442383,-0.0014570951461791992,-0.0018631219863891602,-0.002207040786743164,-0.002460002899169922,-0.002599000930786133,-0.0026073455810546875,-0.002476930618286133,-0.0022083520889282227,-0.0018106698989868164,-0.001301884651184082,-7.071495056152344E-4,-5.7578086853027344E-5,6.116628646850586E-4,0.0012638568878173828,0.0018625259399414062,0.0023745298385620117,0.0027714967727661133,0.0030323266983032227,0.003144502639770508,0.0031050443649291992,0.0029206275939941406,0.0026078224182128906,0.002191305160522461,0.0017036199569702148,0.001181960105895996,6.666183471679688E-4,1.9788742065429688E-4,-1.862049102783203E-4,-4.5239925384521484E-4,-5.750656127929688E-4,-5.371570587158203E-4,-3.3223628997802734E-4,3.528594970703125E-5,5.500316619873047E-4,0.0011867284774780273,0.0019110441207885742,0.0026825666427612305,0.0034562349319458008,0.004186153411865234,0.004827737808227539,0.005341172218322754,0.005693793296813965,0.005862712860107422,0.005835890769958496,0.005613803863525391,0.0052089691162109375,0.004645943641662598,0.0039598941802978516,0.003193974494934082,0.0023975372314453125,0.001622319221496582,9.19342041015625E-4,3.3593177795410156E-4,-8.809566497802734E-5,-3.228187561035156E-4,-3.502368927001953E-4,-1.659393310546875E-4,2.199411392211914E-4,7.838010787963867E-4,0.0014892816543579102,0.0022895336151123047,0.00312960147857666,0.003950357437133789,0.0046918392181396484,0.005297541618347168,0.005717635154724121,0.0059125423431396484,0.00585627555847168,0.005537509918212891,0.004961729049682617,0.004150509834289551,0.003141164779663086,0.001984119415283203,7.406473159790039E-4,-5.211830139160156E-4,-0.0017306804656982422,-0.0028189420700073242,-0.0037235021591186523,-0.004392027854919434,-0.004787087440490723,-0.004887700080871582,-0.004692196846008301,-0.004218459129333496,-0.0035032033920288086,-0.0026006698608398438,-0.0015791654586791992,-5.176067352294922E-4,4.99725341796875E-4,0.0013880729675292969,0.002068161964416504,0.0024706125259399414,0.002541780471801758,0.0022470951080322266,0.0015742778778076172,5.350112915039062E-4,-8.352994918823242E-4,-0.0024782419204711914,-0.004315972328186035,-0.00625455379486084,-0.008190274238586426,-0.010014772415161133,-0.01162254810333252,-0.012917637825012207,-0.013819694519042969,-0.014270186424255371,-0.01423656940460205,-0.01371610164642334,-0.012737154960632324,-0.01135861873626709,-0.00966787338256836,-0.007776975631713867,-0.0058165788650512695,-0.003928780555725098,-0.0022590160369873047,-9.472370147705078E-4,-1.1909008026123047E-4,1.227855682373047E-4,-2.93731689453125E-4,-0.0014039278030395508,-0.003202199935913086,-0.005639195442199707,-0.00862264633178711,-0.01201927661895752,-0.015659689903259277,-0.019346117973327637,-0.02286064624786377,-0.025976181030273438,-0.028467893600463867,-0.030125141143798828,-0.030762672424316406,-0.030231952667236328,-0.02843022346496582,-0.02530801296234131,-0.020873665809631348,-0.01519620418548584,-0.008403778076171875,-6.805658340454102E-4,0.007740020751953125,0.016584277153015137,0.025549888610839844,0.03431832790374756,0.04256927967071533,0.049994468688964844,0.056311964988708496,0.061278581619262695,0.06470179557800293,0.06644749641418457,0.06644749641418457,0.06470179557800293,0.061278581619262695,0.056311964988708496,0.049994468688964844,0.04256927967071533,0.03431832790374756,0.025549888610839844,0.016584277153015137,0.007740020751953125,-6.805658340454102E-4,-0.008403778076171875,-0.01519620418548584,-0.020873665809631348,-0.02530801296234131,-0.02843022346496582,-0.030231952667236328,-0.030762672424316406,-0.030125141143798828,-0.028467893600463867,-0.025976181030273438,-0.02286064624786377,-0.019346117973327637,-0.015659689903259277,-0.01201927661895752,-0.00862264633178711,-0.005639195442199707,-0.003202199935913086,-0.0014039278030395508,-2.93731689453125E-4,1.227855682373047E-4,-1.1909008026123047E-4,-9.472370147705078E-4,-0.0022590160369873047,-0.003928780555725098,-0.0058165788650512695,-0.007776975631713867,-0.00966787338256836,-0.01135861873626709,-0.012737154960632324,-0.01371610164642334,-0.01423656940460205,-0.014270186424255371,-0.013819694519042969,-0.012917637825012207,-0.01162254810333252,-0.010014772415161133,-0.008190274238586426,-0.00625455379486084,-0.004315972328186035,-0.0024782419204711914,-8.352994918823242E-4,5.350112915039062E-4,0.0015742778778076172,0.0022470951080322266,0.002541780471801758,0.0024706125259399414,0.002068161964416504,0.0013880729675292969,4.99725341796875E-4,-5.176067352294922E-4,-0.0015791654586791992,-0.0026006698608398438,-0.0035032033920288086,-0.004218459129333496,-0.004692196846008301,-0.004887700080871582,-0.004787087440490723,-0.004392027854919434,-0.0037235021591186523,-0.0028189420700073242,-0.0017306804656982422,-5.211830139160156E-4,7.406473159790039E-4,0.001984119415283203,0.003141164779663086,0.004150509834289551,0.004961729049682617,0.005537509918212891,0.00585627555847168,0.0059125423431396484,0.005717635154724121,0.005297541618347168,0.0046918392181396484,0.003950357437133789,0.00312960147857666,0.0022895336151123047,0.0014892816543579102,7.838010787963867E-4,2.199411392211914E-4,-1.659393310546875E-4,-3.502368927001953E-4,-3.228187561035156E-4,-8.809566497802734E-5,3.3593177795410156E-4,9.19342041015625E-4,0.001622319221496582,0.0023975372314453125,0.003193974494934082,0.0039598941802978516,0.004645943641662598,0.0052089691162109375,0.005613803863525391,0.005835890769958496,0.005862712860107422,0.005693793296813965,0.005341172218322754,0.004827737808227539,0.004186153411865234,0.0034562349319458008,0.0026825666427612305,0.0019110441207885742,0.0011867284774780273,5.500316619873047E-4,3.528594970703125E-5,-3.3223628997802734E-4,-5.371570587158203E-4,-5.750656127929688E-4,-4.5239925384521484E-4,-1.862049102783203E-4,1.9788742065429688E-4,6.666183471679688E-4,0.001181960105895996,0.0017036199569702148,0.002191305160522461,0.0026078224182128906,0.0029206275939941406,0.0031050443649291992,0.003144502639770508,0.0030323266983032227,0.0027714967727661133,0.0023745298385620117,0.0018625259399414062,0.0012638568878173828,6.116628646850586E-4,-5.7578086853027344E-5,-7.071495056152344E-4,-0.001301884651184082,-0.0018106698989868164,-0.0022083520889282227,-0.002476930618286133,-0.0026073455810546875,-0.002599000930786133,-0.002460002899169922,-0.002207040786743164,-0.0018631219863891602,-0.0014570951461791992,-0.0010205507278442383,-5.869865417480469E-4,-1.8846988677978516E-4,1.4543533325195312E-4,3.904104232788086E-4,5.282163619995117E-4,5.478858947753906E-4,4.4667720794677734E-4,2.2971630096435547E-4,-9.000301361083984E-5,-4.93168830871582E-4,-9.549856185913086E-4,-0.0014470815658569336,-0.0019391775131225586,-0.0024012327194213867,-0.002805352210998535,-0.0031276941299438477,-0.0033495426177978516,-0.003458738327026367,-0.0034503936767578125,-0.0033267736434936523,-0.0030976533889770508,-0.0027790069580078125,-0.0023921728134155273,-0.0019621849060058594,-0.0015166997909545898,-0.0010832548141479492,-6.885528564453125E-4,-3.5572052001953125E-4,-1.0395050048828125E-4,5.3882598876953125E-5,1.10626220703125E-4,6.651878356933594E-5,-7.200241088867188E-5,-2.9206275939941406E-4,-5.756616592407227E-4,-9.008646011352539E-4,-0.0012432336807250977,-0.0015770196914672852,-0.001877903938293457,-0.0021233558654785156,-0.002294778823852539,-0.0023785829544067383,-0.002366781234741211,-0.002257704734802246,-0.0020557641983032227,-0.0017712116241455078,-0.001419663429260254,-0.0010205507278442383,-5.96165657043457E-4,-1.7011165618896484E-4,2.340078353881836E-4,5.947351455688477E-4,8.932352066040039E-4,0.0011150836944580078,0.001251220703125,0.0012977123260498047,0.0012568235397338867,0.0011360645294189453,9.480714797973633E-4,7.097721099853516E-4,4.4083595275878906E-4,1.6260147094726562E-4,-1.0323524475097656E-4,-3.361701965332031E-4,-5.182027816772461E-4,-6.349086761474609E-4,-6.76274299621582E-4,-6.374120712280273E-4,-5.189180374145508E-4,-3.2639503479003906E-4,-7.045269012451172E-5,2.3436546325683594E-4,5.701780319213867E-4,9.174346923828125E-4,0.0012557506561279297,0.0015655755996704102,0.0018291473388671875,0.0020318031311035156,0.002162933349609375,0.0022162199020385742,0.002190709114074707,0.002089858055114746,0.0019222497940063477,0.001700282096862793,0.0014395713806152344,0.001157999038696289,8.742809295654297E-4,6.070137023925781E-4,3.732442855834961E-4,1.876354217529297E-4,6.139278411865234E-5,1.6689300537109375E-6,1.0967254638671875E-5,8.71419906616211E-5,2.2399425506591797E-4,4.1091442108154297E-4,6.341934204101562E-4,8.779764175415039E-4,0.0011249780654907227,0.0013576745986938477,0.0015599727630615234,0.001717209815979004,0.0018182992935180664,0.0018552541732788086,0.0018246173858642578,0.0017271041870117188,0.0015674829483032227,0.0013545751571655273,0.0011005401611328125,8.196830749511719E-4,5.282163619995117E-4,2.4235248565673828E-4,-2.205371856689453E-5,-2.505779266357422E-4,-4.316568374633789E-4,-5.567073822021484E-4,-6.209611892700195E-4,-6.238222122192383E-4,-5.682706832885742E-4,-4.6122074127197266E-4,-3.1304359436035156E-4,-1.3649463653564453E-4,5.424022674560547E-5,2.4402141571044922E-4,4.177093505859375E-4,5.617141723632812E-4,6.645917892456055E-4,7.175207138061523E-4,7.150173187255859E-4,6.554126739501953E-4,5.407333374023438E-4,3.764629364013672E-4,1.7154216766357422E-4,-6.270408630371094E-5,-3.1304359436035156E-4,-5.652904510498047E-4,-8.052587509155273E-4,-0.0010194778442382812,-0.0011963844299316406,-0.0013267993927001953,-0.001404404640197754,-0.0014265775680541992,-0.0013937950134277344,-0.0013103485107421875,-0.0011833906173706055,-0.0010228157043457031,-8.404254913330078E-4,-6.492137908935547E-4,-4.6253204345703125E-4,-2.932548522949219E-4,-1.5270709991455078E-4,-5.030632019042969E-5,7.3909759521484375E-6,1.6689300537109375E-5,-2.276897430419922E-5,-1.081228256225586E-4,-2.332925796508789E-4,-3.9005279541015625E-4,-5.674362182617188E-4,-7.538795471191406E-4,-9.367465972900391E-4,-0.0011039972305297852,-0.0012443065643310547,-0.001348257064819336,-0.0014090538024902344,-0.001422286033630371,-0.0013866424560546875,-0.0013039112091064453,-0.0011790990829467773,-0.0010192394256591797,-8.341073989868164E-4,-6.34312629699707E-4,-4.316568374633789E-4,-2.377033233642578E-4,-6.35385513305664E-5,8.14199447631836E-5,1.8978118896484375E-4,2.5665760040283203E-4,2.796649932861328E-4,2.5975704193115234E-4,2.0015239715576172E-4,1.0704994201660156E-4,-1.1324882507324219E-5,-1.4543533325195312E-4,-2.8443336486816406E-4,-4.1747093200683594E-4,-5.342960357666016E-4,-6.254911422729492E-4,-6.835460662841797E-4,-7.033348083496094E-4,-6.819963455200195E-4,-6.195306777954102E-4,-5.184412002563477E-4,-3.8373470306396484E-4,-2.2280216217041016E-4,-4.4465065002441406E-5,1.4162063598632812E-4,3.248453140258789E-4,4.953145980834961E-4,6.437301635742188E-4,7.624626159667969E-4,8.456707000732422E-4,8.89897346496582E-4,8.943080902099609E-4,8.602142333984375E-4,7.917881011962891E-4,6.949901580810547E-4,5.776882171630859E-4,4.4858455657958984E-4,3.1745433807373047E-4,1.938343048095703E-4,8.64267349243164E-5,2.86102294921875E-6,-5.066394805908203E-5,-7.045269012451172E-5,-5.4836273193359375E-5,-4.5299530029296875E-6,7.736682891845703E-5,1.857280731201172E-4,3.1375885009765625E-4,4.532337188720703E-4,5.953311920166016E-4,7.311105728149414E-4,8.518695831298828E-4,9.500980377197266E-4,0.001019597053527832,0.0010561943054199219,0.0010575056076049805,0.0010235309600830078,9.565353393554688E-4,8.609294891357422E-4,7.424354553222656E-4,6.084442138671875E-4,4.671812057495117E-4,3.2711029052734375E-4,1.9657611846923828E-4,8.296966552734375E-5,-7.271766662597656E-6,-6.949901580810547E-5,-1.0097026824951172E-4,-1.0085105895996094E-4,-7.069110870361328E-5,-1.3589859008789062E-5,6.520748138427734E-5,1.5938282012939453E-4,2.6154518127441406E-4,3.638267517089844E-4,4.584789276123047E-4,5.381107330322266E-4,5.965232849121094E-4,6.289482116699219E-4,6.322860717773438E-4,6.052255630493164E-4,5.484819412231445E-4,4.647970199584961E-4,3.5834312438964844E-4,2.3496150970458984E-4,1.0144710540771484E-4,-3.4809112548828125E-5,-1.6641616821289062E-4,-2.8634071350097656E-4,-3.8814544677734375E-4,-4.667043685913086E-4,-5.186796188354492E-4,-5.420446395874023E-4,-5.36799430847168E-4,-5.049705505371094E-4,-4.4989585876464844E-4,-3.764629364013672E-4,-2.9075145721435547E-4,-1.9943714141845703E-4,-1.0943412780761719E-4,-2.765655517578125E-5,3.993511199951172E-5,8.821487426757812E-5,1.1336803436279297E-4,1.1324882507324219E-4,8.726119995117188E-5,3.6716461181640625E-5,-3.5643577575683594E-5,-1.2540817260742188E-4,-2.2721290588378906E-4,-3.349781036376953E-4,-4.4226646423339844E-4,-5.422830581665039E-4,-6.291866302490234E-4,-6.978511810302734E-4,-7.442235946655273E-4,-7.65681266784668E-4,-7.612705230712891E-4,-7.315874099731445E-4,-6.787776947021484E-4,-6.06536865234375E-4,-5.195140838623047E-4,-4.233121871948242E-4,-3.241300582885742E-4,-2.2804737091064453E-4,-1.4090538024902344E-4,-6.794929504394531E-5,-1.33514404296875E-5,1.990795135498047E-5,3.039836883544922E-5,1.823902130126953E-5,-1.5139579772949219E-5,-6.67572021484375E-5,-1.3267993927001953E-4,-2.0766258239746094E-4,-2.8634071350097656E-4,-3.6275386810302734E-4,-4.3141841888427734E-4,-4.8732757568359375E-4,-5.259513854980469E-4,-5.44428825378418E-4,-5.409717559814453E-4,-5.148649215698242E-4,-4.674196243286133E-4,-4.0078163146972656E-4,-3.186464309692383E-4,-2.2554397583007812E-4,-1.264810562133789E-4,-2.6941299438476562E-5,6.771087646484375E-5,1.5223026275634766E-4,2.224445343017578E-4,2.7501583099365234E-4,3.075599670410156E-4,3.192424774169922E-4,3.1065940856933594E-4,2.8324127197265625E-4,2.4008750915527344E-4,1.8489360809326172E-4,1.2242794036865234E-4,5.7578086853027344E-5,-4.5299530029296875E-6,-5.91278076171875E-5,-1.0216236114501953E-4,-1.2981891632080078E-4,-1.4007091522216797E-4,-1.3148784637451172E-4,-1.043081283569336E-4,-5.9604644775390625E-5,0.0,7.11679458618164E-5,1.4984607696533203E-4,2.3114681243896484E-4,3.104209899902344E-4,3.8313865661621094E-4,4.4476985931396484E-4,4.92095947265625E-4,5.223751068115234E-4,5.341768264770508E-4,5.270242691040039E-4,5.019903182983398E-4,4.609823226928711E-4,4.069805145263672E-4,3.437995910644531E-4,2.7561187744140625E-4,2.0706653594970703E-4,1.4257431030273438E-4,8.654594421386719E-5,4.2319297790527344E-5,1.2993812561035156E-5,0.0,4.291534423828125E-6,2.5153160095214844E-5,6.127357482910156E-5,1.0991096496582031E-4,1.6760826110839844E-4,2.3055076599121094E-4,2.942085266113281E-4,3.542900085449219E-4,4.063844680786133E-4,4.470348358154297E-4,4.729032516479492E-4,4.820823669433594E-4,4.734992980957031E-4,4.470348358154297E-4,4.038810729980469E-4,3.4618377685546875E-4,2.7692317962646484E-4,1.996755599975586E-4,1.188516616821289E-4,3.8623809814453125E-5,-3.6835670471191406E-5,-1.0335445404052734E-4,-1.5783309936523438E-4,-1.9752979278564453E-4,-2.2101402282714844E-4,-2.2745132446289062E-4,-2.17437744140625E-4,-1.9252300262451172E-4,-1.5485286712646484E-4,-1.0764598846435547E-4,-5.447864532470703E-5,5.960464477539062E-7,5.364418029785156E-5,1.0073184967041016E-4,1.386404037475586E-4,1.646280288696289E-4,1.7654895782470703E-4,1.7368793487548828E-4,1.5592575073242188E-4,1.239776611328125E-4,7.987022399902344E-5,2.5987625122070312E-5,-3.457069396972656E-5,-9.810924530029297E-5,-1.6129016876220703E-4,-2.2041797637939453E-4,-2.722740173339844E-4,-3.142356872558594E-4,-3.4439563751220703E-4,-3.6156177520751953E-4,-3.6537647247314453E-4,-3.566741943359375E-4,-3.3676624298095703E-4,-3.077983856201172E-4,-2.726316452026367E-4,-2.3448467254638672E-4,-1.964569091796875E-4,-1.6200542449951172E-4,-1.3399124145507812E-4,-1.1491775512695312E-4,-1.0657310485839844E-4,-1.0991096496582031E-4,-1.2505054473876953E-4,-1.512765884399414E-4,-1.8680095672607422E-4,-2.294778823852539E-4,-2.759695053100586E-4,-3.230571746826172E-4,-3.669261932373047E-4,-4.0400028228759766E-4,-4.309415817260742E-4,-4.450082778930664E-4,-4.438161849975586E-4,-4.2617321014404297E-4,-3.9184093475341797E-4,-3.414154052734375E-4,-2.7680397033691406E-4,-2.0039081573486328E-4,-1.1599063873291016E-4,-2.7418136596679688E-5,6.0439109802246094E-5,1.4328956604003906E-4,2.162456512451172E-4,2.752542495727539E-4,3.167390823364258E-4,3.3783912658691406E-4,3.371238708496094E-4,3.1375885009765625E-4,2.6869773864746094E-4,2.034902572631836E-4,1.2135505676269531E-4,2.6226043701171875E-5,-7.712841033935547E-5,-1.8334388732910156E-4,-2.866983413696289E-4,-3.8170814514160156E-4,-4.627704620361328E-4,-5.252361297607422E-4,-5.649328231811523E-4,-5.788803100585938E-4,-5.651712417602539E-4,-5.234479904174805E-4,-4.5430660247802734E-4,-3.5965442657470703E-4,-2.429485321044922E-4,-1.081228256225586E-4,3.9577484130859375E-5,1.94549560546875E-4,3.510713577270508E-4,5.029439926147461E-4,6.444454193115234E-4,7.704496383666992E-4,8.764266967773438E-4,9.588003158569336E-4,0.0010149478912353516,0.001043558120727539,0.0010443925857543945,0.0010184049606323242,9.675025939941406E-4,8.945465087890625E-4,8.033514022827148E-4,6.979703903198242E-4,5.830526351928711E-4,4.6312808990478516E-4,3.427267074584961E-4,2.2614002227783203E-4,1.169443130493164E-4,1.8358230590820312E-5,-6.73532485961914E-5,-1.386404037475586E-4,-1.9490718841552734E-4,-2.3603439331054688E-4,-2.6285648345947266E-4,-2.770423889160156E-4,-2.802610397338867E-4,-2.7489662170410156E-4,-2.633333206176758E-4,-2.4819374084472656E-4,-2.3186206817626953E-4,-2.1660327911376953E-4,-2.040863037109375E-4,-1.957416534423828E-4,-1.926422119140625E-4,-1.9502639770507812E-4,-2.028942108154297E-4,-2.1564960479736328E-4,-2.3233890533447266E-4,-2.5177001953125E-4,-2.7251243591308594E-4,-2.9277801513671875E-4,-3.110170364379883E-4,-3.2579898834228516E-4,-3.355741500854492E-4,-3.39508056640625E-4,-3.3652782440185547E-4,-3.2639503479003906E-4,-3.091096878051758E-4,-2.846717834472656E-4,-2.5403499603271484E-4,-2.180337905883789E-4,-1.7786026000976562E-4,-1.347064971923828E-4,-9.02414321899414E-5,-4.589557647705078E-5,-2.9802322387695312E-6,3.707408905029297E-5,7.30752944946289E-5,1.043081283569336E-4,1.2993812561035156E-4,1.4960765838623047E-4,1.6295909881591797E-4,1.704692840576172E-4,1.722574234008789E-4,1.6891956329345703E-4,1.6117095947265625E-4,1.4972686767578125E-4,1.354217529296875E-4,1.1944770812988281E-4,1.024007797241211E-4,8.511543273925781E-5,6.842613220214844E-5,5.2809715270996094E-5,7.772445678710938E-5" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="frac" />
// Retrieval info: 	<generic name="coeffBitWidth" value="32" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="23" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="frac" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_2_10hz.vo
// RELATED_FILES: fir_2_10hz.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_2_10hz_0002_rtl_core.vhd, fir_2_10hz_0002_ast.vhd, fir_2_10hz_0002.vhd
