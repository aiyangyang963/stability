-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cxG4GDYEInwLYZG/7jT6WmmzGVIKWdIbLfGw0vvux63eoGVt0gOWDTnRd8EdvF37yt6bkHVseDDS
2/fZJI5bLy35MdBMudV6KMxGGft7yLPrEkJs0r+W0/Cq5KDisOaNa78QY39fljvRCVBzVFJWCj1H
5xakuLs+zw0gAB9rSqcQFsQwJuKFphJQqwz0Lj/YWzYtoyRGylIRfJWArpP+nCdG60qBKZEe+Jle
iY091abFsGLvfKeq9B+RGSUR28cOca9m7JGoW4bjIZLmA6xSlujPdNahqlyeEdw5OIBHCL2jDmZC
gWFIlDaktQAtXt9VbFQds6e8sdRDJvAgXemhVg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
Y3bIRN8zzGA7DS16pSCsTxl+pKTn78pd3x2wcGR/A78Fm/uxert7giXvJuu8BiRuCRLR/CtdxfPv
kqMbaPgMBOeEjJOHgy8CdZqu428c9O8aCdexscfh0Um6CsZEQY3xNwTKlG4hTWUSHx6OsTSbem7E
SE/vPe8rUBCdrzP4o+yBRQ0r0bG/WJ/vpVey2sBrLFcDoSnlMs/5X2K4gsg8oMmwExgrIfkChP0m
R+IMmpKecyLaNEyPuI4AT1IMErrMwBk7ZSPX7nA/vcI/DsGpPrWPYs/MnjcS7Jix2l+48q/M3I4z
xdT1aEbw8hUcXOI082YS2vF6aoAfafrvMhds/Os2Pn4E9fnYh8ygEDXfSlNPWI6JsijlWRQO4v45
HCE2cqX1mhDOMuF2/QP/aDZ4WC/Ma/lKJYKpjlpbHhEmIGfyN6UR47luHPjiACR2RbldjjyUO/u/
2QlD08dVYmoI/LUgJYYQkSmOUG8knRvhDDLZOkF0OwmexxVcuGfm8wOsVA0RLqXfGc88Gu0iAkuh
5e768zMmeaii86islUdYEBtrt+09/o+7gb8dpOEHm4epdQNwTl92nc92xDrV3uEqbiTNaN9rFQUe
+qnSbvBcfljYyipKIW5LLdJV8KABK2Jz2bh/Z3jPg1fhOO4CPFhUQ9aBnX7Uk8xZn3kxCKIA7jbB
TX3bqxIzG8tzRBb6BTSJcxCiqnx099PWYoAks37fzK9MrItUyQc2Kyl57uDm87GeJwYWYDbpcVP+
do7p4gsjMRNhbrZ7cqQGRV54PY/XqkBuv5KSE1C972NygLRfJ+K+t2CWWnBZFNr2pG8cav6WG595
QNERh5H6f+MryIK0qBPSVTX7vxrWsEQxCxlgj4qvkbG6DfPl43JCWyzI9YuiZaFk3ngnJKKPQiSV
kNMcD5nyYORsge/1ZmEpnfEnvYKp/VQzzzqQGbjT642Nopa5LsapHLC2rDpcmbrvQymEcYEMGTPH
qNwt7Fm974sD85sus/uWz+uFqIzi94G6FyXdQiALg5cdLdsyIQL0Zct7NOpF3Ds8cS4XBr6Cd1Zu
KyrZw/Th0AoFWG2uocbKDV+VMwnXSUKcBRqsW5NMe+lPfF48r8v37XD9I/1K2rO1BFyWN0kqySyr
BkRKjBN/2VIkh0vvgj7YlekoD+ggPNiLx+vl3/4vucsJmgicxgyYv1L8FAPFBp6OO8Ehr16dTnyF
14AKcz/nXHkW3rCcORqvk8i6GNAGoXpjNMjIRTQsi6+EYp2AAl/jMgjLlj8GcjLI5YieL0xP63IN
fegChVoiYr2Cnwkr+QS4tgLWupaE6A+a1WVmEftBc8GCQIVdc57bUhD4iWtUpuBiWzfyUQGlrFcQ
Jyo1ROIijm6YAN8LlrFY5/hK+cUhvsuPGGA0ngZonffpEJc+1beQKbn+3uLuxiJsBgL4wYYIViGW
vMoi4R9+DETe1WfKXUxuQPsjIm7JnZmvcas4f7ETnsVGdM6DkEBaNIpzQC7s8u7eFISFtQqpi/cW
3u2AxuKcjLbc+VGaOWNYj49KJ3UHOZxnMMX5mVvnWJ3LQHGH1J+Ht+64IJbpndvCiFl07RFjKDTD
yCwYl+aVo3movu15qXGwXNHcF2NMs5Xsoj7v2BvJnhXgE/Bhilwjl5UxOCYxxlNfDqB3UjqIetJc
TvQs2MmctYlwzknlyx2wgt0NDM65FNDmuieZnsU2BQFACRLhABf3ZB+fVYWpbRHqFkC+R0P9BcLO
spVPX8WyKkUXu2LsN8sQXj2QuEESi1sFb2HMQ7QHoR+wjbHYpSXQD7gDLpsjkS9bbgEU74+hQEDX
X+fFe660FNp9ZjHPTP3AIuTiWgrxjwFtpyfH3OUMBgcBMmMR2Q0/UHv4yYCTDbb1i7uk8YBKgVZB
6wlxbJUGgOGAdlwRPj+CHemYCWFdA52j+kP4FHVSLELobpgbspkF33OG2+ZNOyhOYl6FmZbL5GUv
5bVH2z7gq4dRlW/i0f9+wiL/YwBBKuGoV0Jl+KyicJQpYR/1gmmqedBaSkNlrf+xoEKPoLXdPxYj
ItwquYEzOcHnCcuI+d271XvqaGYXw0HS3PvdUhMP4GaEDtNgWx4X0rJDwy7jj2b5j3kgIDybi0Jc
5SFXyjJv6Jsk2Zf3R79DK6tYk0x6Zesy927UtZSxKW1sEQ+PNI0lVWXZ9sRi94dUQUIYBEvY1fnL
FqDwSv0G90wBYBKyFKSJumDK7uj6FpQ9EOtOChVvMHx7aguDYN+1XoHuuT1ze8syoUThQKNa8L/v
ih34+GEYNDBCQkT2dWx+X6mfvDLafgzahwyakk8o09ar/3xtgZPGeYcsQKGfgjxz6kyB05N2Eigu
WX20ySyAyGSqymQHPaMTnZLOS+jjEZ8w5nckbQT3Cyp8p8eqpWN1U8e9XvQp2IN+aUqa4TQ5dCoz
pRCQw/1DXAHlNKhBRBN0q8Wf443RJWR9lLT8MJ1AabudbzsjspjNtvQj4Zc6mJm4DUzJ5MntSPk2
XoQ35IISidjAl+bP6sYCXP8hTkq0V/GjsIvkwiRGMay1BVe3em093KpAqCxD6FH7exx7O9Wqc2Zw
/9oEFMjnRjuUjWSl4s4md8MtwNI6qBMaahXToG3bwiJLVeyR9yCFKZLtviF9/9iTqFaHeEDhKVDG
b51xlTIUEsV7Q7ZoQ99wZnkEglV9NC/3pkHSyJS/99M3e/MJBfCKbX+PYg6PCGcrRYkvtVK+nlvC
aIPgev1t3RxMIKqzlxy2QRvdMvn4kLFtftDDLo1WHDp+be3PcZqEz4ji8MbuTzKYaKgiKD+ofYMe
zmZwwIxoKemjp5/bMXEe+RLuigKaU2H13mji+9DBFtacZszmGi+Kfwv8sRAdJx6QGBGtuLYGWEMh
sdNbeYhcqcYfHGb5z0VTEn8O2vGj3rHGYJZsk/nlTi0xnygu7324oc5r9CJb4XJSPCXt+dZAoL09
HPDA7xs1ymO6OFM0AUi7OZiMaddXVknczhKCIHMjji+D5xvW0+V8sTRM4axt3XgysCT+0hRG8ikk
RSt/q4yziRpCn/emyJY/H3uuNb9WAoq/kJ5s/lSlPQ5QcdsMymZg5+YcylCc7QmIeIkNToBK8luQ
2niCvUTffENLsbyn/w8ejLDCF8WfoAnzokGAEL7wRYwPUWEVU277duxlkvJU6Ie2WshQvaGoKNCC
JNxhuiNyV7gY8WQyH4068YhtLOB9Sl+wvlLSOj1Uwck40iW7im5O2PsY0V5oIfuAmUkqJEuRZVuz
VPJISkbWWHcVhkoRpxKbrr2d8AbCLstqYs/PLvHA6d3bFjW/R84ngX1AjKnWOxsSx5o5uZ8qQFHf
VsDpnCkp0c+y+1FNG+IOINR5zW1Hfh7uPC6isVco572OniBsG3gbBwydxRFbxZVJTdoLr7lSKqm4
fjdDy08zPaGiJk7ohZJz+vJN4pX1jEKzhW2KP7dli9Vxa79AmECUdTbnaW0NFcDrSHoJydW1MDS0
AN/4HgH1NuDj5DTi/rQl30W7K05gdyFytHRqvTK0OgXfitJe1ekc1Wet2/lPp4E6b0UuvXPTbhQV
qkjggu/mjJRh0TBFqYfXM8c8Lm6weOMiagMs9pZbio3j54VqzNgkKrdCf8tTmKAFXYtuSegSaNrk
FWzPr4u8/K58Je94ecpv9EfBwDUZqlzhpuogsEM75bqMNfqFwezM+aZssHBY47B+2VG5yqdQ4QN5
IqoFeSiJCGHiLjKKu3C0USbpapcNEIbqqEEl8rIdmR/jiTbKgDFj9nrxgtpmmsILYeyJpMt0yJf/
gjBkPP8djGcFWX2HrPWVnkiWVIKzJxBr4YCM+ZCHJ4+TU65zU3Lsva/np1gWpv4y7pdikBSiOlrt
sFPjSoN7kVeCaIdJ2mvmXnYgPlW5yz2aiQjsdcBP5a+axMeZliptA/J+G2jhLKhL1MkM/iRsO0+x
SUfkHK21vWTgTEEEvjV4qlVPNDZE5hg8sq7e/HbRvFITeH6AquynIVHC4jLonNYSz4YSS0PmU+Fu
CSpjJCiI+MBf0DNuOEJ2CL0PJMd8hpDgccqkLpOf1asFnAkDU5bqJoO/9hArCI6pIy9DtqYGz7F8
/HtRpWxKT+3ZlAxoaqZjbTk6K91PoyqK7EDMjaBV0fWKoWauXykVRPD27oM8R98mxi8Erzm8xB5B
oaJ5+/bFYTFX8XrVZBJwLzTB8JLm05QhbDJMqaaCyx0XIC5T77tbG5sOXlrnB1y+Sy/LUxwcadnh
UuoDXeoK8cnP1DGERXaq2s8iyGvw0of/5NX5NJPVTMvBwoEzngsuPQzWK8Ld1NRov2tNbeFuM5XB
kKBzVj5J7AJB0HL/ySfi3oL5Gvc1jDPn4HiaeUM0gUGknTjkCkzSziLxhHgQ82LF3DPxSh0rblwf
EUBXtp7C/PboYq1yD8cA2QNl+hbo0bsVDRnMxQVxkaGy4rf6ZHyIMzPzcqdF9uhuU3jTIqYAvRQU
hiP4CrdqTvJC08xeWp6Np0Zs8WuSpsz520k+Y1KmZOEcaqvR/Ft8+LAiMlX0JhB+GYMSA3cA2v84
K5L6lgmA8ZmJtv/r70q/wPgWhyza1h0pvXdy2c2gR20oAFD0WJo1mHD9sMDstbNljrkKs63+lyl7
sehTaQiqkmHASobG3sIHbeL4JZQd2orL0ykvOWEn0CFX4DOV8r4HUT4EqX17i76xDXX7TsrLkxR5
aTleRqnMx7cff8wvhfpdVf/uxvMUy9vcrntklvS42pQFXoatrDaZv3+VgXzoLIvUVEMW992LmiBT
6Px3EEelbb9vq+FyA3n3X5Z3v11k/axG2oSmkgwB60p6yhqb6XUQnK9KpX1Fxv05Pha0fq7LvU11
Uxg/AcMXpH8IcmAvdvrmgxoLhoGj4mYYwA+JsxguU+LHcvqEwmxhB7xDfGEpgy3rsxPitDpyRC2b
vSZoOHtK0hugUzVXhv9Ruv4sKFSEV4UUexuCINB1kjNDYkjIYC7x8jPGdILHryfYlJQ52VE3OwcO
o/2oR77BfLtb6HNq44Nbo9PtiuSicIsOn90gpAoXKl95yQ6emdo0C4pJTNONVNKweR07hjIDJovv
UWLlgiV/m8XIsNFdPZN6hNxTqX9H1cE5APM82IaFOblU/79aePtJ8ERMXAOM8+5pF5AFHa0NARat
mlDswqk/nKQyTlbVc+Ow9/VNmhE40dFFpTBVm2D/NGH8pULm0I97qF9BD72qAsRIHrxPeLlbAz4Q
3jqDHJnEpoSAQnAb9K2ZmuqKPWF5/Wwbr0rKhmRmVpW6HQWTA1ngS8YwWdR602jFyi0V6nCuiDPi
F4kGOi7kuPVgpkA4uA/4XgKjHHGUiC6FT2UTIMbSaQ9l37N8L7IPyeekU6lx3KXmhaDSMXyljlU4
VCgtsq26kdBPb+K9bVza3n0K4/0vZpOHezwxpnWKKwmBniYof0MlCSRURpN8brrihUYsNMXyRU92
LRvy4+qyjECXOFM7/8h5fQS18y45lizhCZOjFsCRddK9xMsjYIctPn+5RORjQYeD9B69KEhwxtG4
3UpO6P1EuJCby2SmEhZOcstqNFMNcrnxGOPHQWw0k1yOxo5YMCDICnMixtZgvTxfyHGptaLfQKcS
o61kIkMVC1+NAF31PAoI7c749OhL3I86HYWg05T5DRcmeoQClda6Qd3Xsx2HQg1kGPnndU/Cbc7E
93GFh7eWCFvKAddPqukNjK6qo/Y88l/IG7ITrYZpu7jmS2G+JIQG047aTxkGbBqLPF259rabIzKH
GLcISQVp7cfczoomSR4XDpG0HPwq9m0fTwrbzDIdcH5bXtXH0hWGKd2xD4OP+OgfE6Ubpu91Bz8L
+KBEm4dNN1vnWTpAVLfaZXL/j1IWrHnGdZQ/oDR+1a1iHlvO6Q60RZzHZVbUtE3d9Yqn+TFRynD9
ZQQ/v+ykX/fzsaydv/4zcJpXfiJmLU3LAJ5ld2mP5+LBqGPm2mtQ5WdhUWcWfZfR9gLQtyDHurH8
poCA+QahP4GqHXgAl9uBecGKMYNVneu2631Zwj1js2D38L50LhNGQ4+YbONDsiNYrru1yrz6lU+M
JHp21mwpUpNjxcxv+x7J6in2NstLOC4ZCOdCAVr02TOjKfiPOxlLOQAAZrHke8AFlf3UQnMIgTEH
h4Yo6MzWKnX4d+if9FbWzduckqtrr5r5o2hw0vy6dxw+2A4O3Y90Us6b1AnzhEiiVqDdmUseydTp
tErlM24t35078Udmzka1yK7RBRST4zWnJsd+9t42C6/J06M3sMva2BmhH3oBH6GS91KcFdJ4cMGo
/MIqJZaCBF/MPmfHieoMX8F2dAbXZf6/StrLdRv1aFsq/CxYm/H4sOnSAvsZ9C79Ex4S0J0PlitX
y2NDllddAKlFUt+XXsqMvkrUsHvOVhv37xYN8aurZiLMkBRvYrEijGX9w7LRLDL6WJteywCZlxbT
A4LpfB81sCeFB0Xon4yY8q8xlsZZs4pa83KJ8DQjAFGXiVImlq4rXAAIG13HCWRuXGCW2NnK3MoV
RlVH/ZZTzEN6jzh6A/LFImyde5BU/1hShsBlOd2KMBeQv5FGKhqdEjBpnzFnsKUv442E0DE8BBKN
CqRjUp/Ob9brwbU1Vi9UvUZi3QhBkgQpheR7nsq0xQLgTA4gUhVr1eDTG/2o7rE7QDCsv4mT7sJV
ZvB6ZoAYQ0Hq2lhEid+pZGBXQzpIrJqx9iZOUv8y24hecx6AHOIEJ5ooSQjc09/gc+Ljeoat+x3v
eHlterIhaKXF6sgVfXhOhf4vUsuh0fPoypwWi47bo5Lq2Lj4Iks4iHFIPoDmVwXSn2T3yCxb0ge4
oUW8ZbImtG3wHvUc260ac6GomjMP7VOLHfAjowy6Lmp13a0KPx4XIdnC8yRLhLSGIQkhu9gCcjDA
hDPsVtm1Kt33gbPJrm9zWUz795bu9MElOoXjox3up3cd8FrsXcEgbXHsOGvVu8lUD4nF24sYuYVu
j/nCE2TDZr3h9eqmmXFNKtl8i/tgigEVg5Dhy/cRJrEjP46D6glyzeH6dp1pti2Rlr0hASOd7apb
D1dfeJVXf7HeSbohK+jYQHjWUQtiShHznfVeeb6vEmnO+zOYy2bO7Hm/wreqUbfGId/GoJT5Ej+m
1LxN1YNk+HJZ6YB1ms+F8iLazOgjXLHI9/ol5mbDOSmxRIxxPejrmMQ5D4UCQ4nelsqkfdokP5Gx
0hPw4e9IG63lUhaLNjqMBgF+hpYaaD9KwOF1ZiuInYnCI/fSUMyAZ9FpmSy3r8bFvmIoE3QRjwXf
7CpdfbUPkv3yK2Cnp6A938kfxTZXWhWBREXl5SS5ybAb0Fe5IOnuVwwTixMnrXdqv1eS9v45OtIf
EFJiG5nc//Ry9lXDCPHzrS5ksX6XbE55XZljlOkRuia81uFqdxI7PPsoQN/C0zRkTDzD5rP3ur84
eOaMXzuwnZsy0thjyvfqchbduID8fQOjb5U3m5LQ1hcRkxymJi2/tV9QfTog/8GvBWkH7QgxwoIw
EaX5Xn5iRKlB1Y2jydEY8x9qU46oH+bv+WPj4cbDIJVDaNFyd7s5ZIKoziYXcO2p9b6BWwrHKz27
i8x12itTCimzIZ8mjRJabOa00TbdSHbTccIhMxUoZBcdFe6QnkYe8VQ1Z1TqlGXeHBo0AlEIyIbl
DAGXcuETI2zrL5bgrNwfIArCYCH9elnvOuXSyOOqMvWDCmWuU+Ezp+lSb3bBlrFMnpwJRvbCoiVB
VMvx0BAkCFPr6yDNBt5NbDC546GGkr14hTaMDT32URI7yBdp2vnEb1dfWS7WBw93twHRZVLJdEip
R30dVBDI9942ipSqj58Tgh3QSAAJw+xpxThX8wQycXHiLYo7u7iXp/FLFGo97VkBeIlYOr9KxTkc
jVU1rkGCu1jce+BvljBT5AjvOnbvr9goqNc42AmNKl0QdDpjow7s6FY3WhXViEpKQ4jVhwJf7DMU
wSUzV1wiDM1nGNsI68tbHUgEWYPXQLQLNg7VhR0v5snkFWKC/Mw/X96BNVvr5NMbQ7qIVRJfc/8Z
GCtrB3/WsutwUydNHpbc76F91/0JoEUkb7HuC+WkmGk4qdIpFxLy0p2pZdcYIDdwzNZUwOgfTKHk
K7m1bgIeekjtqjHZ7CTxOiOABCBwQ6qgP2/b+JZ7deH7mLptSkILB1a22ZBZ2b1CcaQR160G5/Hy
87+5cNO2r0xjZ5rb7Ne8mfLwCSYZLnvD6ce+zRXaHkL85z4uSgLIGv7VoQnMMcmx4rkmZlmHVqkO
s7gdmd8TKLf7/IvrzGX3mTVuzN2hVDZR3nkzrt6Geo9xn+W6T8u3IH9k2FQQlQUy0tS8R6ckaKzM
xLEL3lSFn689wGwMF10w9Q7F8D0rUU0108IkUqjdq1DTR4m+uKRyaPTTJDFwoVz8aPeUUt9QMZv2
S+Pt1klkFZYvn/78sBeBXDbaRUsmvUevuNttfReqPE+gVLq9oRa4ZCsbydWoNNh7accOh7ccN9cR
36tTrse7HpmRdb2wFVRN7DkTtg9lWDb/NV3wSU0Xk4hIvIuHcTTdjh5PxeCI0TX9pOxoNBDpy3dY
nyTGG2zlRu0rRnmKxKvd9Wot/VCcKsna238sPyU7rNNhoDUQxQp0/aq7K2kOmyJUAWlnzUkhOct6
zUaJOyi1fIXrRjPna1r23xtJkSTZqWcRtDT6Da9PvnlS7yyrS7W/MvciD+Auh7yE2YBSMaqZb0do
UOyUzZNTrs7rXW9n3Ghz9FiNruod1b66ZOxs94Jgk2bdAjw2CLQ0wVdWbeboJ6ozUOIEK0cxMUtv
vrALN6OfdTK5E6sNZa6R3rdhFEDAb4XSbzOBqHNTRiUl+u78yWnzYj2LnfFGMmvNo/OsbFLdr1hZ
On5tnYmcetAJrAaQ2rI9q+pPzl1HhwFgf5yrNGxI1V3iwNomwPxz0KKRl1DKE1uy8zKFEVpa0IRr
AlVNnvGgkMITr7ADhao6CTwfZ8RCMTi3PDTGDeriE8Dg0/BilYetVx8dJ+uyNBZASNfCBJzYTZAF
gasN4nOB75q0J1epitvZTC0hJ2/jya4Onvy11r2GZrL7GxtDNDakGzeo1B8KRt6Z9poCdAUHaGHN
BwsFPqwC8wSdcOhcLMSHgxveATL0ah3Rv50wlOc6FdH4shGMckgrw1sO2T0CYb/50+Pn5f8EteBX
lti3yluth5rL6P1mtS/vroXjSoLPLBULuj3oB2hnhXcx7UlbmzwKXDMZzX8vMP1Cu0mxOcuwRRKy
PofHjTu4xEyVYeC5UvAA6aRMxhFaN3l96+NmUjREQjNdKsENIYDAKVuEoIRSki7yvk551O1xQDTA
m/9T198f8wFGa9fzE8kniELI4N5vezraSezZJCEdxlPkHWWvkZWepkqMmHZrNj0j38hIyJDoBszv
Px+mTeZs69m2QJGDVGE7EaxJRVzCz9btqE3QXuUIxw7i95KNeYDGgoCFmSH0ug6kOZ85ZZEw8ZGH
+sZJrrrrYX/hBORUprezyuwEA+zoi649BHwrpVD4GSWXM2IqsEaS6p4dq+8FW3VwBrjxcXB4tnjd
7vcc/2LlbheBWS2fjkHnY6q2O6DxeKC7Ho1hyfZQfsJHcRKJR9SrVDmJXbF23ElyEw9SkVlS7dOt
IftB7SiE21Z6Q0TVhVhfWa1s5GJHLB7NHz4M67t0jG5xVyC6QEdZx3AImYiSwtxFYXDVtV+nNnsB
W6VIzLSfH/hrGkQV6vzeu4nKBj0SIv13HoS39gQ/N2VToxj3REM8Wr5UPtKWdyFXKjYh8HEh0JiB
LNrB3dEiIuaJecoHWofqbKl77N0WpdbaVScuujhvk6Yv5knIC63T+qJIc7XTqfYLh3z1thwSCGtR
lZhzeKNl5LFTYODTa5Osn9Xz7QS2Qu1wUJ4IB9OK0Ab6frGQQ5xN7ypfnfFTBNApJ63En2hVU20e
v0FfohhfbzcDDMy7nEACeU5CER22T5oNtX5tHsSR41QZv0FFv+BmU2Niv6I8M4d1hwgjt+jnGvu6
XpRZAE5V2CCvhdLhVcSqjLEUklXdcCGD+kLW0+Olw6aCPx8UZ4hEJqsswPDYwHbMVNEfg9zBi70k
T7xg5WF2uXPXGBj7SY4AvTqYJSjx+4GWzcnf97jzFXo7Dd+qiEcbuf2DDcFGjYbegw/Y7j+VJgd2
yRNwQPmNeTgE0ZjFZNoW0KpCOB+YKtJ1MME=
`protect end_protected
