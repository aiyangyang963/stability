-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
auKJckdr0m0yTnn0oLkdh0uEgVncU0KqqGWAxgp8l1wOgCGj0jjMwCNVSCjQe70oj5kCGn3ronCz
y+ngn+8fiSOuEI1asDAbjwBfgQAa2NHg4jTnYyYSDrqjDdLbWIOIOcn2DuHdgsDwySHEUl/RCcbT
DAanTH8yMdBsNl3mo7qRIRe72xN12uIRS3yOhTZsIA6adNMTcOntNbLLxYoghToR0psSGHVklkNS
NxEgcJPNOiUbTJjjUoitX8l2daqrmaBViIRuzV3hWgnv6JBqmEYCJjBhhswndzIEXoKT6IYH4Ehn
+7jq/JG31OHtV5+ANBFUu7nDgZ9t7aX/1ja+2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
ej9Ns18JXlcvUut2KaRTU4yS6zBgtMTZkX2rAJYNKe6nyUpYNNDOcMVbwF/1ruoTxq29QkKeQ12a
f1UXA9meSIJert5Z3Vag4LgGtB2tPhLuSAxjTdnzXlT5AdL8mX396hJ+u4NVZc6uPTsl3auhtfZV
raUv7RgZ9WUqprMnPdrO+ENGC+zkAfxO3lZfnmcsWk1L1EhFLaiOtVday8JZpiN3bFMn8v6sV02k
fUYspk6Bsmv6XWUH8EpMLNXDpR/Qq/8E5bpaxieMS1Ee/iUpDq1NI68iYyF1+Q7b9jfGLH2taYFi
FQvrozozGQMXMyGmevA56CfCl4B4Lj2f8j//y13dQxh8E3rghDdaBM6FQbEKsUyKgZ7uIe9qG0jY
UqWc8hCmKnCTmp2XDTKq9ErOL77I4ljd5hUA4MJ1CO2g5Tm/uvWlHghP8GX+C+D3ZjeLuCfOdMWM
2PmxaNRrD33o2CuKt4rHSwNFnE+wj/cdsXiCPiVQ70xGtY0Wa9HyPfJm7e+sLBfabzikD63ts36g
3TA1UNKRsSjFcPOOVTmsuVmItPmfxVB6NJKvrTX1DjwDncLsy3ZGpqYzZsI5Kv9poGGFoIUz23km
rg89WlOHpx8fLfgrCUyW6ocTR7gd0NlUl8m5WCebNwB3btfhRisXE8azzwl0LMieD0TU+DJd1ZRX
MjKIHl1k+/XEKPJbYC+pm/8H3TYdfpqJIqk/zTKZoVcUZFCY5RPuuF7gh/C8S8cT1dZLBGAMp62N
Y5HM2rRTsuiWBV+H2t0WEgV1w94D4JhxHun0RyYwuM1XISQ3egypSrd4uxuLGd05M0Cnr90Jtc5Q
ayT1GvPBNxnaK/ljL6O00ZJd1ucok/Lz414FYjQjwJITsb+aZBXa6N+Yj6eKEcgUJEFc656NVu1m
wsFh8EABPGBLbpZhHCqJzQ8OOw14XIZn0p3H6HCa72aOhZ350M4L8wnJW73vHQo4J5OVQtndce6Z
eRf6EB2xSGq8+H4SP99yb7cyy0XcZCL7bZP9slVqwltYv+78nYdaEmYmxi8tkAg6rWQ++XyJLexE
OAQ3PV9Fdq7KhEdixCBQpQvtfiaWeuDsjIh/cZlD3QNscdL1fvniEtDn9gUL8ygqTvA5+zQZnjAD
77mXIVpGveLWMfluT4zI+4m2N1eFo9N88vF31YimjHkDg8RhsvM8e7Jq3mKEVPLpdtxh9xNuA1bL
vSfnNJifLMwMlVWPJXDghalM10dtS1DIpuHq4FqLl2bryVY92F7BryNqln+WnMbme49yOG6Paj/m
VQ75FMlnGGHHNBz8XxG0ci9kGqbxuq3C88USPWQB4B5B6C4JmXauYX/OWBYDP/wvYAFlOdIaw7IO
PGl3RoUgyyoYbfT15lacdxZ6HRNL0PZpy780Ywww6X/azjGJ9Ta0ESR4EXqF/7PMyRcJFzsLP3CX
S3cM3aHX3IJWlonhE1WJSsdff3qrRodFzHij8rf9z8GhxHrmlDo2N5GeNnM8ahTyLbUHGxhAwmvZ
kGaXJCImdFgqEhTnp1c95zLOwx0ThlghqehNUgUJXAFLc4nkJ4qC+m2wxWRnARVBPZYHU+x9T/PX
QNuoIZuKPl0lYK3Wvu1KfMBKRfIxJPJlIZnXxH+0Vbkm1JTR12sSKgw6AXTyD4K31C0m3lCuNnam
aprtnV34qwZ+J7ikhpDXDPXk0e6+WM6ePd/zFMKk4TL+iYyZwORF9R7CuTj21o+H5qBz8/JWw/ma
XomEWOypmBJQY4vV1lhRd8HCWmHnX0eD4AkR8Lsid+cLcNOefNSLnYN+XhV5bYR+Nz9gNE9ZeRhh
oTQL2Yx71XIRvpxbLQNX+eUWaa5BSV0aa/lCTLzygq8/DaWxJCsqui3eylrlGpiQ6vBM8Q7XzXUc
L8gKXY3JkpxVVsYGDX2OkbaseV4pNuaj3ocxoQPO9KD3ZRNqs89CSwXPV7P1YGtpJ6xxh4wiIrxB
gXw2t8AIXBRkFS9xjq0JERzO32DgjTtwKMMfI8KE9pUI99a5ZwmNThKspC6ZFr4rogvCvcsBIT6g
S82JwXHAGH7BGmuqcK9UBBHAicxWAP3IgCVFvDWSvXa1IVVwiyZJdHa5NvOPnG00aMPUHNrlJny8
/iSO6OT9PYcQTPnx+e1gj1mKcO5+KpNNOmQ9N55JvyhLRTq02kKTrYtJsYIeaQKli0RmKGsbfv+t
X5HAVj0htLvziEJcTq3hL1GiapYOFe8uWo3CpXwuqfFWD4bCUXaKAdDXji7QDzebqN+1oJzCSKRX
UCz1otdP02weVd4KTTjehiA+PPr6xPXmCRKFIvtLvvMK6xMiGB+bYK3oFLs/qcm5Sr3gxWW5IadU
d+R0P08Vo6R3Ha7wb+QmAJVFOVTIdvCzG1/SotEF3i+HAFAesRjdcWwxmKrrLivF7oySdC5aOnlD
izqdOk9kvsrmfJ5CHeWG71Fd9BcaG3GpE7AHeZTxSSMe5ZSRR7FrrpUpBOmiX/9i6jXR9ghCiRFl
/txjBRlg0VI5lWbGXHllwfkc6KWSSkhU4P56MR7p6JJkEJQzOvF61menyoTrmAxp8dJb784IolQu
nCjtegK6SJkk5zPDqa1H1U4yukOf1cMy6TLizllJ0B15LVnW7883BEUZMKyg+Z+OIAf9n/ttNTHo
c4/ISI6Ci/nhFhT0fE07glc5+LqRUEDNkFrseBcnzFwiaOv6LofSwu6CmImWHlxi2XkPBcQT7hOd
qfVRfjgKGhrTzcCKPXWBV2ulmx0DxsiOHTpTOCA8MnGlKBeqLmLTBuuwNVOfhXbgcNSmc3As3Lbc
ProhhcYmFHslWpjUrA4gj626FI2kalWjJE4IjjCd1ZeDqxFqCT6vBOANp21lSsg/YFIf6G8R+Fow
rl24gCj4ApEuFxk9VR/JkwBAqBnZ3XEIpvEg0v0wut01gcSUsVGB8lF9ZOpmpLnU0d7ETQ2lwXkd
qpdFvcdxzxlo52UGUcdBaXeX/jl3+eMJIWbjQljD+/2iukQZDNH7Xj3NHALZJ4897wlXLWYhIXdp
TiQocYybEP4EUmV5zl6tfu7qP0DEwnSJWscss2u6OCNTibOJape6kdMI5hKVfdyujp3BI60ycvUt
KnroXfn9YZq1GBV0VxERyzINS32j9eFy7jq2fBXuGW2+pl3HFvzpCXEUlUzTlpaoX69Tj42TFldH
7UOTebxnyoOGbbZUm5HUL8HMzQdBzfFfnBpNMzuNWU894SfuOnvGDQruTDz6CettFteYsENy4iHU
EiyHRDGGOgMU2ks38Ki6dAW+m84LtYnUR2dSuHBJ+hosVeulbAFjEN10LlF2jX5Sx65yYFPg+3P/
n8pnr//W1InnSR8skkVjgcwrVlY3MqquDLy3pfJ6JvZT9QEcucRBfGILB2PWKYNH3VPIrQwqYph8
J0WMy8uH5NwLoDY9WGu9NsPSbb+gPX/vI2G+1ZGCvDADEDJLIxXd7olofXv+lLaR2NDV3swz2awJ
qDsMeerUPjEr+iJzouE92RWVcIwgTOX1/Bkyche+uXpDlFudRHj14i3Zz2MkV/gabX8PBe0n5Z46
HdpZ50oUr1xFN+kLrtHn/cg+SkP6PKz3iwtltO0zapyea1kih7ZKtNQMsRQ6Ihs2x4noQ9I4ea2d
aPnHH8Br2dbqiQIt7LmAM62W9e4+SNknUe0s5z4e94/IfTL1km2cxMIQnh178JGlbze7Dbet4VRx
Fv+mpU+K+tr0iGPOACPgB2VGZfxNuAGFhBjHxFWv3mdM3VUT3sPFLUq04uEbU/bGVThFhY/QgOGY
efL8bP4Um4k2/JVQ/USH3y4c59bGjDEnYuD2cpoAcCp4YL3z7xhM6lemM2Wi6N3s9gLrkhUpSLun
aaEWpZq6TVtfzW3ELgZTzYFYDuXtYnUzztoiqEj+QCyyiRKjMTBHJ/bmgOd1H3/JmOU/1BuM04g7
RVaG9O3vNHMeVHUfs0krPEXKsWrjB3YfevlpKD4l2kxLZto6XMrVmi2PTonSuynh3fZVJzFiXvce
8crLApRJghoo455Jq8Fxi8zrNaoEu3giASja/6p9XzUHCjldp798LlkQd7RpYSV1qCquldKL8Xfv
pS0K4UzJYUfJ2M1roYoc0fifViZm7zFWg4g3gcTE/qijz2IM5guT59wA5SoIqL0048ENljb+M6gj
IshXuhLBIN/QHeGbW6WD+pYxN1E8z4jTu3F1fHI/I1IoU+vQcU45y2Y0u4V6OxMwz0jeDmb79G/T
H2YyKhqjIKv4cqvdwi55OfsOwWbRR3cboejQ4oUcfv0VUbiPm+1Z4pYOuyc4uJEegXjUTDx14D4f
KKDG52zAK1VJHSJNUCfaMBNKAemklU9ZpM0pyU0D3bEJoVlDyHoZH2FrpithVD1h8ARBveEQC3Ii
WeexHx2THwhs19MjwvY2ipqZXeUw9rfNbFL+CpMxfcvDLnprTpc6vyvEubo4Rgi1voe+ml8HDjlw
vgNpeRkrmQViEEq6hBEfbcpOgf7m3L1fuOiC8iaiMOZWzmGV/HIRxOKJLt85Yih93who7nMuCsVM
Q2wBcwb1WRAG7rqS42Prp4YSifpXT2D/tTF3kc7m9XBDRPYUhazHqB443dhQK12k95W+8IHN4Wtg
AYplhXdGh4+Fgw4Ye5/FxwPrzj16G6Xdo1/bK0GKn5nMBAdK4BnG7+EiZn0IePo82B4sGV4R1TbY
61Yp2fBcLEPpu538W8HcQIrngTtsWhkOoHzBygYYkDJfYsLAxwL6lX84OVuHnsfIMzBjA3xatWr9
muzfiIzkCVbwiCGW5MeQ+sSaJu9VEijuq3R0gH7P9fyIH8yzDD4yztlZMm98kNNd1Yq9eDDb7l6H
E+IDnDz+7Inf283A52b3HaFTwuhT51x6QQ8alQXKiESRWOi6WZ7lJxspyBqbDyi3tyJV3CtOrfhY
Rdzg2REHl3GMeXCsq/So9UT1REVCjGTDmzOd8iyJlJ7XXAF5UeIbXzOudE9lILSq+saOJqAKLyb8
1atFmbtBKzVEQSq9iaMBE/MuDR1bCZD//0XCH2oq2Hv2AGfOrZkapznCxHIV3HDyMCCRY43V55/v
NzomuOkbX1vnaJFZQ6+Ao1ZBr0mw7sUYeXOBVCNiCGhMXF75tVk8sny8KooQkO5xTSob+gBsbzAM
gMx0x/eU4My0koxxwd4jsACdW02SzknJ5g1QigrloWAc1L6UPKjfjNvCyFYbYAYSb3w6dP7uf8uo
A6zgndwTLej8HfWLIdJRFtt21mImi0H0jPSqiicsRKnA51nNMSx7i4xeobrjWdagSLHeD3JCCz83
0ThpzQ78HVb2KCiIQ6wENKtlXRehPrqED8d9klrhQavxKt6K9hZTq2qxvyiBLCLdLeWHNgnDucPE
FqKaKYZFsaw1/WyfoFm5tB2HkSWpkbliZgbqZLIQHHmeFa9Kgyq+kGt2mE9TMCn+4tVqgwxM9F6t
QwnnbPBar4FGBPwbjgwnZYcWqBrgsSn9vdEsO/9Kb7BISax8Vpn7wXTLrDa/WFKtIClejbH6MZfY
aUn6BxpZrWSE2Z01h8ZaZMLe4voo7QvmSwf9HS/68PY/Ar0bkDNmtBZ5VZfiHTGpzrH13rzIJqdq
VKex4AmK8OanyJ4QXMf5z0N3Zl3vjSh/LC7oQfnIKpCMCwMPQnI7iILWbdMLLsiwbsN2xqhcamse
RVVlrXlinK+2d/r546GxjNf3WE6iZ6pkSs8xrMAjqsMIrF62PEJjpayM/dmrZdZHoeGtDww3j0gM
87M1I08SmHqXpqHGGK0k8aHocYynNoTec5fLMvh17U4C8egFmZ9eXrvXJyrjHT00qEcC2jozeOA8
Wjl3wsuoGfT/DI3y5b1t6OH6T8PtpjIDRCykQBME+15RIKYl0R2QpvoiTVvjwVWVnau9hXS6nA3Z
fD57QYl2SksPXTWRXMXhSlPu7QeEZ/+W6C40AS1IWfJioUl7+OqRgsobrCWkU7Mn7QukdTu0/+HD
eWPu7tsC/cxAwGD4Jwn/eNvSfxYsJVsiBjpZfgJOss3uOUWvlAYJXrbkkAGIkbxXMqyMe4ETHI72
rPRCJnNoptqATw2g/e6Iaqoa23/1kHHSuNVIFE3DUTR04I5EOWMSW5hsNu3krWrpgpyNb+jNbYrR
mUlF5+IRtP12qHkmFIZPysC+2Z7oFbz0yXU62aKAC98dfqPJFlWl+ztPR5TKTtToWKpBArkn9EPl
LYCl0GZPCdEaiNMURzEiLNbR+nGzXHhq5K7NraKH8sSzx+gOO2X0txmK7XwLyl0DROY5UvLwi20j
SN9HrlT52PlJcnGwofzFerogWBqK/SB6FoG9ISQ+l4++Hofrr8ym3yLN7QN1RiRIcZ5jg1it+XfO
oXzTajsb7zIP0m9tWNO+0i77amR64h0nGJ2R4fmtssh0zZQmZ+ZCpV1hrW3rPI4KWTAp2cTC/pfz
aVZt+CyhNne3reQLLPqgTe0chVeEqFUkD935gwSIvpAJe4VFDj8oCpzB4W75CikrFWIZ82GTAa5K
H7Hv1Tj798XDtDIrsP/HeiwDz1GKW1Xlsbbch0EvtZ42b1NGgrg/+8l9LlcFlV2cCvMtFRwnqSIY
sjCh00rmEOt+AMxlIrodabsVwhnrROa3P1oAesER3/0yckvVxzAXvIGA+cjpSLgF1vmzusCliKMv
UA1Xw9l0mEEOVPZ11nOTT4B89pDFubOOYHbC/Zwmms1OrJJsTkoqsgJpMux9s4LUp8iqbKC/amsL
t/iFn1+j4YYXPRxVK9Qi76UdJeBSlMuKybzv+uGDotiXni2euZYti3AHoDwgUGReJYNoTuxPzLMy
yJPtapvVXmo5V5jshPsP5DQP2fR1R1c/cwZd9TkOZG5LHraOnN3+dTl3jIrwDnEnPEpq3k6c+g4s
wizrwy+1DVQ4SM/L4LflcxNKmm1BLWPpehadmxuUrQjjt7P7KWogmWh4YJT4qF7pAcaILkqUTafO
y6/2iqzcIybuSvsRfCveTJ88U3Xarfn6HMvZcsDg3TKAjZ5RK2WSOZe4C475Vl0yr2dZrlRCCxrd
CafIRcBDAf02/M9XZ+zy8OEXhwm2BAEFb7/sYdivnKFhLFcD654H/GXL3CyB/pn12QixKLse2PhH
mAgksSWTevmdLxIxiuV2IS36CjOpsIf3gorusIvdnwOvzsTLgI700zHIaAVMdob1tSO5kz3Xcl0l
IDVbc8AgatI4eVRmrQCaFXcPBve1Tp+TgtmhGrXb9MH3/6bNcIYLVUWeMayg3ZKK0I4dtXW1Vm58
XxJdW9qfCIxPzXBvtvY+FIhs//Apl99eYgw9WUEEzkEy2l2mLBWPHJ0+XDXEO6Tm4yQh3gQnBLwm
uuoXijuDzwLGJlKsnRLzHrj/7aeVucFK0TlDoSrmqrJKZCRxmTgHxKp5PdOr6t1lvhmKhBVl6eTf
on66zj5IlLbGbmKG6iwGgqGohCaMjdZlWFtbJrInzYyRREToTIlIBEtUCRiGmiuBy5s+Vru+mHC4
PZRH3mx6K8QN2Px6vk8dEuUH8cJ2ljK7fqDwNSV7bH+OaRVct2rEQPADxN34dr4A1DrP6FCYaUMC
2H7iSpPTvHMemKb/N5+8GP0eeQCYvKwYhBYz6Snn+gP5t9EWntc6BCHGBT+EYrGs/mwVLaICSeA4
xccjG3Tf/M0DSEbA93L5nJyip3Bm/RpW8BDC7sW523luIHjXa3UgnkQPMmKHUOGbwEFUzetVkwBM
40p4mw95z+6ikGsi/Gzr5/ZXmSrQk4/2Sp4jKn23gdVo75xXsX8LSU0g2Xc4ooNyEs+WnElkUqWT
FtUF8wimRLy1IYA1OxplrYyQiVjdMeTCQ87vLMEJhE2K7hwImNCFgx5ClR0eF646dUI2F328i+a7
vLg3Aen1qeXz4eZo5pLEl1a7Z7lrrRQs6gupTkjoLyA5+vpBSBTKb+hLJzQLbTTDUlxCSU6ALZsZ
+1lQlLKqSEyhi1yGVs5ZIgLvsZmbmuyqvswXAErE+m5gtgOQ0+wu+vzoeJnSFuSk9ZGK7NGkKCtr
fiCcv1xcVePLLGoB0vq0zNlE/LkvDAtI6rU1tdki0OxgWVc0j+hjeLPGlj1cj+FRa4DR21Lo9WiW
ziO/VoB4e1JAOjZWu1kAcYRAjZD+JY61bDlHmRnYYYqcPRrZPdL8sjawPixhDjE3m/8RhXnb+YXB
BFzqOUTsoQid/hiMnUPLEH3AOOLGvuMOEXHpHahq70nDCIgakbRJtsiVH6hCwcxIVz0xcs7WqU+y
Bi2WjVwT1kt3qeYZhUSo6P7J6BTD8mQHKqlJ4rSKKRJT1yDSUT0DZOTBJJ7nzT5t1kgCNeykG1RH
y2OcQsF4X+O1uf8amxd+cB9fV0kwUcC2h+YHhgZ9Ag1ChyTPOEfUHP/hRDwainekupGB5DYSGkA8
JyBBaQRI0Rq1qrR7nD8Vg/6UJUvYyVEMoG7PsFE8GVQXz+hujqevn5jrd62bjHR0OLfq2I6UnXCr
Y59fjAWxwhEwNNZSAUzSizNd1qC6OT6rnDfYRsmFnCxUQDSPSJOIZ/4RI77ot+QnQOazCDbvKMsn
C04x353A9n9oGlRmXyMNOhbs87HBAsr96rVezKEIKfV86YdHQe4+BRsEwQaWwEDa+tYpEDWmTS1T
/1zLutuce7PqRd0aN62zTvTKqXnQtGGilL8+ARhYriBuY1U4aQCckl8Mmi6B55db8XzcHaqCpbSA
uXUZ9rbYUoW99WYZVI9VhrjIP9j1mesAVq675ufH/U65es5oShZ/lLCHNaEFjwelgTi9mEFDJ0aK
MO0Ll2HngNy9QB47yd1xkm0ueZr3HpqospSzEKK0v/8YmOHQ0qm4Wvq1XLSvl7UKhCk10WpkYPGM
IjtMtMGa714jqnVGIhVp2TRf+Y1a6jgtgXmE+CEamxK//dd2sNQoJajomaAOTYpydC57Yeq6MjSY
ftEtDTZ7hj/F2jIhGgh/Q52LKX9Sv9QIiYDTrCbo5vWqiLoH4PP1poc0gvlckNVJwcyGVc08eOWG
2olII+k3y7uX//Jomw6rc6YasrTD49q0qVkRkWPr3eXG0KXeTQ9RrS6lhDpPijDvdOmmbub4cNRX
AfbUD68JE2+CMNpqQsieF+R2AkKmzqWRB51IJPb7mphv6QtvR2faDizGU7iKWfJ3RqPKNYcK838t
q537Ew6DzTHN/UlVvyI23/qc49f8AybUU4dMiLtqGvqLUb/JODEznvIDp76uqMfvf5fkeNcZXx3j
UWOLIaPytiqWlalhSMqr8JJI2IGrsfFqK4oBATHxf5sJ83CLGJfXJxqR/lTgbbV9W1fxnh1gCata
5UO1GdbaF+pjlcnGb52/rCf5Y1Tjnk9V7aYFTuQQUn9aWoURxYqHvMbN01Cab14tdBlvqtby5Omm
ZtpbF6mGeXfF8/sukSlRs5hpsGSPGOyowQ6gLVDKILcbu5bfnYRB+8MlDP/7kim0DOhsbaYVksV9
7+eKMvOnygX6KlRcOCGYGy2RK6zjmTVB+ya5L4A+WXwZEReHUpqeYlK52f4hxxzjHj7NTuIcbKVG
PU/NEyPggZITlfSJFzQJLrJxQlCDHhmjwXXAsUe8ue8514DN1605qQHrPndCKcXLE1xs7sA/FU3Q
C8W60zp9XTetCmJqcTRN2oXJsKz3a/Dl+QSyimBAv6XLlD1WsAX82juy1MGmgCeZCQRehd1vykd3
TTSz1VyL2JQHQzHwlV4shxx6ioo0P9TpvhSAVhD6WaqjMwG1QjoIhx2jgjJ5P5oMk7Bjo+fMusOj
crE5tDUaLeMKVbdBELUaT3Y/eVPh9ODnVJhpoeSYGUmK1BW1662+6JbDsZGLGkvGFU8nDoFp6L4v
ql9rB/MVfjK0di+eQSih6N9XLXXjkvT9FLKmB4exoHVhOXtECYMmNoEDgH0sFoTNanRcIr96ajdr
5SthJRuVQy9b2vto/1ZYUzmDnX2QNWmhG9Pivzfg2p7s4eRgi5Yy28ap+MhdvdOD3r1viqJtSbYU
SEPVA4B7p+SWCCEpvMVfSHGVVdGJX/db5wSo+TSdZzW6LuhmFBGREYNJANHwQZFVchaNWFNCfFtP
2HXZgAkn1pe1W29G22bd6F9dIGI4mR3pext/Gmf/7v0p6tzCtkpZXoy+cQJq99msxjfdrqOapaFQ
VLoM1kbQQX4dH89DMQVtbySx9iTLSvJAlNKbyS2OJXz9xvi6HwiQ7nWfTh/LzsTLzBIN8lQilh3X
SQ2OPAjWkvK2NjlMUpiMGtI6CeXvnjLnE0rdsyu7ji0WgbtSj1vv/ir8AnHlQkeB70m4SYOTfhVm
2+53GHLE7A0+RqTwicKUSWAytU1lVKNWtE+0tyNnJJwzQjqaf9DGyY3IcNotQBwGZDz5yL22HNzd
W27GDDUWkTOsR7AdJdzyirbKtWbo/7chCODb2ll9VmYJemZofWsmkti57plDkooP9MBHg50cPHZQ
MCSMSM7+rVY1DXUy90kqWy65EoLEEFKxEI2eEEqkOJg+53xehP9bTq9p0niAzKdi37KnqKNztXhy
Tp/1xBFPTMupJGJM3A8qIysJamc3Q2tNVbt0dNQnBwBG4RxUPUhNekUZ0gHTXD3nipese1eM4DIC
uf53kiKZaL4RAYcX4xOEN6ofHQsF1SNK4Ecn3C/Wu1SQmRXKtTNe+TUBAtNcnmjCKeOQS5lRFvXQ
rEKjuVx5PnKN37ijMTxgU+SqGlv2wjV6zZZW0D54K3ZvXwgvdjiPOtkYIT9qOmOui9bWj3WwDhie
u9OT3V7vBlqirQwaCviiETIYGOi42De0BM9LBaPmjuUyD/3YeThFV/v+pbJlUmFHfNg8vE1IsFha
gvzY4YuA+Jkj5xI/z8+CamV+y+8h6UwM6cIFOHXoe7xSoUFwzzDFd7L7MTPrzvIfR+wNpFbTp9GM
J76AuuhuielSV4jyigOzQZR4/6dkdknioLLKLjR25pzB91z5pwPY0BMQ4RKIE4Ow32E4TXavqNYL
yPpXpdnktyF/dIFj0JwZutYVf+X3LsQDfCC8QQ8+Qc1ZazR6EDrGE46vaimg70LX8hCGZmij+9oj
56XTM16JnO7UHi6uwYfrAW2+R2ts/FY5yYTomAfYqbre6J8vt6q2s1m6Zo+/kdRck9nPRoaiup5M
nzhcWM2z61Hx6l7DqRg0UJfTv0LHfKw3iRTyxREhxcScuABzIOJO7IvoXU2fkllOxQW4KJJr41kP
8obHvX6duXI6VAqvI724asX7lWz1/kQktwe6Vo1H/icw0mIoeIF6grvrNx0xCCtoVMsTweUFIYYb
KU294macIJpp0Xw6fFrU+HJSnwR9gFLiy63Ry7mlQOoiU4UnU568EyIGHz2TsnuwkfEn3oWQ7wqD
v/0pHz3z8rFGWMxlLitbhq9xXQklv6VFupex27WI/odwOIgPYYmr4lJt/q9hpCcdi0QsaPFce1wD
Qm/fvz6EA+sLKDGvBEx71JfV/hB5MlmZw8Xrl0kg0yGm0Ta3QelYG4Kp395RIQBuvJhfySFgPLk9
x3Jtk/UZyFJ/d8F+ihGCaozjpjob+i4R8isxXoC1MPMgkCIhxNUP8XQjQKxeKjrlTNMIFnJqvJtk
lCqT5vB+LTWbE6TWGlNZMxNvWDQemBoAxlPJekbNokICQY9n0Cj2Y5EHob6yNzxWickgnZOcjp79
vApGgIoAL+OrdDfjqtoamcqgxVnOnR66lzA5deymnMiBILVeqGfgF1Hd+yW3I6eGpw3gpUZ19Nx7
4gBk/MewssMPeabAVfMnJt53FJYb8tuZ20N3Rm0fcc4o9hUHQMev57QVMczF1uHxiCuPAaPbST7f
ywMbb2g9aWwH/LZELl4U0D26oKvp6GkAa4Sfr77adv4wt1BuTMKSPGHnUIAtYVFayod81nzzOH5R
efIgkgpHf3Ywrx+aIarWnfvNnBqp2qpoku/lzoP6CQQkDXnPaK9wfM3lCpihqLFFX7FbgR9WtT11
w3q0QWn+/r3oEnhO+63cxRDcUwRgdYOT4fPKuKAGdpnv2X5btEc7sMgizzAlGWh8eKfsIAWo3tVv
nC6098QvSPZ80Me5WQ1FDKPdoLXg8op2kcOeGq72xUsqd4ZRxJCSo7ykgeYlPKoYX1kRb+PQPcWb
T5fEr5DfC10nTULT1gUPMcLiT7s2XPKppvzXkHwrGlJ2KWh1qqJd2WgLaUu8awtCiEihAL3CpZJL
EKChgZAgblz49dsZWlCtIWPSm+oLBGYmaZiPHH/XzwDtqS0mOYypUJyufb0cG5v6Kn0qtGFElRYV
HMEAEelZYAyU+Z0QOdlNwyaE6q+KJOlm+ZxCRgylsOCZXrP7462UkcI5rDMB2OPzpA3LtMekHOa7
68FibwgsWN/nq5R1aIAn8KqeX3hKx3xcgeeL5bNqwKmD/WxqIJIc2hOh1lGTbZnv1MzIFJBn7udF
wXIvMvq7FMFZyjZKDB3+jsAWrhsDPvTtLgSag2M5QBziOeakWyPDyo/uryPEoTg7zBE+zVLRESUJ
1O32pKyVCFLovap1GLqPXvw15olBvTzJPSxg2PsGt5K4i0LQvdPKafuEbqb5CnqO+KkmLzLM1TMx
bOR9H/OwQR18eZskELn6UViIrjCRm1I3Jvz2xX6hSJ3bYS11fwuzMG5LPxyz2LSpjmHh144+Qaon
tqocKwhKyESzLqtjFFf/njXkkAniQVZ0rG/7UTf7EpYsCseTPi1jEor7th6/wNVuoiErrnMvl8/G
d6Rx4CVpaE7m5h6HCtyRIgEMJ137hEjesJAWeUpdaayFlqs6aKVzgXLfrxqRC2gJOfMaKGGp7hrH
qNuH81iKKCQbL4380q7l3U3EH1wAjRupJIzwONF4WMZi0JpfRp3ysp+29J+NGc1Yw93GHPOTzwye
04jEdqQgUid6lHipD4NnDemlToEaQHasWtJVRaryJqEE3lALOxRZSSLeEcHVmbN0MfaGgWfN+nUz
Dr/UwWAjxuQoL+7LdyJ1/Lo0DUG4j7rHkiZf8tX6ffQUFGNVUjREjBOZa16p5BPC7R9iR4lhwnZQ
0PJaXWJK5hxEWtNXqHnT+T9Ru4B39i0UzmhA0Y/kmSQrqdEnKmQ3Feuax8+tpo8T6oWx/BEZQ4aw
h+Rw6Wh+KbZs8WAkWwtdc0issCMJUir5Np3Ywfn6MCvefSR/EumOPUMr+KmFmnFtggrBbbAFEsBF
AU71XCubQrNlWxIh386bGLf0ug7pFJZmLiac7o1+bOWPWf4C0jg0lns0w9Ho0OopVZ4NSwa8tXEI
9kgAWfutgvdvJPJ6KSg/xgpRr7QbUErnlxbjOppn+AdJp7ffJujHzwsQm0vmLMieIkMPXSrnwtLq
UyH/hfieaORRc0bK4BlR/YeOGLgJwGuiUJ6zxoLYDq03hamawpbuxuHeIKc7ANjkLMlAE4ooRqMA
gNb6LriYKY2bQpWkMWJF2aqdmEfU2zUVL850sSg9WVZxQRUfFu+HpJYm0QF/4tHBntFbRyf6GV6a
sqEhDagUOvzGxzWztY1D7IB1PTknpdvR5XCdLX5yCSMdHmcGIi6dzmzR6MYX7p4PkaZd9JYa2Owp
/T3N5KY44uIF5k/1vGBJWjqSx1dQhpmaX1dOQcOr9lDfTsH08r9qDRIKEFHATK1+/xgAXFFrA142
aYc91doiWwylO4Dz6lGzypIZMvMDwVlAeVjr2k3ybm/kV8oqvtiHxVHLEt2r8TM9CmdIfRk8TKDI
SPCmnCiPbeUPX5qBfMt+aWXPpxAqWog6JJ6tUHHNw7Yph7dmivJvjOyjjwQP47/7vwEbWqPFduW9
dtTiD1AnvqE58YEnQrev8W4craSFAWbwj2OACGHlTnyr9Hku07WQvnqsap42k89WzEEbm7Bc4O3v
4AvrIUNJCHxdunNoL+HH0PxDK7/TWrhfq493omg0Slr825a0vGHIjiHky+FTni5sLJTGIRCjn1PM
lqZ4FfdUw1GDU7GuSoQW+9ht8D1v3b33d3ULypjQt3tB5PCX4tq2xHneWT/vj55Cn6K+qgLfJaa5
yrv4l0F/dXXT5CZ2Y7Zfv9tPERautqNlgoLVM7hkQQ6ebCl/xvRoY7YdKrHdp3fSdsOIp445eEhc
H2iuR3/00NXt3DUClCbg7kmmzYq8pVTnIjqzecdmd1XTFs0XVv/Ec+L/yvC/qDTjWwnDOxtSfNMm
s97mgTJ1QdVs/yBuTnf/PzhwGY4M2iF2y6J37PINMDVFVUcIjr0c9aRjwHY6yQlB92jCQsSKbg5r
RYFioViIiWADO4m1lvq4E7Bv7rL10ons7kXworCUbeLwMkY49/LhVZs2XrgNXKrKodgIN3XKLBtH
uRe2zqjyE2F26kC6rw1PsiCl+LrI+hlV7QCfxScnZzdoL0gVGR3ZY7MY01jrJKzG2qRnGprATC7a
A1GyEK76WmuGl/ssJejaOq5aMoCGfmkYDUxFNsm9mU3BDR4nrbBXIbe55bQAv012Hq6GmFaTcFaz
DEt7Fxu7B6TP+fkYs0lWqSntdLWBLcBn1kVh6G/9yMNRK27stnLeaFYVtsoySowtO1XEIOKsf6zD
wLzcJv03OTn+WkNZyxEDFF8IUmvsrEcbD28xNZJS3rAwdiOAIxAK4bZztJnhnY65uoXU3ZKwDxx4
fbxDKRHzr0UY526kSpys+rk3E6LmIf4NONy750dcPW79QDhun4B81V1Hx05MEOuxBzBCezagZNa7
KXAY+SUFFV8PO+Q2Gc79fELzO29VzGwUnRMW1zjJVK8Ynrw5jxc84hGpkDqBrpw9tz9EsV1Orvvs
07iPOx4aV0sY1t0sbqe94E75qhfBMuoZ57+gXfGwAqqHfA3t9kUD8RhdVLxnSOHBH0TxorK4FBVj
G5i1REs+fqucEXZxRdFbGeLHPMWb5pbND9fRcjPMcPqNmuHBSbphvFrvv/Jl1u9PUaEPvOUMfOFZ
93ON7rpqy8YzSpbqYgFvVt8dc2SplBrpo7UmrGOa3K6yErPDInmktB71vKnWdKqyKd53/v0Yhg9X
CpdNxSPY0wS/N4oW20dHhFBgAoPHbPqatM3NPOuJPC5BFfIIPTlkkl8XCTcTo4UeO8yj+2FgjrVT
VhJnjfkOH/IDziISjcugw+QyD0BUIVOlMfbMfAu4+y6sbJw1ngENscZIeK9KwN31gS0xgp/KtxAh
kTQ7Oh8xCRQpitqix7flIGshOTctxpk2KIZgLB+pn9hfWHOzGYBecF/JA63JN31lwv6lotPqv01i
jwwD0Dy8tIbrYtqALTk9FMSTmb3aq8EOJOFsKDIkJ1O7IViA5WR8yNv4JMuokaMapimDIESAZlgr
sgD4OmhX8FOV4ZAHarAAAUrDKWPpezEdwjof26m3J/M74CJxOMuRERl9gLYgNBoL/A9U5f2ermed
XAoUklKEz06bnRfz/N1xqrd/RDiCsoQ7Rp2jQvCj9HOlPCO4fXs3Sda4/m1enXlONXtKBtSMcFcq
4aUFZws/u3MMEAZ63S2AmVLQKZlm7TsRfcK4rZkJZHfhDpgeRQ1QZzNfZfOQauAkHsy+XFVKy/G4
qzXNTOvJMwg3MIvbmSiw4HeWV1P6/0rhY3H5iq5orIaQinO5LSeNBnqsTYLUdiH4Tg0yHvHVf5Nf
jzFG/t1xmV6gtMT0OLg1ykkq3wqME46SgAVEyRRhCtc8fMWsyp0wH2jWV8efR73bJKYtSriHuq1p
WtydVYkIYPZlP08B0PgU1Lr0W9QV5pE+o9L//DDB9J10+ykdUaRCGht88OLOYuSUuu8/rEfEF985
FaBp387eS7rHHHplhJ4k0P8OcOLRfwk9JyIWpy8tGFRfpifzSpBfD1cv/sz2VY+xtrRhefqvoZUl
DD/s5INBLp6ypROpmroKsfg0wIW7dNe57x0ZIqwATglRpiwGXzYTwIr5XcLgBdtH7ZCncI/CuZXH
DcpbchTCkdupwc+TWn1GeUck8S46MXi1aWA3G1vGBI53F+Z5N5dYBr+zuLdqcNo1ZyVhJnJjwDbK
cNTS3wnkse8lMpxbUDCv9loKB8hW2Q+BhN1Uw1bxy0sOdQ7CVbtltr2VVdNVO9lC6nj9bk0yVNOW
krbWUrW70hRbdqPUe4/QiFi4916O5INqqmrnyaxjFMrWJBmljJDwPhgqeAxHFqegzEYCtilJ8PG4
m6ArHsb7JSdzFy/ie4ytiayvjK15FQNgBe9ldQk8ASsvJRXGMkfZ7CoqaACZCc1av4a6E3thOTsS
Q+stquywpVoNBVYL2C/XElYmu2PGwM5/GPezyiHjuPih7RSCPxdJ2GojYvgtfRyoTzcCZEzbgRhQ
Y5jEIYPPqLnG8oxswNktuRBem3pMsS8tTIMIoYnMHS5hDEg5ui8M540SzRqhFC9hDIXS3rLlYZhE
nAVwmweyx4n4MAelrsf6chzUA0GcSasYMMy+3kIEZYA3YaBOW+v2IU6U65UsO/ZqA+AHhP2gqUIq
2uwOcRO1H52Hw1Xep0ojevfOzQgtgIYAJbhKPnb00OcO2hjxFFSPdhsdZccv6D+d9wkm6ck3XgmD
L34YkFJzAtFnz11/k2KCdqYo52VqXS7P6X9U9JtqeUAvU0ZXbWqssYRMgC9uzQ9yrk6krRky2nKP
FW1xarLuL+4KfmgWXoXvY6TWthGdYh+z4TBU9LH+ScvQd7U+qmaY3ceTy1ACTamhzt+aa66Ipi/7
lu5YhzmUprTKIY6Hxwtumg4l5IPwliP5mhRZI/BI4Fv4D+c2MGfGVnmzlXbCT+wT4uX9e1Eq3QAF
+gGW+15KiAOOAL9NR7m6shOlkqgpfyfZj4kC5i5kQzXNzCiEQCa8Ep4qq0JgTQCm3HqTCwsaZe13
E0R++0iQcpC8fahee745xd2tJ3t/k/Gbi8QRJ2IBfpYQYTkUuBgvoG8CyzZS9Bjx+a9gGT6UrQDs
db+5zlaug2N3BzYb0b1MBvvVTKobecz4Nkid43nN9RHfeo4UtmiXLFyN0PFVsckCu8fvnqcbEUAB
VhFr7z7bBY7YH0K0bh2rkcTDfZj0hX0GqwiE9xkw/b3ULQa6jtvG6kOjTunXJWpPm9Yplk1it2tE
3XnqT8ADc57ZzpNGt0KC6r0nM8ss7ttgoSAj/WDzdSFM/5Qjon2vM0pMHSeB5/8DZpK50COmm6mM
nXQwLm/WJYnr8VFujJRCvQY+CRWw92/rGl5ARs8XEdXx+rwDeP27xpDfvWSiWRUXFTXq3TpbO5Dq
hHieprhvFrzu5tvYZ1+0Yiu1pGGfngeLJnlrwMbFz9JzTFOwGSVB/UNaRiaRid5bKiqFAyQu4yOr
MhuPzvKv2l3QRqKRz10xUWgpAE+5CC+gbs4c0qj8Q2swOztz9Ih8iQwYLCZ2C12vFHggzSvFumeU
btb8wbGb8tFcssYH43nRLeJydzatt0JT3zemzWnzIQ8gCD+P9Cxbuj+QgMh3SwLlhu8CmrEnMfUT
RayfIrE7jOB1MOnpfEEfbUw9cBS8bR29oJtNvM6KqhQSbXfQ9yqyKOjye1oqxZhGpJpOQ4JnSQy2
OyYKc0rIKhU5IWDIhIgW/J33Lznwt0rPQ4NemDl4WOntpFledr59h3crooGC9C5hLQBgOvCVr1up
ITLR2Y9TuQW+cupAwUINKE2QH9SsvQU+hzEWjbkFC1o//C8cA927U5Z7TZ3t/P0rDDCOmqzIdfXt
Ge81xSK4eNLrjdxbLtL3iYRH85fL5NRe4rhpIg2YySshohrSN1PLt84qv+pdCcpzrP/bM5qsHdNN
M82VapB25LKJecdyv4t6WFqTaNVD+jNkuv+vTF1SoVvsOfj2inSDbSwIUUeRceKGXdbB5mTBNPf1
53bX4vZkKTp1xn8xazAUAL33wVtXbfBdUElDZ5n86xkJLIfdxq0+tEyki+1c6MkcwDikltV1ipq2
Fr6dWWhn7LS9B8cPP2Y6CLiz+yDY59cdKi1WtbdPxk6edJBE5qw8XRaB7VxzYjiD65bPhTu1Zrg9
MFcFaRduseNGED065Pmft6O3hmL54SgFMbF9kWvruDp2oSToonkGl2SU9PxzOaL/ykSngxicZDje
PX8MmftZo9Kk42ZZtSbMHJ1d+zt07m+7wV/37FPdChWPeI3Fel2RpOC1W3qZB35qnsoiVQ4VzzYA
z89HcnTldI9NpcAX48pNka+YbTqbXZovnuKN/tglFTfES+0RVlVKYQPdklD5nPdPscH3SBxsjhbU
RT/diSjc8FCZzTioZOnaeK4WNxtyN1t8eK1KkPf7GZpgofmPUskZ3ALHwiTE4ubDgS4iqcjjnaxg
5KeEfmKAheLCqy+2kF66aouS2uzttlTsBEYSerdhWrvK4s+Ha3fEGbLQkoNsZwR/ihJdYFHwZ5CF
g5Gq0nnKEI7Ti1cUxUYDlECj4puRR3PqpX5TMOmtMYNEcxcxBhdAvPk6j4UgcdNuIkdAjT4iTz7J
eOGdsxEDsEGXylD1KemIVMle8RmP6/v+60wNdBh53kW8APQcagiyl5sfRfZqFBBVxFyTc/5tyBwx
N4MxM5UtCin1M5ZPTIdQePcXdx20SfPY0q03dZ7HYWImQGXEU07125wjyZ7G1rb4+V+c8Gs/o3gU
g2SOpUIK9qUKXXglg9StTy8XlE++BitYgqXzj/VxdOVGr+/yUL6sdivrfJMkojJWF4QE8Q6jp9Em
Qgjs6yoRcJt2FR1k7/uln8+1T16G8t6+DHvAfigZOYl+3CPTkciic8wZKK5CYI01jjb7klaJx+wP
SYLNnPscpu2guLQHepNdxh4/Lpr5QEf9IA5Zp62nA3HXy7e+vsfpCCkJCceKYAfb9q1w0aOzBQL9
rCLjoV+3NDB0+C7SULcVPKheBqVZxWA3NgfBfP4O73Pr9fQlW0HOu+Dn49nsz7VQYjAkZ/R0cOOy
SgyPYXmvl1ZdTKlPoLM2fzgFVJZeCY/bOwWXIzrBBFzgXvFe1Xf7NnZ4FeLzh+CpnO+ycnAFBLJE
562TP68wAgOmS46QoMXOyhRHE8g/ZtvG3052+iSo5oPEqzU2yozETeeSGYO/edcSTuIV+foC8hpF
t/KIqRrbDO8TFsGCxkZ1y1RgiBxaethHNd8NmHHtC1/S7RPPcdMNpqtDP+nl7Yw+SSRPwj2vQcF0
f6pQKPrd7R/fdnrtC83CJpj4PjJpeyXJc4cuIOFuiteCe77TLifssGrgbrYG4zYqHD/4i51+MMhC
MJMWZfjNH685MP3uVJl5BjH3HQpSz/7l1AU2peLYBu7y6oQuzMP+oC9GhY841z3rCq8fDq2OPR3u
aA13IDQrygWfaihRPhTVvtBOHng3XrYtYP/eVaOSHex6erhH9RVJWVazLnGDlWCCjQQrMWyNHC5h
jysW4oWcCZXHUfiTEXOVZJuPbJJACU4PwqugGRil/51Z6om8KH1RGLAKrNR78O5R3E0H8AnbxHv2
DOwTf+rhA95yuUTjJiMSpax1oPTG92U3IryB55hbgem5YVLqa9mJzpUIgnn3WhCYEcR2y0kh8dJ7
AWWVWieVUHOm+idWFVzlclXz/JETW7DeZb4q1aJzUp7h8QtqKiiCqesGULmQkXIQVpwOlf/VNe6v
XPGQpLCZQwmyLE/VWs6V55N9AIDwJN8t/bQ96rWOV7dbSlx3Zp4GtypVKIeNaLMw+gyRthZfm+E7
LerDgb/vpgdNP9xjB+Cb04431XtF+5jXe0/bRDAljZ3Ulm4YX3O3Hdnygpr0l4muThBqG+kxpa0n
zcTM407mG1bWEuJM+aYyCyuN0ALzLtaKR9zRGm/x9DGdfBDiGfnZXcwvi3n637il/rza6G87xWVE
W1S5kwNgw3CJqlzPYgxbrM99AVOrHpA7/RPAkpL/F8rHfzxQoY+hzlbOQJvVQKHOh+fyRM2np+Vr
W3dtqbLTBMyvJFcvZGVkv2cYvwS9zNlXQMVT3lBMGfpjS8MBLQrF4upIxMWjatsI6RupXaAl+aPD
sVC4zWgfv/f/osIB0FCXOx2MDHuoc9d9gA2/Mqvk+eTBMqDoUXoZHdt4b7L0IEDhTjrAeYA+01jK
XZiGRboUJKg/sB6JcCM6AcQ8iIzx/9GPnh5MO+xOm/IG4oCpWQa1MncTk2jXAZPbJACfN9hQoaoZ
XuJWFCG1XKJ1K3Z1bQ1aSRFnzVCIVTWjPwYFRMBkI80Su27E0YMqGYmPH8/Xf5tg75A94pmQB/hy
/oXaBrlFMYyyw+R+rn8OJDziS1xU7EZ67tF36/XDEU98ePLM1PLIaypBsLneC5B4k9CvdUHt1ShM
b4ZokBSEmL4wpqCACd2B1ZdSrTiZM/FWGtjoJrugaS49NtXFEEPD5ph3gvoRoI+zSYQTj5Q3/LMh
wNWdoaq7QonQF5P3X/gUm1wnBFL5UQXbWsgVhUSPEhzo+bQImxIeSEJPQj8Zuy0ZKKY549gwb9K+
iz8fp6D1DZ4QcYTuk2UqpDck9l0lUJlIXm7zxLBEX2vx7vN/LPJ25KeORrOmfY8s7RnRMs9KbBpx
il+faAF5wZ7YFCaLKI00SZZHL5I+Gv8hNE5AQRmf8Gj7h6nlXkGaIKs/6leEL4uLuxKF7NA60SRK
/nARgVw4Ppn/KUyAr23Z1/yB6IkDgMHZ860uirVmIvnSNUZvmI8lueqMEOR0/z+aiAdd3w0FFLWN
WQ+dTK0JZFHV0bOI1WhapgTVy4vaHA6Aok0mSxXRdJ+s6AS/r0u9VndJs1H1olIVESpNwQLipXZ3
ctWTCp0V5+lk9LNCOjA0u8X3grqd9xORwb2iQfL6PDFTBR80btsDLJpYyJyjlgtfOnQ4e7CzPXBj
Ek7omfBqIw8VsghHfuD4OvslN2E944wAy5wGeQFR/55c5n+Zt5R2+QiXryiXYm+V7Zhc9v/aKURe
TIxRyZqTbhaSAk9dWsxj3kXqx7jLThhgSgZ/52XLLOjqvSjqfMpC6UVu7f2cODg+ozcIu3vXQiLk
Ga9nxlEX6/10PGVzvek8qDBA3G00OxMhsYEmDsJ9o/dUW/gVPu0GkrKVq7RaziVbkGzbSG1PYMj7
85t1j/f6GnkHpXttiuDBbdOlw9lS+WNDcB38qGKK0OPdyw7xZbuf3EknrEx8lJrPgTHUAIbxSe9u
y2YAsNUy1SIwYur6qyBsUFmyim60W7Ekz+NkXieWxOexFftXRJfenM+LxpKo3Tu2YeUb5dPxtx4B
GvvFiIM3gAODlnd1hMU39+Zzb/MW1AH4/BQcSjblYZ4pdRt7WNWOHJNNC67ZEvR01HpAged21Yth
TDmMQ9pG6TQ4A/PpoTrCk9iwk4LXeTs65mpMVfY4UzAQCRkRVyjzrG9w0svi8oq4zJjUajXVc+zx
7m2CGa251oOz4Ahgqm2HwDz3Iygkt+725QpxQ4QHB7kl3Uuv0Ni03RjjJ44mOavpBAxZP2dzCBUE
8p+zuw4FhH75pEPUU+kp1puEzADFNGZMmafwT5TsKg39sQV5sDrp9An1UF3rZ18QGjgWApjzTgRl
HvQ/WKf5y5U3mgJ+zFx0SjKNmlmXludkEiAspWUp1nPVYQzHtrS7bl4qqmM1sKIiuX1xqswdCG7A
cJg+E90mMhwMyCJ1Ey9dNBFaLtB30F6PuxF+/a4Y7IeH/MbqyeOc0OrE9N3I9CQr/93U29MwHh12
VL0wFEU7U0mGl6/vJm8tKy4Wbni7RaTNOtkmMUS6Qm1N8S0CTWShDVpxG46mh4TBa/c+uNKalEi8
OhmzNy5Lfg0FS/UEpBtGO10Jo8abNWG7egCH7VuxRhoxXf6fHKbH4v2YdO7YmVtqHJ3Mn5/K5RMe
LrZ4YZ92h3ubEyyejJc6HKHx7Bo5Z2XLv9EV1/YpQmp8k99TbaHehJoPD2wQxoOjVgx2tW5/LViE
mFw9QpRA/afGTbC/jyUo+1eJHTsRoa85d/HYTKQIN5nRZY+MnmwWO+pfnmNZVHIx1e26wOLILzJ2
c6afO748griO6/fpxBb5Sl7nOUt2bKWQJCDy03Zu0l0Op5RJ+97F7Gy8Xn7Nbyh6qO99HX9pFiMr
1E206O7nvgf7kfF1rsLzNlEQWo0VcuzaGGBVVN5rwRe/Fd0rFHf0hKs2mBacNXjBESoiVU744Dbc
IlKXd7BziNKHs1nFOj/edni16X9iDJIlhS+IFeRnsR7O68Fa5N8YW5/vGZvKXIO6cH8jz4zb0HrO
nTaPt2rZMJ6GJO2FPhUuPdGVIRhe7ZIQxb+Ex9A7gak/NOHg7pDeacZJnU5ZSsctApMCThdqSLT/
D/M92qVt8gYn8yEbf8uno/qsdT8GVIVhjBh8G6VxdW015caDmLGe+S390+OlovPq98Yj8GWxmQxQ
kbp65jwO5Ap1BdBDSY9+Z3mC8rtPlgKJEP8gL6lor+Ld8yK+3q91cEzd/JT3/AdmkY9Sw7UDYkuU
M3G2nZ8sO1k8LMZl43Y6RCJEqnC7C9qksIUymK7ThT0cMpuXAPg9ZVsueBiMvSOVU1pjwyHmyiJW
qkw0iiVeUyV89Zjx/AxwPm6HY0/n8tXB/IjAIyV2l539DfEelAYADIhA5A36qYBtIYenZYXTtjPN
JN6I6GX+7Voc1pl9TwDtQOJXcOLbMljz90Fx6i5uCb2aeFVM2fgpc2JTHKJt9CA09iomKTgIrl4S
VebEq1+/oKMi3oPwoTtwelyTUezvLrYdJ+3spbnT0b+pbzaf+ZG4YdrIUgcNRGBDoOiYTJqFjSMQ
n2IpkhVr0StDJ83u7061++wtYR4K5zW4IKGHDxQp+2lBPcNuT+gQi3ExvMvvMrUl+7miSiAapqP7
pYoc+0jk1MykLCJYARJfqYv767e4giaNaqPw2JNRVRpjEELDCo9N5wUGzdDAAvBSwr5rg4SN1are
5m78TX2dgeUYb/6UQMULRj4jWk3V2vmmS3NxK9PP+dUn4REC9XdBPxmfyvyaDQ7JhrAC1df56cPc
/TZrBLPQci+fECenXhxYs4/mf8+142vkL66I449eQ8sKHSVALisqLSfpifBmKoPG5pwrqoBwqoVY
xQs+1+tNOz769mILCYgTDfQI8Ymz4sj7E4Ty7/0SETnuTtfysh3FvUlv+R+JweYtsfMXVlD/KUWr
ElJP6cXH3XdarQGijRKNiGmFGTPrY8WTXZyB82mxS2+75x63AlMNbN5k+erQPLOrZrUrlsrnR4tk
9Rynw1VHZClQd2eUAQH5sEMFbuOlURGDePfwSGpvKhcvJ8+eb3xEdDIhWkfowkC/skpHjf/zJ5eS
GnkXM5SdPeE7V5raUboNS+SDssQYniPrKdS0w+Y65DR85DxkqTK9siAheGONhc9X5pgEhCMYQ8wn
nT41xI4id7tJVAZ04FdbqQWJcFQUGBuIrEqCUKgxNVAIU1TXScf3XPsDVu8kW/xDZrIenkyYMnKP
dyuM0y7HUS3ulHQ3HOjM0xT/vA1n8aZJyaLqQpgZN3Gmgsru2zRxteDhY75FFD5susdLieuP4T4P
7OKwgVBDh0s2cJ13L38u3WD2V9hCaTt81iOglTPrEh5qdXnN6DzLbMb+oIPhGlI5oFkbjZTxfIpB
1gWkcCh/yg6tynqx7DJV3h1vXfB0nMZFNTKgB8K8w8bMRNhsccm9E3t5KUd1LCpoBcOx5miWualJ
/rfa1xnlrse/lit3BVNCRoUbTJBA8Ftj9/n20hc1cnn47LIBo5e5XrvQB50OBABRm1ev4hwzZwWy
k8LzqRTUiZw6otA8EqvSnZSY8PWHaCzyhZ3APP2i0e8vyjeNoeWhDWEC2HdKvTANMun24kEaEqhX
lxgNI7a4yfysUTo6dLQ6E7zrPHBlGHYDMW6pbcu4B/b5PLd8GoxC/nwYkl/tCQq6UMCe+wVtmLgF
BV8YLMO+Gt2av97su+sBXPrV3hUK9e0up3VjiStfFLRF6Ee/eBA3KU8pbukPkIujPq1lmCZwkI53
LP17Pw4iK8IcGmjP7UJ3BVCkECvetpc3tdDLJSuY/UxtGMrBC1kRR5ht385JN6uLXn5aoXBjQ0h5
6F+ZVEKbroVw8/RGZ5QjkrzG1YMuoZfdhzgo3dTllP8ppUd6lywqfNpn/6GbTahnz5K0r3zmHrPV
d2UqU3KmR1KL8mLQq0ptS0J423CV+ypyLT1ScK2PUDZvSeCNGE0/iDned2te3T7MLTGRQkiOJ330
bUJ/eL+sF/8IO6BQxkS8hadvUe73S6eG//i6GJwrO6hZ0pdU5+WUrMHl/L/3ema3TOYIJUZUwdlE
/OnnqHkx1Zykhh/ubwCscWZM+XgyPQtcMX9GYeD/MVwfhIHyedwGeWSnhna61ZrbNQ6Lbf1K69ey
BLl/iA6/HKn41gXcRneKkTQjI4NqNVgOMHlPFMdHE857hz9sV/Yk/3d36B1EhMBmD3S5fox3TGdd
gU/M7mB3rY5jl51mA80wG5gTc0ibyx6BCvjcxnipWx8vaW0ra1jZa/+BkokuM8fxFkAqfZvsgkw4
UWVUkkL5p9sWTIrbwKQj56Aq+hy/yv8rGarL0B7Rbr5RfKnTtn7YqhptlZ3MQDjs1AwU5jQbHx2w
uIZ54S4g8s9ncFOpNVvQsk0n0fkLGzkK3GDUdKYhGRp8cBciGpPyVgBRKfdnN53gVDl+CQUiB3G0
Ez89AyXZvzt1OTxnZ7FUQz7bxNqgTnG1cB8SOBQppV+k+RdMCFaiz7e9eEtwea2m+loq3Y/NgIat
nL4wxGYkjPRLKZox8TmzKpoMxdHsHCDDiV3LovPq+oaAlvNTp1tvQ0440YvMbAU9RjfnakwytWzv
6Rr0ztZK6oIBy1cqVAyIrkOU7DGgJteWkZiNQV3bblPoXGDpWk8EngWOBzR4OR6LgHdpED9FyzrY
rKBEA7x6JgLPI460Bd095DrcbOaf2u15YnXIqiR9TSRDuf8u4VhXQ/2FHhGzhVh2rAhsODkKVK3H
yBGcshLtDAHubbsdFZp4c/z19saCRWj48i8Lsv9YOJRdKETifVEAXxlHHzG6Tx7g2ow2k6lp3z1n
G0ObcPG1T6qAvrMV6orMfdBtauMJhhJn9y8vt7+lNq1abBTNDQTcZEtrO6dIM8dkwyz15wOVxaf5
U326CI3kubBlwjKEcDu75+tHmbCrqhOd9zy5n7upWdAdHwTrM9jZa+WjISDBjXxUMxJ07gZaAfpo
DsivTS78xNVHW5nUv6lDqPn9iMLTATVB7+CfVsp6ACyyV7BdYf2HvkbuSVLlDQmkWOexoBmEv2YF
solDZctHQ9l7RA082p2fp5HWuGuDfvp5kT9tZif0KJe//WUE3V8a21+XL+Vxmj+Gtn0NZ9m9hIpj
T1wgTAOLInER/vbbLFZ42KCSxSCcAC4qsf1owUy5hMf0HKD1+gQmSybAG4gNE/ykY6WxFA72FTFv
4lhWNWCXVb/+wfT0FWJbmOr1tZ+8scQWnWIgWv8hjbn4UJ28R9npdW1yLam7CUV2r9LZ97jl20u1
gw4uImaWnpj92NqRTc+AucwsQWU6iLAL5mYbuV7uxlRyBaPAcAJjvm8ILCxt8mO++b0O+OebSLDG
DNHVi/cCVq2mrS2qcu34tCuoIsk0PpE3ebIZfz6D0GWt8VG7YWeKg5yLG5NOR8+5LZCCJDS3SpCs
BSSZnnt5Na/sqqv1zTQoNOotaY70Y7nrrP3Lu70NxJoJd+h8Gb/+TkqSEsFEnIxY082VZ6Xx5NPm
JAaLllwR+vwN4C+fv0qachzg4KFmuFJAonKEvoTAMau6/RIUR1iBQOeEeyP0Ap5/h8b8sIHyFj60
Q+SFuid2PB+LPN5VVlR5TEYbDhzT9RYC10SVj3nACIvikKgoYM7allO8sbDpJHJNX6a48Gp5ejlu
o3YeN0qSAxSgm3XJ6VJEQmutmGSUt1XNw8qC3V4XMBFavVLFN/j9ghlKOhyWJOfmOERiACNFzlqj
CQzRSkIZY1T31ZmQq4F+c9K7tdV67xDQ+UiAVb0YN2CCh8+roW1ui7NEOPsBmuaiScLYoWuG73r/
MbF3WAADiATNmnSMgn3f2dfRNLITY2jO2flmkU4VQnlCiEgzC/k6LQnjfYJPHd/60g0GrXWkHDwC
ktMJWBhpEH9HKcqNb5zgbzOrThtELekeWdZvgn4qZSOGcMmhFrr4VRDflAyGqlV24UmB01We8ebr
Yu5i18dtBVRwT0jZBrTu3EKE7AAm6RdNcWaIdKSpnf9xf9+npXWSb3hog6rLcX+fUe/6bOgxiWcr
f0Cv5yeqMYuENt0+7pyXSVfHFfKv02zyk1DWn0krU/30PAFPYQAQKSvftSWDOFcAteiUoAtOKkVW
DxTS+AumwNx0uxN1oUJ1BONo6CwBAPj9FlyAws/FprIUSSebYGVHeQOPEBqwwY7278TaW3Iatxry
UofzvJJNa/qfGb+Qdk7kL9QsmnJsFV9glC2V/XdEeW8IBMAkryvVqK0nJIsRcJFB0qum+ZknYyK6
e6RgDgaZqh57dot1pj1qhiWvjd79OYap2FwSbleMgUn3BRVpHYTaQCgDMxfHQPBVTORB8d1dFIov
eWWMER/A7X/4d9qoRL0VGWdLHxRTw8IIR2RSSaGE4pMNY5aOOcnPzuyHbErtbKkCTxE/S261dBm6
eBLen38BeVnwZHutCBfiQjyuxwrgBtOgv3T763+vExlCifdkxAsAT+ZcMjlmY0svIgDnDhq5ItyX
kDw5XAkAa7UWvtZBG8CyzIpx4K9Jn0EwHHJGak6/3EXp5KW+WXXgvSsr3W6i9nPH0lmNyNxU9iuQ
UfXwy5gQcbIV7Jk/CJxmyG0GOZJ9Ny0LfT3Sch4UotdY6uSqFzqg0v1vAswBTICLVsYHZm7vVT8O
F47Tca4sWvMxoV7TleRJJlf8YdvczvBfoq/KqAGd78iTeFuzuMPm4JpROyTeifwjAKfmTBV6dK1O
fD5OokuqRu+cb4u9aViZ8oljmtIzVe2Pni1Yv3gfI1QpIih86qLytHO8rykUSid0So3vC9NckvTg
6fE8vbeT1CG5FyPkUjpJG3cbuX5a9qL7VzQOWsu4/1TrXRZFhs4mNYCg0r/3Uk1LTobE0SO9wIxB
cPgZ3YElwJEMQl1fqQvdOg0U9V24F0vVHYq+BOR/XDd/AjunxPEhZUf0u0pKIaWhgQ0/aulKu9YU
QtnLZ5QqOG+AzhBiEizKqdhQiC7O3EEzl0mx95v3ngA1wWJZjxX++F0ezPX6r7v1ha7rVBhutzBD
rilZKraU1dUae/uYlEyb8tbS+HHgI475NEj5V2jk1wvfLPXma/06PtahDzrdUxunJO2LmYtFPFNn
Gi1GAu1TKBLGrB4W1a9UorqjV/qRNJtRNQks4PVhaNNRP1Axbm0ov0CLOUV/o9z9RqAMFTH6BQIW
63JNvWq0jCXGQ/YIhmJkwpxNh/GANUiNjk1+OV78lA23dXk9iu03pjwj5Hmdsmd5Rz5hWYWesdut
7Z7aqpQZFe2tQ3tCOcmGKuv9QKaFsjn73Tdgpa7wo/yWUYkddR6Xn/i0cjSsr+YGRvBpKd9OZyUo
2d2rA5kf8576A9ufwsLtzwgCx/d9LdpPXNaL8AFBF4kMz33PJMqN1nTMnAFh1mGQkprzV8VsM6m1
1MsIms2PuvCsF1UYri5dOIqoPRz6Vn8dQZJruIpcdujbB3CLP4zdB0jP49fH5WUFyy+ww505vMpE
UxD4vEcDEdlJpSa1aEoGUqHeM47td01XOpYqRpxDtzVlr5LA082pXI34Uhx+47wxY/7YQjXjZDVe
ouSqY9ut11DMrxXjCvPHag8eex9JjIyMHfE8cyTR7AazaoCCE6ca8jurIWBvNhmcz0Og6DpM4hqB
j88etXnou53OewwOItWq87BjR1LA1ZW2Do0tAk3QK4DPkAj3bfkaK93TKYT0Fb/YrOJZ1w2qI7zK
1K+bF1o1vSnjRPREtfC8fcJJildnToyxcku4SLKJouxlf9RAj/nhGjRLWcz/adoIzI/DE+gAdnjx
niWi2+MYjwzcXj4xi7Kr3i7EDU11BZkskMO+r34qHCPKS6ZDA1zkhGC9dFDjTjK7Wj5wVLOkkL8m
V1/0NV5iM+R5pR4KnOv8vYaJr29EzI7FnvuwHzDzFplCOmY2D663jMa7PN6EIf5A4mhhcUp6OSZt
/j7l7PPhEbLPz2iD0wLAOFXYwHw+CqFMD+2ttEdVjsFDCAUY/3qiGI7o7uWMDvRigMG6v04yAPOJ
GpdxPsGheHcalzyxoyfJY7hmXo4p
`protect end_protected
